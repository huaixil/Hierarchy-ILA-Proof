module DECODER(
__ILA_DECODER_grant__,
clk,
eq,
irom_out_of_rst,
mem_wait,
op_in,
rst,
wait_data,

state,
op,
mem_act,

ram_wr_sel,
ram_rd_sel_r,

src_sel1,
src_sel2,
src_sel3,

alu_op,
cy_sel,
psw,
wr,
wr_sfr
);
input      [4:0] __ILA_DECODER_grant__;
input            clk;
input            eq;
input            irom_out_of_rst;
input            mem_wait;
input      [7:0] op_in;
input            rst;
input            wait_data;
// output      [4:0] __ILA_DECODER_acc_decode__;
// output            __ILA_DECODER_decode_of_process__;
// output            __ILA_DECODER_decode_of_stall__;
// output            __ILA_DECODER_decode_of_step_0__;
// output            __ILA_DECODER_decode_of_step_1__;
// output            __ILA_DECODER_decode_of_step_2__;
// output            __ILA_DECODER_valid__;
output reg      [1:0] state;
output reg      [7:0] op;
output reg      [2:0] mem_act;
output reg      [2:0] ram_wr_sel;
output reg      [2:0] ram_rd_sel_r;
output reg      [2:0] src_sel1;
output reg      [1:0] src_sel2;
output reg            src_sel3;
output reg      [3:0] alu_op;
output reg      [1:0] cy_sel;
output reg      [1:0] psw;
output reg            wr;
output reg      [1:0] wr_sfr;
wire      [4:0] __ILA_DECODER_acc_decode__;
wire            __ILA_DECODER_decode_of_process__;
wire            __ILA_DECODER_decode_of_stall__;
wire            __ILA_DECODER_decode_of_step_0__;
wire            __ILA_DECODER_decode_of_step_1__;
wire            __ILA_DECODER_decode_of_step_2__;
wire      [4:0] __ILA_DECODER_grant__;
wire            __ILA_DECODER_valid__;
wire      [1:0] bv_2_0_n9;
wire      [1:0] bv_2_1_n15;
wire      [1:0] bv_2_2_n21;
wire      [1:0] bv_2_3_n6;
wire      [2:0] bv_3_0_n124;
wire      [2:0] bv_3_1_n122;
wire      [2:0] bv_3_2_n123;
wire      [2:0] bv_3_3_n121;
wire      [2:0] bv_3_4_n125;
wire      [2:0] bv_3_5_n230;
wire      [2:0] bv_3_6_n490;
wire      [2:0] bv_3_7_n119;
wire      [3:0] bv_4_0_n823;
wire      [3:0] bv_4_10_n961;
wire      [3:0] bv_4_11_n965;
wire      [3:0] bv_4_12_n886;
wire      [3:0] bv_4_13_n850;
wire      [3:0] bv_4_14_n933;
wire      [3:0] bv_4_15_n894;
wire      [3:0] bv_4_1_n957;
wire      [3:0] bv_4_2_n848;
wire      [3:0] bv_4_3_n826;
wire      [3:0] bv_4_4_n828;
wire      [3:0] bv_4_5_n852;
wire      [3:0] bv_4_6_n913;
wire      [3:0] bv_4_7_n866;
wire      [3:0] bv_4_8_n906;
wire      [3:0] bv_4_9_n880;
wire      [4:0] bv_5_11_n283;
wire      [4:0] bv_5_13_n307;
wire      [4:0] bv_5_15_n149;
wire      [4:0] bv_5_17_n45;
wire      [4:0] bv_5_19_n302;
wire      [4:0] bv_5_1_n47;
wire      [4:0] bv_5_21_n146;
wire      [4:0] bv_5_23_n51;
wire      [4:0] bv_5_25_n152;
wire      [4:0] bv_5_27_n67;
wire      [4:0] bv_5_29_n294;
wire      [4:0] bv_5_31_n143;
wire      [4:0] bv_5_3_n138;
wire      [4:0] bv_5_5_n278;
wire      [4:0] bv_5_7_n280;
wire      [4:0] bv_5_9_n299;
wire      [6:0] bv_7_107_n225;
wire      [6:0] bv_7_113_n76;
wire      [6:0] bv_7_115_n403;
wire      [6:0] bv_7_11_n208;
wire      [6:0] bv_7_121_n79;
wire      [6:0] bv_7_123_n213;
wire      [6:0] bv_7_19_n389;
wire      [6:0] bv_7_27_n391;
wire      [6:0] bv_7_35_n408;
wire      [6:0] bv_7_3_n210;
wire      [6:0] bv_7_43_n394;
wire      [6:0] bv_7_51_n418;
wire      [6:0] bv_7_59_n219;
wire      [6:0] bv_7_67_n156;
wire      [6:0] bv_7_75_n411;
wire      [6:0] bv_7_83_n216;
wire      [6:0] bv_7_91_n55;
wire      [6:0] bv_7_99_n222;
wire      [7:0] bv_8_0_n247;
wire      [7:0] bv_8_100_n681;
wire      [7:0] bv_8_101_n382;
wire      [7:0] bv_8_112_n109;
wire      [7:0] bv_8_114_n367;
wire      [7:0] bv_8_115_n100;
wire      [7:0] bv_8_116_n675;
wire      [7:0] bv_8_117_n181;
wire      [7:0] bv_8_128_n88;
wire      [7:0] bv_8_130_n326;
wire      [7:0] bv_8_131_n29;
wire      [7:0] bv_8_132_n38;
wire      [7:0] bv_8_133_n228;
wire      [7:0] bv_8_144_n687;
wire      [7:0] bv_8_146_n184;
wire      [7:0] bv_8_147_n27;
wire      [7:0] bv_8_148_n589;
wire      [7:0] bv_8_149_n377;
wire      [7:0] bv_8_160_n370;
wire      [7:0] bv_8_162_n355;
wire      [7:0] bv_8_163_n424;
wire      [7:0] bv_8_164_n41;
wire      [7:0] bv_8_16_n94;
wire      [7:0] bv_8_176_n329;
wire      [7:0] bv_8_178_n168;
wire      [7:0] bv_8_179_n908;
wire      [7:0] bv_8_180_n61;
wire      [7:0] bv_8_181_n58;
wire      [7:0] bv_8_18_n73;
wire      [7:0] bv_8_192_n135;
wire      [7:0] bv_8_194_n165;
wire      [7:0] bv_8_195_n794;
wire      [7:0] bv_8_196_n592;
wire      [7:0] bv_8_197_n199;
wire      [7:0] bv_8_19_n584;
wire      [7:0] bv_8_208_n193;
wire      [7:0] bv_8_20_n559;
wire      [7:0] bv_8_210_n196;
wire      [7:0] bv_8_211_n815;
wire      [7:0] bv_8_212_n556;
wire      [7:0] bv_8_213_n70;
wire      [7:0] bv_8_21_n171;
wire      [7:0] bv_8_224_n82;
wire      [7:0] bv_8_228_n550;
wire      [7:0] bv_8_229_n350;
wire      [7:0] bv_8_240_n85;
wire      [7:0] bv_8_244_n553;
wire      [7:0] bv_8_245_n178;
wire      [7:0] bv_8_2_n64;
wire      [7:0] bv_8_32_n91;
wire      [7:0] bv_8_34_n32;
wire      [7:0] bv_8_35_n575;
wire      [7:0] bv_8_36_n667;
wire      [7:0] bv_8_37_n313;
wire      [7:0] bv_8_3_n581;
wire      [7:0] bv_8_48_n106;
wire      [7:0] bv_8_4_n564;
wire      [7:0] bv_8_50_n35;
wire      [7:0] bv_8_51_n578;
wire      [7:0] bv_8_52_n670;
wire      [7:0] bv_8_53_n316;
wire      [7:0] bv_8_5_n175;
wire      [7:0] bv_8_64_n97;
wire      [7:0] bv_8_66_n187;
wire      [7:0] bv_8_67_n190;
wire      [7:0] bv_8_68_n678;
wire      [7:0] bv_8_69_n360;
wire      [7:0] bv_8_80_n103;
wire      [7:0] bv_8_82_n159;
wire      [7:0] bv_8_83_n162;
wire      [7:0] bv_8_84_n262;
wire      [7:0] bv_8_85_n319;
wire      [7:0] bv_8_96_n112;
wire      [7:0] bv_8_98_n202;
wire      [7:0] bv_8_99_n205;
wire            clk;
wire            eq;
wire            irom_out_of_rst;
wire            mem_wait;
wire            n0;
wire            n1;
wire            n10;
wire            n1000;
wire            n1001;
wire            n1002;
wire            n1003;
wire            n1004;
wire            n1005;
wire            n1006;
wire            n1007;
wire            n1008;
wire            n1009;
wire            n101;
wire            n1010;
wire            n1011;
wire            n1012;
wire            n1013;
wire            n1014;
wire            n1015;
wire            n1016;
wire            n1017;
wire            n1018;
wire            n1019;
wire            n102;
wire            n1020;
wire            n1021;
wire            n1022;
wire            n1023;
wire            n1024;
wire            n1025;
wire            n1026;
wire            n1027;
wire            n1028;
wire            n1029;
wire            n1030;
wire            n1031;
wire            n1032;
wire            n1033;
wire            n1034;
wire            n1035;
wire            n1036;
wire            n1037;
wire            n1038;
wire            n1039;
wire            n104;
wire            n1040;
wire            n1041;
wire            n1042;
wire            n1043;
wire            n1044;
wire            n1045;
wire            n1046;
wire            n1047;
wire            n1048;
wire      [1:0] n1049;
wire            n105;
wire      [1:0] n1050;
wire      [1:0] n1051;
wire      [1:0] n1052;
wire            n1053;
wire            n1054;
wire            n1055;
wire      [1:0] n1056;
wire            n1057;
wire            n1058;
wire            n1059;
wire            n1060;
wire            n1061;
wire            n1062;
wire            n1063;
wire            n1064;
wire            n1065;
wire            n1066;
wire            n1067;
wire            n1068;
wire            n1069;
wire            n107;
wire            n1070;
wire            n1071;
wire            n1072;
wire            n1073;
wire            n1074;
wire            n1075;
wire            n1076;
wire            n1077;
wire            n1078;
wire            n1079;
wire            n108;
wire            n1080;
wire            n1081;
wire            n1082;
wire            n1083;
wire            n1084;
wire            n1085;
wire            n1086;
wire            n1087;
wire            n1088;
wire            n1089;
wire            n1090;
wire            n1091;
wire            n1092;
wire            n1093;
wire            n1094;
wire            n1095;
wire            n1096;
wire            n1097;
wire            n1098;
wire            n1099;
wire            n11;
wire            n110;
wire            n1100;
wire            n1101;
wire            n1102;
wire            n1103;
wire            n1104;
wire            n1105;
wire            n1106;
wire            n1107;
wire            n1108;
wire            n1109;
wire            n111;
wire            n1110;
wire            n1111;
wire      [1:0] n1112;
wire      [1:0] n1113;
wire      [1:0] n1114;
wire            n1115;
wire            n1116;
wire            n1117;
wire      [1:0] n1118;
wire            n1119;
wire            n1120;
wire            n1121;
wire      [1:0] n1122;
wire            n1123;
wire            n1124;
wire            n1125;
wire            n1126;
wire            n1127;
wire            n1128;
wire            n1129;
wire            n113;
wire            n1130;
wire            n1131;
wire            n1132;
wire            n1133;
wire            n1134;
wire            n1135;
wire            n1136;
wire            n1137;
wire            n1138;
wire            n1139;
wire            n114;
wire            n1140;
wire            n1141;
wire            n1142;
wire            n1143;
wire            n1144;
wire            n1145;
wire            n1146;
wire            n1147;
wire            n1148;
wire            n1149;
wire      [1:0] n115;
wire            n1150;
wire            n1151;
wire            n1152;
wire            n1153;
wire            n1154;
wire            n1155;
wire            n1156;
wire            n1157;
wire            n1158;
wire            n1159;
wire      [1:0] n116;
wire            n1160;
wire            n1161;
wire            n1162;
wire            n1163;
wire            n1164;
wire            n1165;
wire      [1:0] n1166;
wire            n1167;
wire            n1168;
wire            n1169;
wire            n117;
wire            n1170;
wire            n1171;
wire            n1172;
wire            n1173;
wire            n1174;
wire            n1175;
wire            n1176;
wire            n1177;
wire            n1178;
wire            n1179;
wire      [7:0] n118;
wire            n1180;
wire            n1181;
wire            n1182;
wire            n1183;
wire            n1184;
wire            n1185;
wire            n1186;
wire            n1187;
wire            n1188;
wire            n1189;
wire            n1190;
wire            n1191;
wire            n1192;
wire            n1193;
wire            n1194;
wire            n1195;
wire            n1196;
wire            n1197;
wire            n1198;
wire            n1199;
wire            n12;
wire            n120;
wire            n1200;
wire            n1201;
wire            n1202;
wire            n1203;
wire            n1204;
wire            n1205;
wire            n1206;
wire            n1207;
wire            n1208;
wire            n1209;
wire            n1210;
wire            n1211;
wire            n1212;
wire            n1213;
wire            n1214;
wire            n1215;
wire            n1216;
wire            n1217;
wire            n1218;
wire            n1219;
wire            n1220;
wire            n1221;
wire            n1222;
wire            n1223;
wire            n1224;
wire            n1225;
wire            n1226;
wire            n1227;
wire            n1228;
wire            n1229;
wire            n1230;
wire            n1231;
wire            n1232;
wire            n1233;
wire            n1234;
wire            n1235;
wire            n1236;
wire            n1237;
wire            n1238;
wire            n1239;
wire            n1240;
wire            n1241;
wire            n1242;
wire            n1243;
wire            n1244;
wire            n1245;
wire            n1246;
wire            n1247;
wire            n1248;
wire            n1249;
wire            n1250;
wire            n1251;
wire      [1:0] n1252;
wire      [1:0] n1253;
wire      [1:0] n1254;
wire            n1255;
wire            n1256;
wire            n1257;
wire            n1258;
wire            n1259;
wire      [2:0] n126;
wire            n1260;
wire            n1261;
wire            n1262;
wire            n1263;
wire            n1264;
wire      [1:0] n1265;
wire      [1:0] n1266;
wire      [2:0] n127;
wire      [2:0] n128;
wire      [2:0] n129;
wire            n13;
wire      [2:0] n130;
wire      [2:0] n131;
wire      [2:0] n132;
wire      [2:0] n133;
wire            n134;
wire            n136;
wire            n137;
wire            n139;
wire            n14;
wire            n140;
wire            n141;
wire            n142;
wire            n144;
wire            n145;
wire            n147;
wire            n148;
wire            n150;
wire            n151;
wire            n153;
wire            n154;
wire            n155;
wire            n157;
wire            n158;
wire            n16;
wire            n160;
wire            n161;
wire            n163;
wire            n164;
wire            n166;
wire            n167;
wire            n169;
wire            n17;
wire            n170;
wire            n172;
wire            n173;
wire            n174;
wire            n176;
wire            n177;
wire            n179;
wire            n18;
wire            n180;
wire            n182;
wire            n183;
wire            n185;
wire            n186;
wire            n188;
wire            n189;
wire            n19;
wire            n191;
wire            n192;
wire            n194;
wire            n195;
wire            n197;
wire            n198;
wire            n2;
wire            n20;
wire            n200;
wire            n201;
wire            n203;
wire            n204;
wire            n206;
wire            n207;
wire            n209;
wire            n211;
wire            n212;
wire            n214;
wire            n215;
wire            n217;
wire            n218;
wire            n22;
wire            n220;
wire            n221;
wire            n223;
wire            n224;
wire            n226;
wire            n227;
wire            n229;
wire            n23;
wire      [2:0] n231;
wire      [2:0] n232;
wire      [2:0] n233;
wire      [2:0] n234;
wire      [2:0] n235;
wire            n236;
wire            n237;
wire            n238;
wire      [2:0] n239;
wire            n24;
wire      [4:0] n240;
wire            n241;
wire            n242;
wire            n243;
wire            n244;
wire      [2:0] n245;
wire      [2:0] n246;
wire            n248;
wire            n249;
wire            n25;
wire            n250;
wire      [7:0] n251;
wire      [7:0] n252;
wire      [4:0] n253;
wire            n254;
wire            n255;
wire            n256;
wire      [6:0] n257;
wire            n258;
wire            n259;
wire            n26;
wire            n260;
wire            n261;
wire            n263;
wire            n264;
wire            n265;
wire            n266;
wire            n267;
wire            n268;
wire            n269;
wire            n270;
wire            n271;
wire            n272;
wire            n273;
wire            n274;
wire            n275;
wire            n276;
wire      [4:0] n277;
wire            n279;
wire            n28;
wire            n281;
wire            n282;
wire            n284;
wire            n285;
wire            n286;
wire            n287;
wire            n288;
wire            n289;
wire            n290;
wire            n291;
wire            n292;
wire            n293;
wire            n295;
wire            n296;
wire            n297;
wire            n298;
wire            n3;
wire            n30;
wire            n300;
wire            n301;
wire            n303;
wire            n304;
wire            n305;
wire            n306;
wire            n308;
wire            n309;
wire            n31;
wire            n310;
wire            n311;
wire            n312;
wire            n314;
wire            n315;
wire            n317;
wire            n318;
wire            n320;
wire            n321;
wire            n322;
wire            n323;
wire            n324;
wire            n325;
wire            n327;
wire            n328;
wire            n33;
wire            n330;
wire            n331;
wire            n332;
wire            n333;
wire            n334;
wire            n335;
wire            n336;
wire            n337;
wire            n338;
wire            n339;
wire            n34;
wire            n340;
wire            n341;
wire            n342;
wire            n343;
wire            n344;
wire            n345;
wire            n346;
wire            n347;
wire            n348;
wire            n349;
wire            n351;
wire            n352;
wire            n353;
wire            n354;
wire            n356;
wire            n357;
wire            n358;
wire            n359;
wire            n36;
wire            n361;
wire            n362;
wire            n363;
wire            n364;
wire            n365;
wire            n366;
wire            n368;
wire            n369;
wire            n37;
wire            n371;
wire            n372;
wire            n373;
wire            n374;
wire            n375;
wire            n376;
wire            n378;
wire            n379;
wire            n380;
wire            n381;
wire            n383;
wire            n384;
wire            n385;
wire            n386;
wire            n387;
wire            n388;
wire            n39;
wire            n390;
wire            n392;
wire            n393;
wire            n395;
wire            n396;
wire            n397;
wire            n398;
wire            n399;
wire            n4;
wire            n40;
wire            n400;
wire            n401;
wire            n402;
wire            n404;
wire            n405;
wire            n406;
wire            n407;
wire            n409;
wire            n410;
wire            n412;
wire            n413;
wire            n414;
wire            n415;
wire            n416;
wire            n417;
wire            n419;
wire            n42;
wire            n420;
wire            n421;
wire            n422;
wire            n423;
wire            n425;
wire            n426;
wire            n427;
wire            n428;
wire            n429;
wire            n43;
wire            n430;
wire            n431;
wire            n432;
wire            n433;
wire            n434;
wire      [2:0] n435;
wire      [2:0] n436;
wire      [2:0] n437;
wire      [2:0] n438;
wire      [2:0] n439;
wire      [4:0] n44;
wire      [2:0] n440;
wire      [2:0] n441;
wire            n442;
wire            n443;
wire            n444;
wire            n445;
wire            n446;
wire            n447;
wire            n448;
wire            n449;
wire            n450;
wire            n451;
wire            n452;
wire            n453;
wire            n454;
wire            n455;
wire            n456;
wire            n457;
wire            n458;
wire      [2:0] n459;
wire            n46;
wire      [2:0] n460;
wire      [2:0] n461;
wire            n462;
wire            n463;
wire            n464;
wire      [2:0] n465;
wire            n466;
wire            n467;
wire            n468;
wire            n469;
wire            n470;
wire            n471;
wire            n472;
wire            n473;
wire            n474;
wire            n475;
wire            n476;
wire            n477;
wire            n478;
wire            n479;
wire            n48;
wire            n480;
wire            n481;
wire            n482;
wire            n483;
wire            n484;
wire            n485;
wire            n486;
wire            n487;
wire            n488;
wire            n489;
wire            n49;
wire            n491;
wire            n492;
wire            n493;
wire            n494;
wire            n495;
wire            n496;
wire            n497;
wire            n498;
wire            n499;
wire            n5;
wire      [4:0] n50;
wire      [2:0] n500;
wire      [2:0] n501;
wire      [2:0] n502;
wire      [2:0] n503;
wire      [2:0] n504;
wire      [2:0] n505;
wire            n506;
wire            n507;
wire            n508;
wire            n509;
wire            n510;
wire            n511;
wire      [2:0] n512;
wire      [2:0] n513;
wire            n514;
wire            n515;
wire            n516;
wire            n517;
wire            n518;
wire            n519;
wire            n52;
wire            n520;
wire            n521;
wire            n522;
wire            n523;
wire            n524;
wire            n525;
wire            n526;
wire            n527;
wire            n528;
wire            n529;
wire            n53;
wire            n530;
wire            n531;
wire            n532;
wire            n533;
wire            n534;
wire            n535;
wire            n536;
wire            n537;
wire            n538;
wire            n539;
wire      [6:0] n54;
wire            n540;
wire            n541;
wire            n542;
wire            n543;
wire            n544;
wire            n545;
wire            n546;
wire            n547;
wire            n548;
wire            n549;
wire            n551;
wire            n552;
wire            n554;
wire            n555;
wire            n557;
wire            n558;
wire            n56;
wire            n560;
wire            n561;
wire            n562;
wire            n563;
wire            n565;
wire            n566;
wire            n567;
wire            n568;
wire            n569;
wire            n57;
wire            n570;
wire            n571;
wire            n572;
wire            n573;
wire            n574;
wire            n576;
wire            n577;
wire            n579;
wire            n580;
wire            n582;
wire            n583;
wire            n585;
wire            n586;
wire            n587;
wire            n588;
wire            n59;
wire            n590;
wire            n591;
wire            n593;
wire            n594;
wire            n595;
wire            n596;
wire            n597;
wire            n598;
wire            n599;
wire            n60;
wire            n600;
wire            n601;
wire            n602;
wire            n603;
wire            n604;
wire            n605;
wire            n606;
wire            n607;
wire            n608;
wire            n609;
wire            n610;
wire            n611;
wire            n612;
wire            n613;
wire            n614;
wire            n615;
wire            n616;
wire            n617;
wire            n618;
wire            n619;
wire            n62;
wire            n620;
wire            n621;
wire            n622;
wire            n623;
wire            n624;
wire            n625;
wire            n626;
wire            n627;
wire            n628;
wire            n629;
wire            n63;
wire            n630;
wire            n631;
wire            n632;
wire            n633;
wire            n634;
wire            n635;
wire            n636;
wire            n637;
wire            n638;
wire            n639;
wire            n640;
wire            n641;
wire            n642;
wire            n643;
wire            n644;
wire            n645;
wire            n646;
wire            n647;
wire            n648;
wire            n649;
wire            n65;
wire            n650;
wire            n651;
wire            n652;
wire            n653;
wire            n654;
wire            n655;
wire            n656;
wire            n657;
wire            n658;
wire            n659;
wire            n66;
wire            n660;
wire            n661;
wire            n662;
wire            n663;
wire            n664;
wire            n665;
wire            n666;
wire            n668;
wire            n669;
wire            n671;
wire            n672;
wire            n673;
wire            n674;
wire            n676;
wire            n677;
wire            n679;
wire            n68;
wire            n680;
wire            n682;
wire            n683;
wire            n684;
wire            n685;
wire            n686;
wire            n688;
wire            n689;
wire            n69;
wire            n690;
wire            n691;
wire            n692;
wire            n693;
wire      [2:0] n694;
wire      [2:0] n695;
wire      [2:0] n696;
wire      [2:0] n697;
wire      [2:0] n698;
wire            n699;
wire            n7;
wire            n700;
wire            n701;
wire            n702;
wire            n703;
wire            n704;
wire            n705;
wire            n706;
wire            n707;
wire            n708;
wire      [2:0] n709;
wire            n71;
wire      [2:0] n710;
wire            n711;
wire            n712;
wire            n713;
wire            n714;
wire            n715;
wire            n716;
wire            n717;
wire      [2:0] n718;
wire      [2:0] n719;
wire            n72;
wire      [2:0] n720;
wire      [1:0] n721;
wire            n722;
wire            n723;
wire            n724;
wire            n725;
wire            n726;
wire            n727;
wire            n728;
wire            n729;
wire            n730;
wire            n731;
wire            n732;
wire            n733;
wire            n734;
wire            n735;
wire            n736;
wire            n737;
wire            n738;
wire            n739;
wire            n74;
wire            n740;
wire            n741;
wire            n742;
wire            n743;
wire            n744;
wire            n745;
wire            n746;
wire            n747;
wire            n748;
wire            n749;
wire            n75;
wire            n750;
wire            n751;
wire            n752;
wire            n753;
wire            n754;
wire            n755;
wire            n756;
wire            n757;
wire            n758;
wire            n759;
wire            n760;
wire            n761;
wire            n762;
wire            n763;
wire            n764;
wire            n765;
wire            n766;
wire            n767;
wire            n768;
wire            n769;
wire            n77;
wire            n770;
wire            n771;
wire            n772;
wire            n773;
wire            n774;
wire            n775;
wire            n776;
wire            n777;
wire            n778;
wire            n779;
wire            n78;
wire            n780;
wire            n781;
wire            n782;
wire            n783;
wire            n784;
wire            n785;
wire            n786;
wire            n787;
wire            n788;
wire      [1:0] n789;
wire      [1:0] n790;
wire      [1:0] n791;
wire            n792;
wire            n793;
wire            n795;
wire            n796;
wire            n797;
wire            n798;
wire            n799;
wire            n8;
wire            n80;
wire            n800;
wire            n801;
wire            n802;
wire            n803;
wire            n804;
wire            n805;
wire            n806;
wire            n807;
wire            n808;
wire            n809;
wire            n81;
wire            n810;
wire            n811;
wire            n812;
wire            n813;
wire            n814;
wire            n816;
wire            n817;
wire            n818;
wire            n819;
wire            n820;
wire            n821;
wire            n822;
wire      [3:0] n824;
wire            n825;
wire            n827;
wire      [3:0] n829;
wire            n83;
wire      [3:0] n830;
wire            n831;
wire            n832;
wire            n833;
wire            n834;
wire            n835;
wire            n836;
wire            n837;
wire            n838;
wire            n839;
wire            n84;
wire            n840;
wire            n841;
wire            n842;
wire            n843;
wire            n844;
wire            n845;
wire            n846;
wire            n847;
wire            n849;
wire            n851;
wire            n853;
wire            n854;
wire            n855;
wire            n856;
wire            n857;
wire            n858;
wire            n859;
wire            n86;
wire            n860;
wire            n861;
wire            n862;
wire            n863;
wire            n864;
wire            n865;
wire            n867;
wire            n868;
wire            n869;
wire            n87;
wire            n870;
wire            n871;
wire            n872;
wire            n873;
wire            n874;
wire            n875;
wire            n876;
wire            n877;
wire            n878;
wire            n879;
wire            n881;
wire            n882;
wire            n883;
wire            n884;
wire            n885;
wire            n887;
wire            n888;
wire            n889;
wire            n89;
wire            n890;
wire            n891;
wire            n892;
wire            n893;
wire            n895;
wire            n896;
wire            n897;
wire            n898;
wire            n899;
wire            n90;
wire            n900;
wire            n901;
wire            n902;
wire            n903;
wire            n904;
wire            n905;
wire            n907;
wire            n909;
wire            n910;
wire            n911;
wire            n912;
wire            n914;
wire            n915;
wire            n916;
wire            n917;
wire            n918;
wire            n919;
wire            n92;
wire            n920;
wire            n921;
wire            n922;
wire            n923;
wire            n924;
wire            n925;
wire            n926;
wire            n927;
wire            n928;
wire            n929;
wire            n93;
wire            n930;
wire            n931;
wire            n932;
wire            n934;
wire            n935;
wire            n936;
wire            n937;
wire            n938;
wire            n939;
wire            n940;
wire            n941;
wire            n942;
wire            n943;
wire            n944;
wire            n945;
wire            n946;
wire            n947;
wire            n948;
wire            n949;
wire            n95;
wire            n950;
wire            n951;
wire            n952;
wire            n953;
wire            n954;
wire            n955;
wire            n956;
wire            n958;
wire            n959;
wire            n96;
wire            n960;
wire            n962;
wire            n963;
wire            n964;
wire      [3:0] n966;
wire      [3:0] n967;
wire      [3:0] n968;
wire      [3:0] n969;
wire      [3:0] n970;
wire      [3:0] n971;
wire      [3:0] n972;
wire      [3:0] n973;
wire      [3:0] n974;
wire      [3:0] n975;
wire      [3:0] n976;
wire      [3:0] n977;
wire      [3:0] n978;
wire      [3:0] n979;
wire            n98;
wire      [3:0] n980;
wire            n981;
wire            n982;
wire      [3:0] n983;
wire      [3:0] n984;
wire            n985;
wire            n986;
wire      [3:0] n987;
wire      [3:0] n988;
wire      [1:0] n989;
wire            n99;
wire            n990;
wire            n991;
wire            n992;
wire            n993;
wire            n994;
wire            n995;
wire            n996;
wire            n997;
wire            n998;
wire            n999;
wire      [7:0] op_in;
wire            rst;
wire            wait_data;
assign __ILA_DECODER_valid__ = 1'b1 ;
assign n0 =  ( mem_wait ) == ( 1'b1 )  ;
assign n1 =  ( wait_data ) == ( 1'b1 )  ;
assign n2 =  ( n0 ) | ( n1 )  ;
assign __ILA_DECODER_decode_of_stall__ = n2 ;
assign __ILA_DECODER_acc_decode__[0] = __ILA_DECODER_decode_of_stall__ ;
assign n3 =  ( mem_wait ) == ( 1'b0 )  ;
assign n4 =  ( wait_data ) == ( 1'b0 )  ;
assign n5 =  ( n3 ) & (n4 )  ;
assign bv_2_3_n6 = 2'h3 ;
assign n7 =  ( state ) == ( bv_2_3_n6 )  ;
assign n8 =  ( n5 ) & (n7 )  ;
assign __ILA_DECODER_decode_of_process__ = n8 ;
assign __ILA_DECODER_acc_decode__[1] = __ILA_DECODER_decode_of_process__ ;
assign bv_2_0_n9 = 2'h0 ;
assign n10 =  ( state ) == ( bv_2_0_n9 )  ;
assign n11 =  ( mem_wait ) == ( 1'b0 )  ;
assign n12 =  ( n10 ) & (n11 )  ;
assign n13 =  ( wait_data ) == ( 1'b0 )  ;
assign n14 =  ( n12 ) & (n13 )  ;
assign __ILA_DECODER_decode_of_step_0__ = n14 ;
assign __ILA_DECODER_acc_decode__[2] = __ILA_DECODER_decode_of_step_0__ ;
assign bv_2_1_n15 = 2'h1 ;
assign n16 =  ( state ) == ( bv_2_1_n15 )  ;
assign n17 =  ( mem_wait ) == ( 1'b0 )  ;
assign n18 =  ( n16 ) & (n17 )  ;
assign n19 =  ( wait_data ) == ( 1'b0 )  ;
assign n20 =  ( n18 ) & (n19 )  ;
assign __ILA_DECODER_decode_of_step_1__ = n20 ;
assign __ILA_DECODER_acc_decode__[3] = __ILA_DECODER_decode_of_step_1__ ;
assign bv_2_2_n21 = 2'h2 ;
assign n22 =  ( state ) == ( bv_2_2_n21 )  ;
assign n23 =  ( mem_wait ) == ( 1'b0 )  ;
assign n24 =  ( n22 ) & (n23 )  ;
assign n25 =  ( wait_data ) == ( 1'b0 )  ;
assign n26 =  ( n24 ) & (n25 )  ;
assign __ILA_DECODER_decode_of_step_2__ = n26 ;
assign __ILA_DECODER_acc_decode__[4] = __ILA_DECODER_decode_of_step_2__ ;
assign bv_8_147_n27 = 8'h93 ;
assign n28 =  ( op_in ) == ( bv_8_147_n27 )  ;
assign bv_8_131_n29 = 8'h83 ;
assign n30 =  ( op_in ) == ( bv_8_131_n29 )  ;
assign n31 =  ( n28 ) | ( n30 )  ;
assign bv_8_34_n32 = 8'h22 ;
assign n33 =  ( op_in ) == ( bv_8_34_n32 )  ;
assign n34 =  ( n31 ) | ( n33 )  ;
assign bv_8_50_n35 = 8'h32 ;
assign n36 =  ( op_in ) == ( bv_8_50_n35 )  ;
assign n37 =  ( n34 ) | ( n36 )  ;
assign bv_8_132_n38 = 8'h84 ;
assign n39 =  ( op_in ) == ( bv_8_132_n38 )  ;
assign n40 =  ( n37 ) | ( n39 )  ;
assign bv_8_164_n41 = 8'ha4 ;
assign n42 =  ( op_in ) == ( bv_8_164_n41 )  ;
assign n43 =  ( n40 ) | ( n42 )  ;
assign n44 = op_in[4:0] ;
assign bv_5_17_n45 = 5'h11 ;
assign n46 =  ( n44 ) == ( bv_5_17_n45 )  ;
assign bv_5_1_n47 = 5'h1 ;
assign n48 =  ( n44 ) == ( bv_5_1_n47 )  ;
assign n49 =  ( n46 ) | ( n48 )  ;
assign n50 = op_in[7:3] ;
assign bv_5_23_n51 = 5'h17 ;
assign n52 =  ( n50 ) == ( bv_5_23_n51 )  ;
assign n53 =  ( n49 ) | ( n52 )  ;
assign n54 = op_in[7:1] ;
assign bv_7_91_n55 = 7'h5b ;
assign n56 =  ( n54 ) == ( bv_7_91_n55 )  ;
assign n57 =  ( n53 ) | ( n56 )  ;
assign bv_8_181_n58 = 8'hb5 ;
assign n59 =  ( op_in ) == ( bv_8_181_n58 )  ;
assign n60 =  ( n57 ) | ( n59 )  ;
assign bv_8_180_n61 = 8'hb4 ;
assign n62 =  ( op_in ) == ( bv_8_180_n61 )  ;
assign n63 =  ( n60 ) | ( n62 )  ;
assign bv_8_2_n64 = 8'h2 ;
assign n65 =  ( op_in ) == ( bv_8_2_n64 )  ;
assign n66 =  ( n63 ) | ( n65 )  ;
assign bv_5_27_n67 = 5'h1b ;
assign n68 =  ( n50 ) == ( bv_5_27_n67 )  ;
assign n69 =  ( n66 ) | ( n68 )  ;
assign bv_8_213_n70 = 8'hd5 ;
assign n71 =  ( op_in ) == ( bv_8_213_n70 )  ;
assign n72 =  ( n69 ) | ( n71 )  ;
assign bv_8_18_n73 = 8'h12 ;
assign n74 =  ( op_in ) == ( bv_8_18_n73 )  ;
assign n75 =  ( n72 ) | ( n74 )  ;
assign bv_7_113_n76 = 7'h71 ;
assign n77 =  ( n54 ) == ( bv_7_113_n76 )  ;
assign n78 =  ( n75 ) | ( n77 )  ;
assign bv_7_121_n79 = 7'h79 ;
assign n80 =  ( n54 ) == ( bv_7_121_n79 )  ;
assign n81 =  ( n78 ) | ( n80 )  ;
assign bv_8_224_n82 = 8'he0 ;
assign n83 =  ( op_in ) == ( bv_8_224_n82 )  ;
assign n84 =  ( n81 ) | ( n83 )  ;
assign bv_8_240_n85 = 8'hf0 ;
assign n86 =  ( op_in ) == ( bv_8_240_n85 )  ;
assign n87 =  ( n84 ) | ( n86 )  ;
assign bv_8_128_n88 = 8'h80 ;
assign n89 =  ( op_in ) == ( bv_8_128_n88 )  ;
assign n90 =  ( n87 ) | ( n89 )  ;
assign bv_8_32_n91 = 8'h20 ;
assign n92 =  ( op_in ) == ( bv_8_32_n91 )  ;
assign n93 =  ( n90 ) | ( n92 )  ;
assign bv_8_16_n94 = 8'h10 ;
assign n95 =  ( op_in ) == ( bv_8_16_n94 )  ;
assign n96 =  ( n93 ) | ( n95 )  ;
assign bv_8_64_n97 = 8'h40 ;
assign n98 =  ( op_in ) == ( bv_8_64_n97 )  ;
assign n99 =  ( n96 ) | ( n98 )  ;
assign bv_8_115_n100 = 8'h73 ;
assign n101 =  ( op_in ) == ( bv_8_115_n100 )  ;
assign n102 =  ( n99 ) | ( n101 )  ;
assign bv_8_80_n103 = 8'h50 ;
assign n104 =  ( op_in ) == ( bv_8_80_n103 )  ;
assign n105 =  ( n102 ) | ( n104 )  ;
assign bv_8_48_n106 = 8'h30 ;
assign n107 =  ( op_in ) == ( bv_8_48_n106 )  ;
assign n108 =  ( n105 ) | ( n107 )  ;
assign bv_8_112_n109 = 8'h70 ;
assign n110 =  ( op_in ) == ( bv_8_112_n109 )  ;
assign n111 =  ( n108 ) | ( n110 )  ;
assign bv_8_96_n112 = 8'h60 ;
assign n113 =  ( op_in ) == ( bv_8_96_n112 )  ;
assign n114 =  ( n111 ) | ( n113 )  ;
assign n115 =  ( n114 ) ? ( bv_2_2_n21 ) : ( bv_2_0_n9 ) ;
assign n116 =  ( n43 ) ? ( bv_2_3_n6 ) : ( n115 ) ;
assign n117 =  ( state ) == ( bv_2_0_n9 )  ;
assign n118 =  ( n117 ) ? ( op_in ) : ( op ) ;
assign bv_3_7_n119 = 3'h7 ;
assign n120 =  ( mem_wait ) == ( 1'b1 )  ;
assign bv_3_3_n121 = 3'h3 ;
assign bv_3_1_n122 = 3'h1 ;
assign bv_3_2_n123 = 3'h2 ;
assign bv_3_0_n124 = 3'h0 ;
assign bv_3_4_n125 = 3'h4 ;
assign n126 =  ( n30 ) ? ( bv_3_4_n125 ) : ( bv_3_7_n119 ) ;
assign n127 =  ( n28 ) ? ( bv_3_4_n125 ) : ( n126 ) ;
assign n128 =  ( n83 ) ? ( bv_3_0_n124 ) : ( n127 ) ;
assign n129 =  ( n77 ) ? ( bv_3_2_n123 ) : ( n128 ) ;
assign n130 =  ( n86 ) ? ( bv_3_1_n122 ) : ( n129 ) ;
assign n131 =  ( n80 ) ? ( bv_3_3_n121 ) : ( n130 ) ;
assign n132 =  ( n120 ) ? ( bv_3_7_n119 ) : ( n131 ) ;
assign n133 =  ( wait_data ) ? ( ram_wr_sel ) : ( bv_3_0_n124 ) ;
assign n134 =  ( n46 ) | ( n74 )  ;
assign bv_8_192_n135 = 8'hc0 ;
assign n136 =  ( op_in ) == ( bv_8_192_n135 )  ;
assign n137 =  ( n134 ) | ( n136 )  ;
assign bv_5_3_n138 = 5'h3 ;
assign n139 =  ( n50 ) == ( bv_5_3_n138 )  ;
assign n140 =  ( n139 ) | ( n68 )  ;
assign n141 =  ( n50 ) == ( bv_5_1_n47 )  ;
assign n142 =  ( n140 ) | ( n141 )  ;
assign bv_5_31_n143 = 5'h1f ;
assign n144 =  ( n50 ) == ( bv_5_31_n143 )  ;
assign n145 =  ( n142 ) | ( n144 )  ;
assign bv_5_21_n146 = 5'h15 ;
assign n147 =  ( n50 ) == ( bv_5_21_n146 )  ;
assign n148 =  ( n145 ) | ( n147 )  ;
assign bv_5_15_n149 = 5'hf ;
assign n150 =  ( n50 ) == ( bv_5_15_n149 )  ;
assign n151 =  ( n148 ) | ( n150 )  ;
assign bv_5_25_n152 = 5'h19 ;
assign n153 =  ( n50 ) == ( bv_5_25_n152 )  ;
assign n154 =  ( n151 ) | ( n153 )  ;
assign n155 =  ( n50 ) == ( bv_5_17_n45 )  ;
assign bv_7_67_n156 = 7'h43 ;
assign n157 =  ( n54 ) == ( bv_7_67_n156 )  ;
assign n158 =  ( n155 ) | ( n157 )  ;
assign bv_8_82_n159 = 8'h52 ;
assign n160 =  ( op_in ) == ( bv_8_82_n159 )  ;
assign n161 =  ( n158 ) | ( n160 )  ;
assign bv_8_83_n162 = 8'h53 ;
assign n163 =  ( op_in ) == ( bv_8_83_n162 )  ;
assign n164 =  ( n161 ) | ( n163 )  ;
assign bv_8_194_n165 = 8'hc2 ;
assign n166 =  ( op_in ) == ( bv_8_194_n165 )  ;
assign n167 =  ( n164 ) | ( n166 )  ;
assign bv_8_178_n168 = 8'hb2 ;
assign n169 =  ( op_in ) == ( bv_8_178_n168 )  ;
assign n170 =  ( n167 ) | ( n169 )  ;
assign bv_8_21_n171 = 8'h15 ;
assign n172 =  ( op_in ) == ( bv_8_21_n171 )  ;
assign n173 =  ( n170 ) | ( n172 )  ;
assign n174 =  ( n173 ) | ( n71 )  ;
assign bv_8_5_n175 = 8'h5 ;
assign n176 =  ( op_in ) == ( bv_8_5_n175 )  ;
assign n177 =  ( n174 ) | ( n176 )  ;
assign bv_8_245_n178 = 8'hf5 ;
assign n179 =  ( op_in ) == ( bv_8_245_n178 )  ;
assign n180 =  ( n177 ) | ( n179 )  ;
assign bv_8_117_n181 = 8'h75 ;
assign n182 =  ( op_in ) == ( bv_8_117_n181 )  ;
assign n183 =  ( n180 ) | ( n182 )  ;
assign bv_8_146_n184 = 8'h92 ;
assign n185 =  ( op_in ) == ( bv_8_146_n184 )  ;
assign n186 =  ( n183 ) | ( n185 )  ;
assign bv_8_66_n187 = 8'h42 ;
assign n188 =  ( op_in ) == ( bv_8_66_n187 )  ;
assign n189 =  ( n186 ) | ( n188 )  ;
assign bv_8_67_n190 = 8'h43 ;
assign n191 =  ( op_in ) == ( bv_8_67_n190 )  ;
assign n192 =  ( n189 ) | ( n191 )  ;
assign bv_8_208_n193 = 8'hd0 ;
assign n194 =  ( op_in ) == ( bv_8_208_n193 )  ;
assign n195 =  ( n192 ) | ( n194 )  ;
assign bv_8_210_n196 = 8'hd2 ;
assign n197 =  ( op_in ) == ( bv_8_210_n196 )  ;
assign n198 =  ( n195 ) | ( n197 )  ;
assign bv_8_197_n199 = 8'hc5 ;
assign n200 =  ( op_in ) == ( bv_8_197_n199 )  ;
assign n201 =  ( n198 ) | ( n200 )  ;
assign bv_8_98_n202 = 8'h62 ;
assign n203 =  ( op_in ) == ( bv_8_98_n202 )  ;
assign n204 =  ( n201 ) | ( n203 )  ;
assign bv_8_99_n205 = 8'h63 ;
assign n206 =  ( op_in ) == ( bv_8_99_n205 )  ;
assign n207 =  ( n204 ) | ( n206 )  ;
assign bv_7_11_n208 = 7'hb ;
assign n209 =  ( n54 ) == ( bv_7_11_n208 )  ;
assign bv_7_3_n210 = 7'h3 ;
assign n211 =  ( n54 ) == ( bv_7_3_n210 )  ;
assign n212 =  ( n209 ) | ( n211 )  ;
assign bv_7_123_n213 = 7'h7b ;
assign n214 =  ( n54 ) == ( bv_7_123_n213 )  ;
assign n215 =  ( n212 ) | ( n214 )  ;
assign bv_7_83_n216 = 7'h53 ;
assign n217 =  ( n54 ) == ( bv_7_83_n216 )  ;
assign n218 =  ( n215 ) | ( n217 )  ;
assign bv_7_59_n219 = 7'h3b ;
assign n220 =  ( n54 ) == ( bv_7_59_n219 )  ;
assign n221 =  ( n218 ) | ( n220 )  ;
assign bv_7_99_n222 = 7'h63 ;
assign n223 =  ( n54 ) == ( bv_7_99_n222 )  ;
assign n224 =  ( n221 ) | ( n223 )  ;
assign bv_7_107_n225 = 7'h6b ;
assign n226 =  ( n54 ) == ( bv_7_107_n225 )  ;
assign n227 =  ( n224 ) | ( n226 )  ;
assign bv_8_133_n228 = 8'h85 ;
assign n229 =  ( op_in ) == ( bv_8_133_n228 )  ;
assign bv_3_5_n230 = 3'h5 ;
assign n231 =  ( n229 ) ? ( bv_3_5_n230 ) : ( bv_3_0_n124 ) ;
assign n232 =  ( n227 ) ? ( bv_3_2_n123 ) : ( n231 ) ;
assign n233 =  ( n207 ) ? ( bv_3_1_n122 ) : ( n232 ) ;
assign n234 =  ( n154 ) ? ( bv_3_0_n124 ) : ( n233 ) ;
assign n235 =  ( n137 ) ? ( bv_3_3_n121 ) : ( n234 ) ;
assign n236 =  ( op ) == ( bv_8_132_n38 )  ;
assign n237 =  ( op ) == ( bv_8_164_n41 )  ;
assign n238 =  ( n236 ) | ( n237 )  ;
assign n239 =  ( n238 ) ? ( bv_3_7_n119 ) : ( bv_3_0_n124 ) ;
assign n240 = op[4:0] ;
assign n241 =  ( n240 ) == ( bv_5_17_n45 )  ;
assign n242 =  ( op ) == ( bv_8_18_n73 )  ;
assign n243 =  ( n241 ) | ( n242 )  ;
assign n244 =  ( op ) == ( bv_8_16_n94 )  ;
assign n245 =  ( n244 ) ? ( bv_3_1_n122 ) : ( bv_3_0_n124 ) ;
assign n246 =  ( n243 ) ? ( bv_3_3_n121 ) : ( n245 ) ;
assign bv_8_0_n247 = 8'h0 ;
assign n248 =  ( state ) == ( bv_2_0_n9 )  ;
assign n249 = ~ ( wait_data )  ;
assign n250 =  ( n248 ) & (n249 )  ;
assign n251 =  ( n250 ) ? ( op_in ) : ( op ) ;
assign n252 =  ( mem_wait ) ? ( bv_8_0_n247 ) : ( n251 ) ;
assign n253 = n252[4:0] ;
assign n254 =  ( n253 ) == ( bv_5_17_n45 )  ;
assign n255 =  ( n253 ) == ( bv_5_1_n47 )  ;
assign n256 =  ( n254 ) | ( n255 )  ;
assign n257 = n252[7:1] ;
assign n258 =  ( n257 ) == ( bv_7_113_n76 )  ;
assign n259 =  ( n256 ) | ( n258 )  ;
assign n260 =  ( n257 ) == ( bv_7_121_n79 )  ;
assign n261 =  ( n259 ) | ( n260 )  ;
assign bv_8_84_n262 = 8'h54 ;
assign n263 =  ( n252 ) == ( bv_8_84_n262 )  ;
assign n264 =  ( n261 ) | ( n263 )  ;
assign n265 =  ( n252 ) == ( bv_8_180_n61 )  ;
assign n266 =  ( n264 ) | ( n265 )  ;
assign n267 =  ( n252 ) == ( bv_8_18_n73 )  ;
assign n268 =  ( n266 ) | ( n267 )  ;
assign n269 =  ( n252 ) == ( bv_8_2_n64 )  ;
assign n270 =  ( n268 ) | ( n269 )  ;
assign n271 =  ( n252 ) == ( bv_8_131_n29 )  ;
assign n272 =  ( n270 ) | ( n271 )  ;
assign n273 =  ( n252 ) == ( bv_8_224_n82 )  ;
assign n274 =  ( n272 ) | ( n273 )  ;
assign n275 =  ( n252 ) == ( bv_8_240_n85 )  ;
assign n276 =  ( n274 ) | ( n275 )  ;
assign n277 = n252[7:3] ;
assign bv_5_5_n278 = 5'h5 ;
assign n279 =  ( n277 ) == ( bv_5_5_n278 )  ;
assign bv_5_7_n280 = 5'h7 ;
assign n281 =  ( n277 ) == ( bv_5_7_n280 )  ;
assign n282 =  ( n279 ) | ( n281 )  ;
assign bv_5_11_n283 = 5'hb ;
assign n284 =  ( n277 ) == ( bv_5_11_n283 )  ;
assign n285 =  ( n282 ) | ( n284 )  ;
assign n286 =  ( n277 ) == ( bv_5_23_n51 )  ;
assign n287 =  ( n285 ) | ( n286 )  ;
assign n288 =  ( n277 ) == ( bv_5_3_n138 )  ;
assign n289 =  ( n287 ) | ( n288 )  ;
assign n290 =  ( n277 ) == ( bv_5_27_n67 )  ;
assign n291 =  ( n289 ) | ( n290 )  ;
assign n292 =  ( n277 ) == ( bv_5_1_n47 )  ;
assign n293 =  ( n291 ) | ( n292 )  ;
assign bv_5_29_n294 = 5'h1d ;
assign n295 =  ( n277 ) == ( bv_5_29_n294 )  ;
assign n296 =  ( n293 ) | ( n295 )  ;
assign n297 =  ( n277 ) == ( bv_5_17_n45 )  ;
assign n298 =  ( n296 ) | ( n297 )  ;
assign bv_5_9_n299 = 5'h9 ;
assign n300 =  ( n277 ) == ( bv_5_9_n299 )  ;
assign n301 =  ( n298 ) | ( n300 )  ;
assign bv_5_19_n302 = 5'h13 ;
assign n303 =  ( n277 ) == ( bv_5_19_n302 )  ;
assign n304 =  ( n301 ) | ( n303 )  ;
assign n305 =  ( n277 ) == ( bv_5_25_n152 )  ;
assign n306 =  ( n304 ) | ( n305 )  ;
assign bv_5_13_n307 = 5'hd ;
assign n308 =  ( n277 ) == ( bv_5_13_n307 )  ;
assign n309 =  ( n306 ) | ( n308 )  ;
assign n310 =  ( n277 ) == ( bv_5_21_n146 )  ;
assign n311 =  ( n257 ) == ( bv_7_83_n216 )  ;
assign n312 =  ( n310 ) | ( n311 )  ;
assign bv_8_37_n313 = 8'h25 ;
assign n314 =  ( n252 ) == ( bv_8_37_n313 )  ;
assign n315 =  ( n312 ) | ( n314 )  ;
assign bv_8_53_n316 = 8'h35 ;
assign n317 =  ( n252 ) == ( bv_8_53_n316 )  ;
assign n318 =  ( n315 ) | ( n317 )  ;
assign bv_8_85_n319 = 8'h55 ;
assign n320 =  ( n252 ) == ( bv_8_85_n319 )  ;
assign n321 =  ( n318 ) | ( n320 )  ;
assign n322 =  ( n252 ) == ( bv_8_82_n159 )  ;
assign n323 =  ( n321 ) | ( n322 )  ;
assign n324 =  ( n252 ) == ( bv_8_83_n162 )  ;
assign n325 =  ( n323 ) | ( n324 )  ;
assign bv_8_130_n326 = 8'h82 ;
assign n327 =  ( n252 ) == ( bv_8_130_n326 )  ;
assign n328 =  ( n325 ) | ( n327 )  ;
assign bv_8_176_n329 = 8'hb0 ;
assign n330 =  ( n252 ) == ( bv_8_176_n329 )  ;
assign n331 =  ( n328 ) | ( n330 )  ;
assign n332 =  ( n252 ) == ( bv_8_181_n58 )  ;
assign n333 =  ( n331 ) | ( n332 )  ;
assign n334 =  ( n252 ) == ( bv_8_194_n165 )  ;
assign n335 =  ( n333 ) | ( n334 )  ;
assign n336 =  ( n252 ) == ( bv_8_178_n168 )  ;
assign n337 =  ( n335 ) | ( n336 )  ;
assign n338 =  ( n252 ) == ( bv_8_21_n171 )  ;
assign n339 =  ( n337 ) | ( n338 )  ;
assign n340 =  ( n252 ) == ( bv_8_213_n70 )  ;
assign n341 =  ( n339 ) | ( n340 )  ;
assign n342 =  ( n252 ) == ( bv_8_5_n175 )  ;
assign n343 =  ( n341 ) | ( n342 )  ;
assign n344 =  ( n252 ) == ( bv_8_32_n91 )  ;
assign n345 =  ( n343 ) | ( n344 )  ;
assign n346 =  ( n252 ) == ( bv_8_16_n94 )  ;
assign n347 =  ( n345 ) | ( n346 )  ;
assign n348 =  ( n252 ) == ( bv_8_48_n106 )  ;
assign n349 =  ( n347 ) | ( n348 )  ;
assign bv_8_229_n350 = 8'he5 ;
assign n351 =  ( n252 ) == ( bv_8_229_n350 )  ;
assign n352 =  ( n349 ) | ( n351 )  ;
assign n353 =  ( n252 ) == ( bv_8_133_n228 )  ;
assign n354 =  ( n352 ) | ( n353 )  ;
assign bv_8_162_n355 = 8'ha2 ;
assign n356 =  ( n252 ) == ( bv_8_162_n355 )  ;
assign n357 =  ( n354 ) | ( n356 )  ;
assign n358 =  ( n252 ) == ( bv_8_146_n184 )  ;
assign n359 =  ( n357 ) | ( n358 )  ;
assign bv_8_69_n360 = 8'h45 ;
assign n361 =  ( n252 ) == ( bv_8_69_n360 )  ;
assign n362 =  ( n359 ) | ( n361 )  ;
assign n363 =  ( n252 ) == ( bv_8_66_n187 )  ;
assign n364 =  ( n362 ) | ( n363 )  ;
assign n365 =  ( n252 ) == ( bv_8_67_n190 )  ;
assign n366 =  ( n364 ) | ( n365 )  ;
assign bv_8_114_n367 = 8'h72 ;
assign n368 =  ( n252 ) == ( bv_8_114_n367 )  ;
assign n369 =  ( n366 ) | ( n368 )  ;
assign bv_8_160_n370 = 8'ha0 ;
assign n371 =  ( n252 ) == ( bv_8_160_n370 )  ;
assign n372 =  ( n369 ) | ( n371 )  ;
assign n373 =  ( n252 ) == ( bv_8_192_n135 )  ;
assign n374 =  ( n372 ) | ( n373 )  ;
assign n375 =  ( n252 ) == ( bv_8_210_n196 )  ;
assign n376 =  ( n374 ) | ( n375 )  ;
assign bv_8_149_n377 = 8'h95 ;
assign n378 =  ( n252 ) == ( bv_8_149_n377 )  ;
assign n379 =  ( n376 ) | ( n378 )  ;
assign n380 =  ( n252 ) == ( bv_8_197_n199 )  ;
assign n381 =  ( n379 ) | ( n380 )  ;
assign bv_8_101_n382 = 8'h65 ;
assign n383 =  ( n252 ) == ( bv_8_101_n382 )  ;
assign n384 =  ( n381 ) | ( n383 )  ;
assign n385 =  ( n252 ) == ( bv_8_98_n202 )  ;
assign n386 =  ( n384 ) | ( n385 )  ;
assign n387 =  ( n252 ) == ( bv_8_99_n205 )  ;
assign n388 =  ( n386 ) | ( n387 )  ;
assign bv_7_19_n389 = 7'h13 ;
assign n390 =  ( n257 ) == ( bv_7_19_n389 )  ;
assign bv_7_27_n391 = 7'h1b ;
assign n392 =  ( n257 ) == ( bv_7_27_n391 )  ;
assign n393 =  ( n390 ) | ( n392 )  ;
assign bv_7_43_n394 = 7'h2b ;
assign n395 =  ( n257 ) == ( bv_7_43_n394 )  ;
assign n396 =  ( n393 ) | ( n395 )  ;
assign n397 =  ( n257 ) == ( bv_7_91_n55 )  ;
assign n398 =  ( n396 ) | ( n397 )  ;
assign n399 =  ( n257 ) == ( bv_7_11_n208 )  ;
assign n400 =  ( n398 ) | ( n399 )  ;
assign n401 =  ( n257 ) == ( bv_7_3_n210 )  ;
assign n402 =  ( n400 ) | ( n401 )  ;
assign bv_7_115_n403 = 7'h73 ;
assign n404 =  ( n257 ) == ( bv_7_115_n403 )  ;
assign n405 =  ( n402 ) | ( n404 )  ;
assign n406 =  ( n257 ) == ( bv_7_67_n156 )  ;
assign n407 =  ( n405 ) | ( n406 )  ;
assign bv_7_35_n408 = 7'h23 ;
assign n409 =  ( n257 ) == ( bv_7_35_n408 )  ;
assign n410 =  ( n407 ) | ( n409 )  ;
assign bv_7_75_n411 = 7'h4b ;
assign n412 =  ( n257 ) == ( bv_7_75_n411 )  ;
assign n413 =  ( n410 ) | ( n412 )  ;
assign n414 =  ( n257 ) == ( bv_7_99_n222 )  ;
assign n415 =  ( n413 ) | ( n414 )  ;
assign n416 =  ( n257 ) == ( bv_7_107_n225 )  ;
assign n417 =  ( n415 ) | ( n416 )  ;
assign bv_7_51_n418 = 7'h33 ;
assign n419 =  ( n257 ) == ( bv_7_51_n418 )  ;
assign n420 =  ( n417 ) | ( n419 )  ;
assign n421 =  ( n252 ) == ( bv_8_132_n38 )  ;
assign n422 =  ( n252 ) == ( bv_8_164_n41 )  ;
assign n423 =  ( n421 ) | ( n422 )  ;
assign bv_8_163_n424 = 8'ha3 ;
assign n425 =  ( n252 ) == ( bv_8_163_n424 )  ;
assign n426 =  ( n252 ) == ( bv_8_115_n100 )  ;
assign n427 =  ( n425 ) | ( n426 )  ;
assign n428 =  ( n252 ) == ( bv_8_147_n27 )  ;
assign n429 =  ( n427 ) | ( n428 )  ;
assign n430 =  ( n252 ) == ( bv_8_208_n193 )  ;
assign n431 =  ( n252 ) == ( bv_8_34_n32 )  ;
assign n432 =  ( n430 ) | ( n431 )  ;
assign n433 =  ( n252 ) == ( bv_8_50_n35 )  ;
assign n434 =  ( n432 ) | ( n433 )  ;
assign n435 =  ( n434 ) ? ( bv_3_3_n121 ) : ( bv_3_0_n124 ) ;
assign n436 =  ( n429 ) ? ( bv_3_5_n230 ) : ( n435 ) ;
assign n437 =  ( n423 ) ? ( bv_3_4_n125 ) : ( n436 ) ;
assign n438 =  ( n420 ) ? ( bv_3_1_n122 ) : ( n437 ) ;
assign n439 =  ( n388 ) ? ( bv_3_2_n123 ) : ( n438 ) ;
assign n440 =  ( n309 ) ? ( bv_3_0_n124 ) : ( n439 ) ;
assign n441 =  ( n276 ) ? ( bv_3_0_n124 ) : ( n440 ) ;
assign n442 =  ( n277 ) == ( bv_5_23_n51 )  ;
assign n443 =  ( n257 ) == ( bv_7_91_n55 )  ;
assign n444 =  ( n442 ) | ( n443 )  ;
assign n445 =  ( n252 ) == ( bv_8_181_n58 )  ;
assign n446 =  ( n444 ) | ( n445 )  ;
assign n447 =  ( n252 ) == ( bv_8_180_n61 )  ;
assign n448 =  ( n446 ) | ( n447 )  ;
assign n449 =  ( n277 ) == ( bv_5_27_n67 )  ;
assign n450 =  ( n448 ) | ( n449 )  ;
assign n451 =  ( n252 ) == ( bv_8_213_n70 )  ;
assign n452 =  ( n450 ) | ( n451 )  ;
assign n453 =  ( n252 ) == ( bv_8_34_n32 )  ;
assign n454 =  ( n252 ) == ( bv_8_50_n35 )  ;
assign n455 =  ( n453 ) | ( n454 )  ;
assign n456 =  ( n252 ) == ( bv_8_132_n38 )  ;
assign n457 =  ( n252 ) == ( bv_8_164_n41 )  ;
assign n458 =  ( n456 ) | ( n457 )  ;
assign n459 =  ( n458 ) ? ( bv_3_4_n125 ) : ( bv_3_0_n124 ) ;
assign n460 =  ( n455 ) ? ( bv_3_3_n121 ) : ( n459 ) ;
assign n461 =  ( n452 ) ? ( bv_3_0_n124 ) : ( n460 ) ;
assign n462 =  ( n252 ) == ( bv_8_132_n38 )  ;
assign n463 =  ( n252 ) == ( bv_8_164_n41 )  ;
assign n464 =  ( n462 ) | ( n463 )  ;
assign n465 =  ( n464 ) ? ( bv_3_4_n125 ) : ( bv_3_0_n124 ) ;
assign n466 =  ( n252 ) == ( bv_8_128_n88 )  ;
assign n467 =  ( n252 ) == ( bv_8_34_n32 )  ;
assign n468 =  ( n466 ) | ( n467 )  ;
assign n469 =  ( n252 ) == ( bv_8_50_n35 )  ;
assign n470 =  ( n468 ) | ( n469 )  ;
assign n471 =  ( n277 ) == ( bv_5_23_n51 )  ;
assign n472 =  ( n470 ) | ( n471 )  ;
assign n473 =  ( n257 ) == ( bv_7_91_n55 )  ;
assign n474 =  ( n472 ) | ( n473 )  ;
assign n475 =  ( n252 ) == ( bv_8_181_n58 )  ;
assign n476 =  ( n474 ) | ( n475 )  ;
assign n477 =  ( n252 ) == ( bv_8_180_n61 )  ;
assign n478 =  ( n476 ) | ( n477 )  ;
assign n479 =  ( n277 ) == ( bv_5_27_n67 )  ;
assign n480 =  ( n478 ) | ( n479 )  ;
assign n481 =  ( n252 ) == ( bv_8_213_n70 )  ;
assign n482 =  ( n480 ) | ( n481 )  ;
assign n483 =  ( n252 ) == ( bv_8_115_n100 )  ;
assign n484 =  ( n482 ) | ( n483 )  ;
assign n485 =  ( n252 ) == ( bv_8_48_n106 )  ;
assign n486 =  ( n484 ) | ( n485 )  ;
assign n487 =  ( n252 ) == ( bv_8_64_n97 )  ;
assign n488 =  ( n252 ) == ( bv_8_80_n103 )  ;
assign n489 =  ( n487 ) | ( n488 )  ;
assign bv_3_6_n490 = 3'h6 ;
assign n491 =  ( n252 ) == ( bv_8_112_n109 )  ;
assign n492 =  ( n252 ) == ( bv_8_96_n112 )  ;
assign n493 =  ( n491 ) | ( n492 )  ;
assign n494 =  ( n252 ) == ( bv_8_32_n91 )  ;
assign n495 =  ( n252 ) == ( bv_8_16_n94 )  ;
assign n496 =  ( n494 ) | ( n495 )  ;
assign n497 =  ( n252 ) == ( bv_8_132_n38 )  ;
assign n498 =  ( n252 ) == ( bv_8_164_n41 )  ;
assign n499 =  ( n497 ) | ( n498 )  ;
assign n500 =  ( n499 ) ? ( bv_3_4_n125 ) : ( bv_3_0_n124 ) ;
assign n501 =  ( n496 ) ? ( bv_3_2_n123 ) : ( n500 ) ;
assign n502 =  ( n493 ) ? ( bv_3_7_n119 ) : ( n501 ) ;
assign n503 =  ( n489 ) ? ( bv_3_6_n490 ) : ( n502 ) ;
assign n504 =  ( n486 ) ? ( bv_3_0_n124 ) : ( n503 ) ;
assign n505 =  ( wait_data ) ? ( src_sel1 ) : ( bv_3_0_n124 ) ;
assign n506 =  ( n252 ) == ( bv_8_132_n38 )  ;
assign n507 =  ( n252 ) == ( bv_8_164_n41 )  ;
assign n508 =  ( n506 ) | ( n507 )  ;
assign n509 =  ( n252 ) == ( bv_8_34_n32 )  ;
assign n510 =  ( n252 ) == ( bv_8_50_n35 )  ;
assign n511 =  ( n509 ) | ( n510 )  ;
assign n512 =  ( n511 ) ? ( bv_3_0_n124 ) : ( bv_3_0_n124 ) ;
assign n513 =  ( n508 ) ? ( bv_3_3_n121 ) : ( n512 ) ;
assign n514 =  ( n253 ) == ( bv_5_17_n45 )  ;
assign n515 =  ( n252 ) == ( bv_8_18_n73 )  ;
assign n516 =  ( n514 ) | ( n515 )  ;
assign n517 =  ( n252 ) == ( bv_8_131_n29 )  ;
assign n518 =  ( n516 ) | ( n517 )  ;
assign n519 =  ( n277 ) == ( bv_5_5_n278 )  ;
assign n520 =  ( n277 ) == ( bv_5_7_n280 )  ;
assign n521 =  ( n519 ) | ( n520 )  ;
assign n522 =  ( n277 ) == ( bv_5_11_n283 )  ;
assign n523 =  ( n521 ) | ( n522 )  ;
assign n524 =  ( n277 ) == ( bv_5_31_n143 )  ;
assign n525 =  ( n523 ) | ( n524 )  ;
assign n526 =  ( n277 ) == ( bv_5_19_n302 )  ;
assign n527 =  ( n525 ) | ( n526 )  ;
assign n528 =  ( n257 ) == ( bv_7_19_n389 )  ;
assign n529 =  ( n527 ) | ( n528 )  ;
assign n530 =  ( n257 ) == ( bv_7_27_n391 )  ;
assign n531 =  ( n529 ) | ( n530 )  ;
assign n532 =  ( n257 ) == ( bv_7_43_n394 )  ;
assign n533 =  ( n531 ) | ( n532 )  ;
assign n534 =  ( n257 ) == ( bv_7_123_n213 )  ;
assign n535 =  ( n533 ) | ( n534 )  ;
assign n536 =  ( n257 ) == ( bv_7_75_n411 )  ;
assign n537 =  ( n535 ) | ( n536 )  ;
assign n538 =  ( n252 ) == ( bv_8_37_n313 )  ;
assign n539 =  ( n537 ) | ( n538 )  ;
assign n540 =  ( n252 ) == ( bv_8_53_n316 )  ;
assign n541 =  ( n539 ) | ( n540 )  ;
assign n542 =  ( n252 ) == ( bv_8_85_n319 )  ;
assign n543 =  ( n541 ) | ( n542 )  ;
assign n544 =  ( n252 ) == ( bv_8_82_n159 )  ;
assign n545 =  ( n543 ) | ( n544 )  ;
assign n546 =  ( n252 ) == ( bv_8_181_n58 )  ;
assign n547 =  ( n545 ) | ( n546 )  ;
assign n548 =  ( n252 ) == ( bv_8_180_n61 )  ;
assign n549 =  ( n547 ) | ( n548 )  ;
assign bv_8_228_n550 = 8'he4 ;
assign n551 =  ( n252 ) == ( bv_8_228_n550 )  ;
assign n552 =  ( n549 ) | ( n551 )  ;
assign bv_8_244_n553 = 8'hf4 ;
assign n554 =  ( n252 ) == ( bv_8_244_n553 )  ;
assign n555 =  ( n552 ) | ( n554 )  ;
assign bv_8_212_n556 = 8'hd4 ;
assign n557 =  ( n252 ) == ( bv_8_212_n556 )  ;
assign n558 =  ( n555 ) | ( n557 )  ;
assign bv_8_20_n559 = 8'h14 ;
assign n560 =  ( n252 ) == ( bv_8_20_n559 )  ;
assign n561 =  ( n558 ) | ( n560 )  ;
assign n562 =  ( n252 ) == ( bv_8_132_n38 )  ;
assign n563 =  ( n561 ) | ( n562 )  ;
assign bv_8_4_n564 = 8'h4 ;
assign n565 =  ( n252 ) == ( bv_8_4_n564 )  ;
assign n566 =  ( n563 ) | ( n565 )  ;
assign n567 =  ( n252 ) == ( bv_8_115_n100 )  ;
assign n568 =  ( n566 ) | ( n567 )  ;
assign n569 =  ( n252 ) == ( bv_8_245_n178 )  ;
assign n570 =  ( n568 ) | ( n569 )  ;
assign n571 =  ( n252 ) == ( bv_8_147_n27 )  ;
assign n572 =  ( n570 ) | ( n571 )  ;
assign n573 =  ( n252 ) == ( bv_8_164_n41 )  ;
assign n574 =  ( n572 ) | ( n573 )  ;
assign bv_8_35_n575 = 8'h23 ;
assign n576 =  ( n252 ) == ( bv_8_35_n575 )  ;
assign n577 =  ( n574 ) | ( n576 )  ;
assign bv_8_51_n578 = 8'h33 ;
assign n579 =  ( n252 ) == ( bv_8_51_n578 )  ;
assign n580 =  ( n577 ) | ( n579 )  ;
assign bv_8_3_n581 = 8'h3 ;
assign n582 =  ( n252 ) == ( bv_8_3_n581 )  ;
assign n583 =  ( n580 ) | ( n582 )  ;
assign bv_8_19_n584 = 8'h13 ;
assign n585 =  ( n252 ) == ( bv_8_19_n584 )  ;
assign n586 =  ( n583 ) | ( n585 )  ;
assign n587 =  ( n252 ) == ( bv_8_149_n377 )  ;
assign n588 =  ( n586 ) | ( n587 )  ;
assign bv_8_148_n589 = 8'h94 ;
assign n590 =  ( n252 ) == ( bv_8_148_n589 )  ;
assign n591 =  ( n588 ) | ( n590 )  ;
assign bv_8_196_n592 = 8'hc4 ;
assign n593 =  ( n252 ) == ( bv_8_196_n592 )  ;
assign n594 =  ( n591 ) | ( n593 )  ;
assign n595 =  ( n277 ) == ( bv_5_23_n51 )  ;
assign n596 =  ( n277 ) == ( bv_5_3_n138 )  ;
assign n597 =  ( n595 ) | ( n596 )  ;
assign n598 =  ( n277 ) == ( bv_5_27_n67 )  ;
assign n599 =  ( n597 ) | ( n598 )  ;
assign n600 =  ( n277 ) == ( bv_5_1_n47 )  ;
assign n601 =  ( n599 ) | ( n600 )  ;
assign n602 =  ( n277 ) == ( bv_5_29_n294 )  ;
assign n603 =  ( n601 ) | ( n602 )  ;
assign n604 =  ( n277 ) == ( bv_5_21_n146 )  ;
assign n605 =  ( n603 ) | ( n604 )  ;
assign n606 =  ( n277 ) == ( bv_5_17_n45 )  ;
assign n607 =  ( n605 ) | ( n606 )  ;
assign n608 =  ( n277 ) == ( bv_5_9_n299 )  ;
assign n609 =  ( n607 ) | ( n608 )  ;
assign n610 =  ( n277 ) == ( bv_5_25_n152 )  ;
assign n611 =  ( n609 ) | ( n610 )  ;
assign n612 =  ( n277 ) == ( bv_5_13_n307 )  ;
assign n613 =  ( n611 ) | ( n612 )  ;
assign n614 =  ( n257 ) == ( bv_7_91_n55 )  ;
assign n615 =  ( n613 ) | ( n614 )  ;
assign n616 =  ( n257 ) == ( bv_7_11_n208 )  ;
assign n617 =  ( n615 ) | ( n616 )  ;
assign n618 =  ( n257 ) == ( bv_7_3_n210 )  ;
assign n619 =  ( n617 ) | ( n618 )  ;
assign n620 =  ( n257 ) == ( bv_7_115_n403 )  ;
assign n621 =  ( n619 ) | ( n620 )  ;
assign n622 =  ( n257 ) == ( bv_7_67_n156 )  ;
assign n623 =  ( n621 ) | ( n622 )  ;
assign n624 =  ( n257 ) == ( bv_7_83_n216 )  ;
assign n625 =  ( n623 ) | ( n624 )  ;
assign n626 =  ( n257 ) == ( bv_7_35_n408 )  ;
assign n627 =  ( n625 ) | ( n626 )  ;
assign n628 =  ( n257 ) == ( bv_7_99_n222 )  ;
assign n629 =  ( n627 ) | ( n628 )  ;
assign n630 =  ( n257 ) == ( bv_7_107_n225 )  ;
assign n631 =  ( n629 ) | ( n630 )  ;
assign n632 =  ( n257 ) == ( bv_7_51_n418 )  ;
assign n633 =  ( n631 ) | ( n632 )  ;
assign n634 =  ( n252 ) == ( bv_8_21_n171 )  ;
assign n635 =  ( n633 ) | ( n634 )  ;
assign n636 =  ( n252 ) == ( bv_8_213_n70 )  ;
assign n637 =  ( n635 ) | ( n636 )  ;
assign n638 =  ( n252 ) == ( bv_8_5_n175 )  ;
assign n639 =  ( n637 ) | ( n638 )  ;
assign n640 =  ( n252 ) == ( bv_8_163_n424 )  ;
assign n641 =  ( n639 ) | ( n640 )  ;
assign n642 =  ( n252 ) == ( bv_8_229_n350 )  ;
assign n643 =  ( n641 ) | ( n642 )  ;
assign n644 =  ( n252 ) == ( bv_8_133_n228 )  ;
assign n645 =  ( n643 ) | ( n644 )  ;
assign n646 =  ( n252 ) == ( bv_8_69_n360 )  ;
assign n647 =  ( n645 ) | ( n646 )  ;
assign n648 =  ( n252 ) == ( bv_8_66_n187 )  ;
assign n649 =  ( n647 ) | ( n648 )  ;
assign n650 =  ( n252 ) == ( bv_8_208_n193 )  ;
assign n651 =  ( n649 ) | ( n650 )  ;
assign n652 =  ( n252 ) == ( bv_8_192_n135 )  ;
assign n653 =  ( n651 ) | ( n652 )  ;
assign n654 =  ( n252 ) == ( bv_8_34_n32 )  ;
assign n655 =  ( n653 ) | ( n654 )  ;
assign n656 =  ( n252 ) == ( bv_8_50_n35 )  ;
assign n657 =  ( n655 ) | ( n656 )  ;
assign n658 =  ( n252 ) == ( bv_8_197_n199 )  ;
assign n659 =  ( n657 ) | ( n658 )  ;
assign n660 =  ( n252 ) == ( bv_8_101_n382 )  ;
assign n661 =  ( n659 ) | ( n660 )  ;
assign n662 =  ( n252 ) == ( bv_8_98_n202 )  ;
assign n663 =  ( n661 ) | ( n662 )  ;
assign n664 =  ( n277 ) == ( bv_5_15_n149 )  ;
assign n665 =  ( n257 ) == ( bv_7_59_n219 )  ;
assign n666 =  ( n664 ) | ( n665 )  ;
assign bv_8_36_n667 = 8'h24 ;
assign n668 =  ( n252 ) == ( bv_8_36_n667 )  ;
assign n669 =  ( n666 ) | ( n668 )  ;
assign bv_8_52_n670 = 8'h34 ;
assign n671 =  ( n252 ) == ( bv_8_52_n670 )  ;
assign n672 =  ( n669 ) | ( n671 )  ;
assign n673 =  ( n252 ) == ( bv_8_84_n262 )  ;
assign n674 =  ( n672 ) | ( n673 )  ;
assign bv_8_116_n675 = 8'h74 ;
assign n676 =  ( n252 ) == ( bv_8_116_n675 )  ;
assign n677 =  ( n674 ) | ( n676 )  ;
assign bv_8_68_n678 = 8'h44 ;
assign n679 =  ( n252 ) == ( bv_8_68_n678 )  ;
assign n680 =  ( n677 ) | ( n679 )  ;
assign bv_8_100_n681 = 8'h64 ;
assign n682 =  ( n252 ) == ( bv_8_100_n681 )  ;
assign n683 =  ( n680 ) | ( n682 )  ;
assign n684 =  ( n252 ) == ( bv_8_83_n162 )  ;
assign n685 =  ( n252 ) == ( bv_8_117_n181 )  ;
assign n686 =  ( n684 ) | ( n685 )  ;
assign bv_8_144_n687 = 8'h90 ;
assign n688 =  ( n252 ) == ( bv_8_144_n687 )  ;
assign n689 =  ( n686 ) | ( n688 )  ;
assign n690 =  ( n252 ) == ( bv_8_67_n190 )  ;
assign n691 =  ( n689 ) | ( n690 )  ;
assign n692 =  ( n252 ) == ( bv_8_99_n205 )  ;
assign n693 =  ( n691 ) | ( n692 )  ;
assign n694 =  ( n693 ) ? ( bv_3_2_n123 ) : ( bv_3_0_n124 ) ;
assign n695 =  ( n683 ) ? ( bv_3_1_n122 ) : ( n694 ) ;
assign n696 =  ( n663 ) ? ( bv_3_0_n124 ) : ( n695 ) ;
assign n697 =  ( n594 ) ? ( bv_3_3_n121 ) : ( n696 ) ;
assign n698 =  ( n518 ) ? ( bv_3_5_n230 ) : ( n697 ) ;
assign n699 =  ( n252 ) == ( bv_8_132_n38 )  ;
assign n700 =  ( n252 ) == ( bv_8_164_n41 )  ;
assign n701 =  ( n699 ) | ( n700 )  ;
assign n702 =  ( n252 ) == ( bv_8_147_n27 )  ;
assign n703 =  ( n252 ) == ( bv_8_131_n29 )  ;
assign n704 =  ( n702 ) | ( n703 )  ;
assign n705 =  ( n252 ) == ( bv_8_224_n82 )  ;
assign n706 =  ( n704 ) | ( n705 )  ;
assign n707 =  ( n257 ) == ( bv_7_113_n76 )  ;
assign n708 =  ( n706 ) | ( n707 )  ;
assign n709 =  ( n708 ) ? ( bv_3_7_n119 ) : ( bv_3_0_n124 ) ;
assign n710 =  ( n701 ) ? ( bv_3_3_n121 ) : ( n709 ) ;
assign n711 =  ( n253 ) == ( bv_5_17_n45 )  ;
assign n712 =  ( n252 ) == ( bv_8_18_n73 )  ;
assign n713 =  ( n711 ) | ( n712 )  ;
assign n714 =  ( n252 ) == ( bv_8_132_n38 )  ;
assign n715 =  ( n252 ) == ( bv_8_164_n41 )  ;
assign n716 =  ( n714 ) | ( n715 )  ;
assign n717 =  ( n252 ) == ( bv_8_16_n94 )  ;
assign n718 =  ( n717 ) ? ( bv_3_0_n124 ) : ( bv_3_0_n124 ) ;
assign n719 =  ( n716 ) ? ( bv_3_3_n121 ) : ( n718 ) ;
assign n720 =  ( n713 ) ? ( bv_3_4_n125 ) : ( n719 ) ;
assign n721 =  ( wait_data ) ? ( src_sel2 ) : ( bv_2_0_n9 ) ;
assign n722 =  ( n277 ) == ( bv_5_23_n51 )  ;
assign n723 =  ( n257 ) == ( bv_7_91_n55 )  ;
assign n724 =  ( n722 ) | ( n723 )  ;
assign n725 =  ( n252 ) == ( bv_8_180_n61 )  ;
assign n726 =  ( n724 ) | ( n725 )  ;
assign n727 =  ( n252 ) == ( bv_8_144_n687 )  ;
assign n728 =  ( n726 ) | ( n727 )  ;
assign n729 =  ( n252 ) == ( bv_8_148_n589 )  ;
assign n730 =  ( n728 ) | ( n729 )  ;
assign n731 =  ( n277 ) == ( bv_5_9_n299 )  ;
assign n732 =  ( n277 ) == ( bv_5_25_n152 )  ;
assign n733 =  ( n731 ) | ( n732 )  ;
assign n734 =  ( n277 ) == ( bv_5_13_n307 )  ;
assign n735 =  ( n733 ) | ( n734 )  ;
assign n736 =  ( n257 ) == ( bv_7_35_n408 )  ;
assign n737 =  ( n735 ) | ( n736 )  ;
assign n738 =  ( n257 ) == ( bv_7_99_n222 )  ;
assign n739 =  ( n737 ) | ( n738 )  ;
assign n740 =  ( n257 ) == ( bv_7_107_n225 )  ;
assign n741 =  ( n739 ) | ( n740 )  ;
assign n742 =  ( n257 ) == ( bv_7_51_n418 )  ;
assign n743 =  ( n741 ) | ( n742 )  ;
assign n744 =  ( n252 ) == ( bv_8_36_n667 )  ;
assign n745 =  ( n743 ) | ( n744 )  ;
assign n746 =  ( n252 ) == ( bv_8_52_n670 )  ;
assign n747 =  ( n745 ) | ( n746 )  ;
assign n748 =  ( n252 ) == ( bv_8_84_n262 )  ;
assign n749 =  ( n747 ) | ( n748 )  ;
assign n750 =  ( n252 ) == ( bv_8_228_n550 )  ;
assign n751 =  ( n749 ) | ( n750 )  ;
assign n752 =  ( n252 ) == ( bv_8_131_n29 )  ;
assign n753 =  ( n751 ) | ( n752 )  ;
assign n754 =  ( n252 ) == ( bv_8_69_n360 )  ;
assign n755 =  ( n753 ) | ( n754 )  ;
assign n756 =  ( n252 ) == ( bv_8_68_n678 )  ;
assign n757 =  ( n755 ) | ( n756 )  ;
assign n758 =  ( n252 ) == ( bv_8_66_n187 )  ;
assign n759 =  ( n757 ) | ( n758 )  ;
assign n760 =  ( n252 ) == ( bv_8_197_n199 )  ;
assign n761 =  ( n759 ) | ( n760 )  ;
assign n762 =  ( n252 ) == ( bv_8_101_n382 )  ;
assign n763 =  ( n761 ) | ( n762 )  ;
assign n764 =  ( n252 ) == ( bv_8_100_n681 )  ;
assign n765 =  ( n763 ) | ( n764 )  ;
assign n766 =  ( n252 ) == ( bv_8_98_n202 )  ;
assign n767 =  ( n765 ) | ( n766 )  ;
assign n768 =  ( n277 ) == ( bv_5_3_n138 )  ;
assign n769 =  ( n277 ) == ( bv_5_27_n67 )  ;
assign n770 =  ( n768 ) | ( n769 )  ;
assign n771 =  ( n277 ) == ( bv_5_1_n47 )  ;
assign n772 =  ( n770 ) | ( n771 )  ;
assign n773 =  ( n257 ) == ( bv_7_11_n208 )  ;
assign n774 =  ( n772 ) | ( n773 )  ;
assign n775 =  ( n257 ) == ( bv_7_3_n210 )  ;
assign n776 =  ( n774 ) | ( n775 )  ;
assign n777 =  ( n252 ) == ( bv_8_20_n559 )  ;
assign n778 =  ( n776 ) | ( n777 )  ;
assign n779 =  ( n252 ) == ( bv_8_21_n171 )  ;
assign n780 =  ( n778 ) | ( n779 )  ;
assign n781 =  ( n252 ) == ( bv_8_213_n70 )  ;
assign n782 =  ( n780 ) | ( n781 )  ;
assign n783 =  ( n252 ) == ( bv_8_4_n564 )  ;
assign n784 =  ( n782 ) | ( n783 )  ;
assign n785 =  ( n252 ) == ( bv_8_5_n175 )  ;
assign n786 =  ( n784 ) | ( n785 )  ;
assign n787 =  ( n252 ) == ( bv_8_163_n424 )  ;
assign n788 =  ( n786 ) | ( n787 )  ;
assign n789 =  ( n788 ) ? ( bv_2_2_n21 ) : ( bv_2_0_n9 ) ;
assign n790 =  ( n767 ) ? ( bv_2_1_n15 ) : ( n789 ) ;
assign n791 =  ( n730 ) ? ( bv_2_3_n6 ) : ( n790 ) ;
assign n792 =  ( wait_data ) ? ( src_sel3 ) : ( 1'b0 )  ;
assign n793 =  ( n252 ) == ( bv_8_228_n550 )  ;
assign bv_8_195_n794 = 8'hc3 ;
assign n795 =  ( n252 ) == ( bv_8_195_n794 )  ;
assign n796 =  ( n793 ) | ( n795 )  ;
assign n797 =  ( n252 ) == ( bv_8_194_n165 )  ;
assign n798 =  ( n796 ) | ( n797 )  ;
assign n799 =  ( n252 ) == ( bv_8_32_n91 )  ;
assign n800 =  ( n798 ) | ( n799 )  ;
assign n801 =  ( n252 ) == ( bv_8_16_n94 )  ;
assign n802 =  ( n800 ) | ( n801 )  ;
assign n803 =  ( n252 ) == ( bv_8_64_n97 )  ;
assign n804 =  ( n802 ) | ( n803 )  ;
assign n805 =  ( n252 ) == ( bv_8_48_n106 )  ;
assign n806 =  ( n804 ) | ( n805 )  ;
assign n807 =  ( n252 ) == ( bv_8_80_n103 )  ;
assign n808 =  ( n806 ) | ( n807 )  ;
assign n809 =  ( n252 ) == ( bv_8_112_n109 )  ;
assign n810 =  ( n808 ) | ( n809 )  ;
assign n811 =  ( n252 ) == ( bv_8_96_n112 )  ;
assign n812 =  ( n810 ) | ( n811 )  ;
assign n813 =  ( n252 ) == ( bv_8_131_n29 )  ;
assign n814 =  ( n812 ) | ( n813 )  ;
assign bv_8_211_n815 = 8'hd3 ;
assign n816 =  ( n252 ) == ( bv_8_211_n815 )  ;
assign n817 =  ( n814 ) | ( n816 )  ;
assign n818 =  ( n252 ) == ( bv_8_210_n196 )  ;
assign n819 =  ( n817 ) | ( n818 )  ;
assign n820 =  ( n252 ) == ( bv_8_128_n88 )  ;
assign n821 =  ( n819 ) | ( n820 )  ;
assign n822 =  ( n821 ) ? ( 1'b1 ) : ( 1'b0 )  ;
assign bv_4_0_n823 = 4'h0 ;
assign n824 =  ( wait_data ) ? ( alu_op ) : ( bv_4_0_n823 ) ;
assign n825 =  ( n252 ) == ( bv_8_164_n41 )  ;
assign bv_4_3_n826 = 4'h3 ;
assign n827 =  ( n252 ) == ( bv_8_132_n38 )  ;
assign bv_4_4_n828 = 4'h4 ;
assign n829 =  ( n827 ) ? ( bv_4_4_n828 ) : ( bv_4_0_n823 ) ;
assign n830 =  ( n825 ) ? ( bv_4_3_n826 ) : ( n829 ) ;
assign n831 =  ( n277 ) == ( bv_5_23_n51 )  ;
assign n832 =  ( n277 ) == ( bv_5_19_n302 )  ;
assign n833 =  ( n831 ) | ( n832 )  ;
assign n834 =  ( n257 ) == ( bv_7_91_n55 )  ;
assign n835 =  ( n833 ) | ( n834 )  ;
assign n836 =  ( n257 ) == ( bv_7_75_n411 )  ;
assign n837 =  ( n835 ) | ( n836 )  ;
assign n838 =  ( n252 ) == ( bv_8_181_n58 )  ;
assign n839 =  ( n837 ) | ( n838 )  ;
assign n840 =  ( n252 ) == ( bv_8_180_n61 )  ;
assign n841 =  ( n839 ) | ( n840 )  ;
assign n842 =  ( n252 ) == ( bv_8_228_n550 )  ;
assign n843 =  ( n841 ) | ( n842 )  ;
assign n844 =  ( n252 ) == ( bv_8_149_n377 )  ;
assign n845 =  ( n843 ) | ( n844 )  ;
assign n846 =  ( n252 ) == ( bv_8_148_n589 )  ;
assign n847 =  ( n845 ) | ( n846 )  ;
assign bv_4_2_n848 = 4'h2 ;
assign n849 =  ( n252 ) == ( bv_8_19_n584 )  ;
assign bv_4_13_n850 = 4'hd ;
assign n851 =  ( n252 ) == ( bv_8_212_n556 )  ;
assign bv_4_5_n852 = 4'h5 ;
assign n853 =  ( n277 ) == ( bv_5_11_n283 )  ;
assign n854 =  ( n257 ) == ( bv_7_43_n394 )  ;
assign n855 =  ( n853 ) | ( n854 )  ;
assign n856 =  ( n252 ) == ( bv_8_85_n319 )  ;
assign n857 =  ( n855 ) | ( n856 )  ;
assign n858 =  ( n252 ) == ( bv_8_84_n262 )  ;
assign n859 =  ( n857 ) | ( n858 )  ;
assign n860 =  ( n252 ) == ( bv_8_82_n159 )  ;
assign n861 =  ( n859 ) | ( n860 )  ;
assign n862 =  ( n252 ) == ( bv_8_83_n162 )  ;
assign n863 =  ( n861 ) | ( n862 )  ;
assign n864 =  ( n252 ) == ( bv_8_130_n326 )  ;
assign n865 =  ( n863 ) | ( n864 )  ;
assign bv_4_7_n866 = 4'h7 ;
assign n867 =  ( n277 ) == ( bv_5_9_n299 )  ;
assign n868 =  ( n257 ) == ( bv_7_35_n408 )  ;
assign n869 =  ( n867 ) | ( n868 )  ;
assign n870 =  ( n252 ) == ( bv_8_69_n360 )  ;
assign n871 =  ( n869 ) | ( n870 )  ;
assign n872 =  ( n252 ) == ( bv_8_68_n678 )  ;
assign n873 =  ( n871 ) | ( n872 )  ;
assign n874 =  ( n252 ) == ( bv_8_66_n187 )  ;
assign n875 =  ( n873 ) | ( n874 )  ;
assign n876 =  ( n252 ) == ( bv_8_67_n190 )  ;
assign n877 =  ( n875 ) | ( n876 )  ;
assign n878 =  ( n252 ) == ( bv_8_114_n367 )  ;
assign n879 =  ( n877 ) | ( n878 )  ;
assign bv_4_9_n880 = 4'h9 ;
assign n881 =  ( n252 ) == ( bv_8_164_n41 )  ;
assign n882 =  ( n252 ) == ( bv_8_132_n38 )  ;
assign n883 =  ( n252 ) == ( bv_8_176_n329 )  ;
assign n884 =  ( n252 ) == ( bv_8_3_n581 )  ;
assign n885 =  ( n883 ) | ( n884 )  ;
assign bv_4_12_n886 = 4'hc ;
assign n887 =  ( n277 ) == ( bv_5_25_n152 )  ;
assign n888 =  ( n257 ) == ( bv_7_99_n222 )  ;
assign n889 =  ( n887 ) | ( n888 )  ;
assign n890 =  ( n257 ) == ( bv_7_107_n225 )  ;
assign n891 =  ( n889 ) | ( n890 )  ;
assign n892 =  ( n252 ) == ( bv_8_197_n199 )  ;
assign n893 =  ( n891 ) | ( n892 )  ;
assign bv_4_15_n894 = 4'hf ;
assign n895 =  ( n277 ) == ( bv_5_13_n307 )  ;
assign n896 =  ( n257 ) == ( bv_7_51_n418 )  ;
assign n897 =  ( n895 ) | ( n896 )  ;
assign n898 =  ( n252 ) == ( bv_8_101_n382 )  ;
assign n899 =  ( n897 ) | ( n898 )  ;
assign n900 =  ( n252 ) == ( bv_8_100_n681 )  ;
assign n901 =  ( n899 ) | ( n900 )  ;
assign n902 =  ( n252 ) == ( bv_8_98_n202 )  ;
assign n903 =  ( n901 ) | ( n902 )  ;
assign n904 =  ( n252 ) == ( bv_8_99_n205 )  ;
assign n905 =  ( n903 ) | ( n904 )  ;
assign bv_4_8_n906 = 4'h8 ;
assign n907 =  ( n252 ) == ( bv_8_244_n553 )  ;
assign bv_8_179_n908 = 8'hb3 ;
assign n909 =  ( n252 ) == ( bv_8_179_n908 )  ;
assign n910 =  ( n907 ) | ( n909 )  ;
assign n911 =  ( n252 ) == ( bv_8_178_n168 )  ;
assign n912 =  ( n910 ) | ( n911 )  ;
assign bv_4_6_n913 = 4'h6 ;
assign n914 =  ( n277 ) == ( bv_5_3_n138 )  ;
assign n915 =  ( n277 ) == ( bv_5_27_n67 )  ;
assign n916 =  ( n914 ) | ( n915 )  ;
assign n917 =  ( n277 ) == ( bv_5_1_n47 )  ;
assign n918 =  ( n916 ) | ( n917 )  ;
assign n919 =  ( n257 ) == ( bv_7_11_n208 )  ;
assign n920 =  ( n918 ) | ( n919 )  ;
assign n921 =  ( n257 ) == ( bv_7_3_n210 )  ;
assign n922 =  ( n920 ) | ( n921 )  ;
assign n923 =  ( n252 ) == ( bv_8_20_n559 )  ;
assign n924 =  ( n922 ) | ( n923 )  ;
assign n925 =  ( n252 ) == ( bv_8_21_n171 )  ;
assign n926 =  ( n924 ) | ( n925 )  ;
assign n927 =  ( n252 ) == ( bv_8_213_n70 )  ;
assign n928 =  ( n926 ) | ( n927 )  ;
assign n929 =  ( n252 ) == ( bv_8_4_n564 )  ;
assign n930 =  ( n928 ) | ( n929 )  ;
assign n931 =  ( n252 ) == ( bv_8_5_n175 )  ;
assign n932 =  ( n930 ) | ( n931 )  ;
assign bv_4_14_n933 = 4'he ;
assign n934 =  ( n277 ) == ( bv_5_5_n278 )  ;
assign n935 =  ( n277 ) == ( bv_5_7_n280 )  ;
assign n936 =  ( n934 ) | ( n935 )  ;
assign n937 =  ( n257 ) == ( bv_7_19_n389 )  ;
assign n938 =  ( n936 ) | ( n937 )  ;
assign n939 =  ( n257 ) == ( bv_7_27_n391 )  ;
assign n940 =  ( n938 ) | ( n939 )  ;
assign n941 =  ( n252 ) == ( bv_8_37_n313 )  ;
assign n942 =  ( n940 ) | ( n941 )  ;
assign n943 =  ( n252 ) == ( bv_8_36_n667 )  ;
assign n944 =  ( n942 ) | ( n943 )  ;
assign n945 =  ( n252 ) == ( bv_8_53_n316 )  ;
assign n946 =  ( n944 ) | ( n945 )  ;
assign n947 =  ( n252 ) == ( bv_8_52_n670 )  ;
assign n948 =  ( n946 ) | ( n947 )  ;
assign n949 =  ( n252 ) == ( bv_8_163_n424 )  ;
assign n950 =  ( n948 ) | ( n949 )  ;
assign n951 =  ( n252 ) == ( bv_8_115_n100 )  ;
assign n952 =  ( n950 ) | ( n951 )  ;
assign n953 =  ( n252 ) == ( bv_8_147_n27 )  ;
assign n954 =  ( n952 ) | ( n953 )  ;
assign n955 =  ( n252 ) == ( bv_8_131_n29 )  ;
assign n956 =  ( n954 ) | ( n955 )  ;
assign bv_4_1_n957 = 4'h1 ;
assign n958 =  ( n252 ) == ( bv_8_160_n370 )  ;
assign n959 =  ( n252 ) == ( bv_8_35_n575 )  ;
assign n960 =  ( n958 ) | ( n959 )  ;
assign bv_4_10_n961 = 4'ha ;
assign n962 =  ( n252 ) == ( bv_8_51_n578 )  ;
assign n963 =  ( n252 ) == ( bv_8_196_n592 )  ;
assign n964 =  ( n962 ) | ( n963 )  ;
assign bv_4_11_n965 = 4'hb ;
assign n966 =  ( n964 ) ? ( bv_4_11_n965 ) : ( bv_4_0_n823 ) ;
assign n967 =  ( n960 ) ? ( bv_4_10_n961 ) : ( n966 ) ;
assign n968 =  ( n956 ) ? ( bv_4_1_n957 ) : ( n967 ) ;
assign n969 =  ( n932 ) ? ( bv_4_14_n933 ) : ( n968 ) ;
assign n970 =  ( n912 ) ? ( bv_4_6_n913 ) : ( n969 ) ;
assign n971 =  ( n905 ) ? ( bv_4_8_n906 ) : ( n970 ) ;
assign n972 =  ( n893 ) ? ( bv_4_15_n894 ) : ( n971 ) ;
assign n973 =  ( n885 ) ? ( bv_4_12_n886 ) : ( n972 ) ;
assign n974 =  ( n882 ) ? ( bv_4_4_n828 ) : ( n973 ) ;
assign n975 =  ( n881 ) ? ( bv_4_3_n826 ) : ( n974 ) ;
assign n976 =  ( n879 ) ? ( bv_4_9_n880 ) : ( n975 ) ;
assign n977 =  ( n865 ) ? ( bv_4_7_n866 ) : ( n976 ) ;
assign n978 =  ( n851 ) ? ( bv_4_5_n852 ) : ( n977 ) ;
assign n979 =  ( n849 ) ? ( bv_4_13_n850 ) : ( n978 ) ;
assign n980 =  ( n847 ) ? ( bv_4_2_n848 ) : ( n979 ) ;
assign n981 =  ( n252 ) == ( bv_8_164_n41 )  ;
assign n982 =  ( n252 ) == ( bv_8_132_n38 )  ;
assign n983 =  ( n982 ) ? ( bv_4_4_n828 ) : ( bv_4_0_n823 ) ;
assign n984 =  ( n981 ) ? ( bv_4_3_n826 ) : ( n983 ) ;
assign n985 =  ( n252 ) == ( bv_8_164_n41 )  ;
assign n986 =  ( n252 ) == ( bv_8_132_n38 )  ;
assign n987 =  ( n986 ) ? ( bv_4_4_n828 ) : ( bv_4_0_n823 ) ;
assign n988 =  ( n985 ) ? ( bv_4_3_n826 ) : ( n987 ) ;
assign n989 =  ( wait_data ) ? ( cy_sel ) : ( bv_2_0_n9 ) ;
assign n990 =  ( n277 ) == ( bv_5_7_n280 )  ;
assign n991 =  ( n277 ) == ( bv_5_19_n302 )  ;
assign n992 =  ( n990 ) | ( n991 )  ;
assign n993 =  ( n257 ) == ( bv_7_27_n391 )  ;
assign n994 =  ( n992 ) | ( n993 )  ;
assign n995 =  ( n257 ) == ( bv_7_75_n411 )  ;
assign n996 =  ( n994 ) | ( n995 )  ;
assign n997 =  ( n252 ) == ( bv_8_53_n316 )  ;
assign n998 =  ( n996 ) | ( n997 )  ;
assign n999 =  ( n252 ) == ( bv_8_52_n670 )  ;
assign n1000 =  ( n998 ) | ( n999 )  ;
assign n1001 =  ( n252 ) == ( bv_8_130_n326 )  ;
assign n1002 =  ( n1000 ) | ( n1001 )  ;
assign n1003 =  ( n252 ) == ( bv_8_176_n329 )  ;
assign n1004 =  ( n1002 ) | ( n1003 )  ;
assign n1005 =  ( n252 ) == ( bv_8_179_n908 )  ;
assign n1006 =  ( n1004 ) | ( n1005 )  ;
assign n1007 =  ( n252 ) == ( bv_8_212_n556 )  ;
assign n1008 =  ( n1006 ) | ( n1007 )  ;
assign n1009 =  ( n252 ) == ( bv_8_146_n184 )  ;
assign n1010 =  ( n1008 ) | ( n1009 )  ;
assign n1011 =  ( n252 ) == ( bv_8_114_n367 )  ;
assign n1012 =  ( n1010 ) | ( n1011 )  ;
assign n1013 =  ( n252 ) == ( bv_8_160_n370 )  ;
assign n1014 =  ( n1012 ) | ( n1013 )  ;
assign n1015 =  ( n252 ) == ( bv_8_51_n578 )  ;
assign n1016 =  ( n1014 ) | ( n1015 )  ;
assign n1017 =  ( n252 ) == ( bv_8_19_n584 )  ;
assign n1018 =  ( n1016 ) | ( n1017 )  ;
assign n1019 =  ( n252 ) == ( bv_8_149_n377 )  ;
assign n1020 =  ( n1018 ) | ( n1019 )  ;
assign n1021 =  ( n252 ) == ( bv_8_148_n589 )  ;
assign n1022 =  ( n1020 ) | ( n1021 )  ;
assign n1023 =  ( n252 ) == ( bv_8_197_n199 )  ;
assign n1024 =  ( n252 ) == ( bv_8_211_n815 )  ;
assign n1025 =  ( n1023 ) | ( n1024 )  ;
assign n1026 =  ( n252 ) == ( bv_8_210_n196 )  ;
assign n1027 =  ( n1025 ) | ( n1026 )  ;
assign n1028 =  ( n252 ) == ( bv_8_20_n559 )  ;
assign n1029 =  ( n1027 ) | ( n1028 )  ;
assign n1030 =  ( n252 ) == ( bv_8_21_n171 )  ;
assign n1031 =  ( n1029 ) | ( n1030 )  ;
assign n1032 =  ( n252 ) == ( bv_8_213_n70 )  ;
assign n1033 =  ( n1031 ) | ( n1032 )  ;
assign n1034 =  ( n252 ) == ( bv_8_163_n424 )  ;
assign n1035 =  ( n1033 ) | ( n1034 )  ;
assign n1036 =  ( n257 ) == ( bv_7_99_n222 )  ;
assign n1037 =  ( n1035 ) | ( n1036 )  ;
assign n1038 =  ( n277 ) == ( bv_5_3_n138 )  ;
assign n1039 =  ( n1037 ) | ( n1038 )  ;
assign n1040 =  ( n277 ) == ( bv_5_27_n67 )  ;
assign n1041 =  ( n1039 ) | ( n1040 )  ;
assign n1042 =  ( n277 ) == ( bv_5_25_n152 )  ;
assign n1043 =  ( n1041 ) | ( n1042 )  ;
assign n1044 =  ( n257 ) == ( bv_7_11_n208 )  ;
assign n1045 =  ( n1043 ) | ( n1044 )  ;
assign n1046 =  ( n252 ) == ( bv_8_178_n168 )  ;
assign n1047 =  ( n252 ) == ( bv_8_162_n355 )  ;
assign n1048 =  ( n1046 ) | ( n1047 )  ;
assign n1049 =  ( n1048 ) ? ( bv_2_2_n21 ) : ( bv_2_0_n9 ) ;
assign n1050 =  ( n1045 ) ? ( bv_2_3_n6 ) : ( n1049 ) ;
assign n1051 =  ( n1022 ) ? ( bv_2_1_n15 ) : ( n1050 ) ;
assign n1052 =  ( wait_data ) ? ( psw ) : ( bv_2_0_n9 ) ;
assign n1053 =  ( n252 ) == ( bv_8_132_n38 )  ;
assign n1054 =  ( n252 ) == ( bv_8_164_n41 )  ;
assign n1055 =  ( n1053 ) | ( n1054 )  ;
assign n1056 =  ( n1055 ) ? ( bv_2_2_n21 ) : ( bv_2_0_n9 ) ;
assign n1057 =  ( n277 ) == ( bv_5_23_n51 )  ;
assign n1058 =  ( n257 ) == ( bv_7_91_n55 )  ;
assign n1059 =  ( n1057 ) | ( n1058 )  ;
assign n1060 =  ( n252 ) == ( bv_8_130_n326 )  ;
assign n1061 =  ( n1059 ) | ( n1060 )  ;
assign n1062 =  ( n252 ) == ( bv_8_176_n329 )  ;
assign n1063 =  ( n1061 ) | ( n1062 )  ;
assign n1064 =  ( n252 ) == ( bv_8_181_n58 )  ;
assign n1065 =  ( n1063 ) | ( n1064 )  ;
assign n1066 =  ( n252 ) == ( bv_8_180_n61 )  ;
assign n1067 =  ( n1065 ) | ( n1066 )  ;
assign n1068 =  ( n252 ) == ( bv_8_195_n794 )  ;
assign n1069 =  ( n1067 ) | ( n1068 )  ;
assign n1070 =  ( n252 ) == ( bv_8_179_n908 )  ;
assign n1071 =  ( n1069 ) | ( n1070 )  ;
assign n1072 =  ( n252 ) == ( bv_8_212_n556 )  ;
assign n1073 =  ( n1071 ) | ( n1072 )  ;
assign n1074 =  ( n252 ) == ( bv_8_162_n355 )  ;
assign n1075 =  ( n1073 ) | ( n1074 )  ;
assign n1076 =  ( n252 ) == ( bv_8_114_n367 )  ;
assign n1077 =  ( n1075 ) | ( n1076 )  ;
assign n1078 =  ( n252 ) == ( bv_8_160_n370 )  ;
assign n1079 =  ( n1077 ) | ( n1078 )  ;
assign n1080 =  ( n252 ) == ( bv_8_51_n578 )  ;
assign n1081 =  ( n1079 ) | ( n1080 )  ;
assign n1082 =  ( n252 ) == ( bv_8_19_n584 )  ;
assign n1083 =  ( n1081 ) | ( n1082 )  ;
assign n1084 =  ( n252 ) == ( bv_8_211_n815 )  ;
assign n1085 =  ( n1083 ) | ( n1084 )  ;
assign n1086 =  ( n252 ) == ( bv_8_132_n38 )  ;
assign n1087 =  ( n252 ) == ( bv_8_164_n41 )  ;
assign n1088 =  ( n1086 ) | ( n1087 )  ;
assign n1089 =  ( n277 ) == ( bv_5_5_n278 )  ;
assign n1090 =  ( n277 ) == ( bv_5_7_n280 )  ;
assign n1091 =  ( n1089 ) | ( n1090 )  ;
assign n1092 =  ( n277 ) == ( bv_5_19_n302 )  ;
assign n1093 =  ( n1091 ) | ( n1092 )  ;
assign n1094 =  ( n257 ) == ( bv_7_19_n389 )  ;
assign n1095 =  ( n1093 ) | ( n1094 )  ;
assign n1096 =  ( n257 ) == ( bv_7_27_n391 )  ;
assign n1097 =  ( n1095 ) | ( n1096 )  ;
assign n1098 =  ( n257 ) == ( bv_7_75_n411 )  ;
assign n1099 =  ( n1097 ) | ( n1098 )  ;
assign n1100 =  ( n252 ) == ( bv_8_37_n313 )  ;
assign n1101 =  ( n1099 ) | ( n1100 )  ;
assign n1102 =  ( n252 ) == ( bv_8_36_n667 )  ;
assign n1103 =  ( n1101 ) | ( n1102 )  ;
assign n1104 =  ( n252 ) == ( bv_8_53_n316 )  ;
assign n1105 =  ( n1103 ) | ( n1104 )  ;
assign n1106 =  ( n252 ) == ( bv_8_52_n670 )  ;
assign n1107 =  ( n1105 ) | ( n1106 )  ;
assign n1108 =  ( n252 ) == ( bv_8_149_n377 )  ;
assign n1109 =  ( n1107 ) | ( n1108 )  ;
assign n1110 =  ( n252 ) == ( bv_8_148_n589 )  ;
assign n1111 =  ( n1109 ) | ( n1110 )  ;
assign n1112 =  ( n1111 ) ? ( bv_2_3_n6 ) : ( bv_2_0_n9 ) ;
assign n1113 =  ( n1088 ) ? ( bv_2_2_n21 ) : ( n1112 ) ;
assign n1114 =  ( n1085 ) ? ( bv_2_1_n15 ) : ( n1113 ) ;
assign n1115 =  ( n252 ) == ( bv_8_132_n38 )  ;
assign n1116 =  ( n252 ) == ( bv_8_164_n41 )  ;
assign n1117 =  ( n1115 ) | ( n1116 )  ;
assign n1118 =  ( n1117 ) ? ( bv_2_2_n21 ) : ( bv_2_0_n9 ) ;
assign n1119 =  ( n252 ) == ( bv_8_132_n38 )  ;
assign n1120 =  ( n252 ) == ( bv_8_164_n41 )  ;
assign n1121 =  ( n1119 ) | ( n1120 )  ;
assign n1122 =  ( n1121 ) ? ( bv_2_2_n21 ) : ( bv_2_0_n9 ) ;
assign n1123 =  ( wait_data ) ? ( wr ) : ( 1'b0 )  ;
assign n1124 =  ( n46 ) | ( n139 )  ;
assign n1125 =  ( n1124 ) | ( n68 )  ;
assign n1126 =  ( n1125 ) | ( n141 )  ;
assign n1127 =  ( n1126 ) | ( n144 )  ;
assign n1128 =  ( n1127 ) | ( n147 )  ;
assign n1129 =  ( n1128 ) | ( n150 )  ;
assign n1130 =  ( n1129 ) | ( n155 )  ;
assign n1131 =  ( n1130 ) | ( n153 )  ;
assign n1132 =  ( n1131 ) | ( n209 )  ;
assign n1133 =  ( n1132 ) | ( n211 )  ;
assign n1134 =  ( n1133 ) | ( n157 )  ;
assign n1135 =  ( n1134 ) | ( n214 )  ;
assign n1136 =  ( n1135 ) | ( n217 )  ;
assign n1137 =  ( n1136 ) | ( n220 )  ;
assign n1138 =  ( n1137 ) | ( n223 )  ;
assign n1139 =  ( n1138 ) | ( n226 )  ;
assign n1140 =  ( n1139 ) | ( n160 )  ;
assign n1141 =  ( n1140 ) | ( n163 )  ;
assign n1142 =  ( n1141 ) | ( n166 )  ;
assign n1143 =  ( n1142 ) | ( n169 )  ;
assign n1144 =  ( n1143 ) | ( n172 )  ;
assign n1145 =  ( n1144 ) | ( n71 )  ;
assign n1146 =  ( n1145 ) | ( n176 )  ;
assign n1147 =  ( n1146 ) | ( n74 )  ;
assign n1148 =  ( n1147 ) | ( n179 )  ;
assign n1149 =  ( n1148 ) | ( n229 )  ;
assign n1150 =  ( n1149 ) | ( n182 )  ;
assign n1151 =  ( n1150 ) | ( n185 )  ;
assign n1152 =  ( n1151 ) | ( n188 )  ;
assign n1153 =  ( n1152 ) | ( n191 )  ;
assign n1154 =  ( n1153 ) | ( n194 )  ;
assign n1155 =  ( n1154 ) | ( n136 )  ;
assign n1156 =  ( n1155 ) | ( n197 )  ;
assign n1157 =  ( n1156 ) | ( n200 )  ;
assign n1158 =  ( n1157 ) | ( n203 )  ;
assign n1159 =  ( n1158 ) | ( n206 )  ;
assign n1160 =  ( n1159 ) ? ( 1'b1 ) : ( 1'b0 )  ;
assign n1161 =  ( n237 ) | ( n236 )  ;
assign n1162 =  ( n1161 ) ? ( 1'b1 ) : ( 1'b0 )  ;
assign n1163 =  ( n241 ) | ( n242 )  ;
assign n1164 =  ( n1163 ) | ( n244 )  ;
assign n1165 =  ( n1164 ) ? ( 1'b1 ) : ( 1'b0 )  ;
assign n1166 =  ( wait_data ) ? ( wr_sfr ) : ( bv_2_0_n9 ) ;
assign n1167 =  ( n277 ) == ( bv_5_5_n278 )  ;
assign n1168 =  ( n277 ) == ( bv_5_7_n280 )  ;
assign n1169 =  ( n1167 ) | ( n1168 )  ;
assign n1170 =  ( n277 ) == ( bv_5_11_n283 )  ;
assign n1171 =  ( n1169 ) | ( n1170 )  ;
assign n1172 =  ( n277 ) == ( bv_5_29_n294 )  ;
assign n1173 =  ( n1171 ) | ( n1172 )  ;
assign n1174 =  ( n277 ) == ( bv_5_9_n299 )  ;
assign n1175 =  ( n1173 ) | ( n1174 )  ;
assign n1176 =  ( n277 ) == ( bv_5_19_n302 )  ;
assign n1177 =  ( n1175 ) | ( n1176 )  ;
assign n1178 =  ( n277 ) == ( bv_5_13_n307 )  ;
assign n1179 =  ( n1177 ) | ( n1178 )  ;
assign n1180 =  ( n257 ) == ( bv_7_19_n389 )  ;
assign n1181 =  ( n1179 ) | ( n1180 )  ;
assign n1182 =  ( n257 ) == ( bv_7_27_n391 )  ;
assign n1183 =  ( n1181 ) | ( n1182 )  ;
assign n1184 =  ( n257 ) == ( bv_7_43_n394 )  ;
assign n1185 =  ( n1183 ) | ( n1184 )  ;
assign n1186 =  ( n257 ) == ( bv_7_115_n403 )  ;
assign n1187 =  ( n1185 ) | ( n1186 )  ;
assign n1188 =  ( n257 ) == ( bv_7_35_n408 )  ;
assign n1189 =  ( n1187 ) | ( n1188 )  ;
assign n1190 =  ( n257 ) == ( bv_7_75_n411 )  ;
assign n1191 =  ( n1189 ) | ( n1190 )  ;
assign n1192 =  ( n257 ) == ( bv_7_51_n418 )  ;
assign n1193 =  ( n1191 ) | ( n1192 )  ;
assign n1194 =  ( n252 ) == ( bv_8_37_n313 )  ;
assign n1195 =  ( n1193 ) | ( n1194 )  ;
assign n1196 =  ( n252 ) == ( bv_8_36_n667 )  ;
assign n1197 =  ( n1195 ) | ( n1196 )  ;
assign n1198 =  ( n252 ) == ( bv_8_53_n316 )  ;
assign n1199 =  ( n1197 ) | ( n1198 )  ;
assign n1200 =  ( n252 ) == ( bv_8_52_n670 )  ;
assign n1201 =  ( n1199 ) | ( n1200 )  ;
assign n1202 =  ( n252 ) == ( bv_8_85_n319 )  ;
assign n1203 =  ( n1201 ) | ( n1202 )  ;
assign n1204 =  ( n252 ) == ( bv_8_84_n262 )  ;
assign n1205 =  ( n1203 ) | ( n1204 )  ;
assign n1206 =  ( n252 ) == ( bv_8_228_n550 )  ;
assign n1207 =  ( n1205 ) | ( n1206 )  ;
assign n1208 =  ( n252 ) == ( bv_8_244_n553 )  ;
assign n1209 =  ( n1207 ) | ( n1208 )  ;
assign n1210 =  ( n252 ) == ( bv_8_212_n556 )  ;
assign n1211 =  ( n1209 ) | ( n1210 )  ;
assign n1212 =  ( n252 ) == ( bv_8_20_n559 )  ;
assign n1213 =  ( n1211 ) | ( n1212 )  ;
assign n1214 =  ( n252 ) == ( bv_8_4_n564 )  ;
assign n1215 =  ( n1213 ) | ( n1214 )  ;
assign n1216 =  ( n252 ) == ( bv_8_229_n350 )  ;
assign n1217 =  ( n1215 ) | ( n1216 )  ;
assign n1218 =  ( n252 ) == ( bv_8_116_n675 )  ;
assign n1219 =  ( n1217 ) | ( n1218 )  ;
assign n1220 =  ( n252 ) == ( bv_8_69_n360 )  ;
assign n1221 =  ( n1219 ) | ( n1220 )  ;
assign n1222 =  ( n252 ) == ( bv_8_68_n678 )  ;
assign n1223 =  ( n1221 ) | ( n1222 )  ;
assign n1224 =  ( n252 ) == ( bv_8_35_n575 )  ;
assign n1225 =  ( n1223 ) | ( n1224 )  ;
assign n1226 =  ( n252 ) == ( bv_8_51_n578 )  ;
assign n1227 =  ( n1225 ) | ( n1226 )  ;
assign n1228 =  ( n252 ) == ( bv_8_3_n581 )  ;
assign n1229 =  ( n1227 ) | ( n1228 )  ;
assign n1230 =  ( n252 ) == ( bv_8_19_n584 )  ;
assign n1231 =  ( n1229 ) | ( n1230 )  ;
assign n1232 =  ( n252 ) == ( bv_8_149_n377 )  ;
assign n1233 =  ( n1231 ) | ( n1232 )  ;
assign n1234 =  ( n252 ) == ( bv_8_148_n589 )  ;
assign n1235 =  ( n1233 ) | ( n1234 )  ;
assign n1236 =  ( n252 ) == ( bv_8_101_n382 )  ;
assign n1237 =  ( n1235 ) | ( n1236 )  ;
assign n1238 =  ( n252 ) == ( bv_8_100_n681 )  ;
assign n1239 =  ( n1237 ) | ( n1238 )  ;
assign n1240 =  ( n277 ) == ( bv_5_25_n152 )  ;
assign n1241 =  ( n257 ) == ( bv_7_99_n222 )  ;
assign n1242 =  ( n1240 ) | ( n1241 )  ;
assign n1243 =  ( n257 ) == ( bv_7_107_n225 )  ;
assign n1244 =  ( n1242 ) | ( n1243 )  ;
assign n1245 =  ( n252 ) == ( bv_8_196_n592 )  ;
assign n1246 =  ( n1244 ) | ( n1245 )  ;
assign n1247 =  ( n252 ) == ( bv_8_197_n199 )  ;
assign n1248 =  ( n1246 ) | ( n1247 )  ;
assign n1249 =  ( n252 ) == ( bv_8_163_n424 )  ;
assign n1250 =  ( n252 ) == ( bv_8_144_n687 )  ;
assign n1251 =  ( n1249 ) | ( n1250 )  ;
assign n1252 =  ( n1251 ) ? ( bv_2_3_n6 ) : ( bv_2_0_n9 ) ;
assign n1253 =  ( n1248 ) ? ( bv_2_2_n21 ) : ( n1252 ) ;
assign n1254 =  ( n1239 ) ? ( bv_2_1_n15 ) : ( n1253 ) ;
assign n1255 =  ( n252 ) == ( bv_8_147_n27 )  ;
assign n1256 =  ( n252 ) == ( bv_8_131_n29 )  ;
assign n1257 =  ( n1255 ) | ( n1256 )  ;
assign n1258 =  ( n252 ) == ( bv_8_224_n82 )  ;
assign n1259 =  ( n1257 ) | ( n1258 )  ;
assign n1260 =  ( n257 ) == ( bv_7_113_n76 )  ;
assign n1261 =  ( n1259 ) | ( n1260 )  ;
assign n1262 =  ( n252 ) == ( bv_8_132_n38 )  ;
assign n1263 =  ( n252 ) == ( bv_8_164_n41 )  ;
assign n1264 =  ( n1262 ) | ( n1263 )  ;
assign n1265 =  ( n1264 ) ? ( bv_2_2_n21 ) : ( bv_2_0_n9 ) ;
assign n1266 =  ( n1261 ) ? ( bv_2_1_n15 ) : ( n1265 ) ;
always @(posedge clk) begin
   if(rst) begin
   end
   else if(__ILA_DECODER_valid__) begin
       if ( __ILA_DECODER_decode_of_stall__ && __ILA_DECODER_grant__[0] ) begin
           state <= state;
       end else if ( __ILA_DECODER_decode_of_process__ && __ILA_DECODER_grant__[1] ) begin
           state <= bv_2_2_n21;
       end else if ( __ILA_DECODER_decode_of_step_0__ && __ILA_DECODER_grant__[2] ) begin
           state <= n116;
       end else if ( __ILA_DECODER_decode_of_step_1__ && __ILA_DECODER_grant__[3] ) begin
           state <= bv_2_0_n9;
       end else if ( __ILA_DECODER_decode_of_step_2__ && __ILA_DECODER_grant__[4] ) begin
           state <= bv_2_1_n15;
       end
       if ( __ILA_DECODER_decode_of_stall__ && __ILA_DECODER_grant__[0] ) begin
           op <= n118;
       end else if ( __ILA_DECODER_decode_of_step_0__ && __ILA_DECODER_grant__[2] ) begin
           op <= op_in;
       end
       if ( __ILA_DECODER_decode_of_stall__ && __ILA_DECODER_grant__[0] ) begin
           mem_act <= bv_3_7_n119;
       end else if ( __ILA_DECODER_decode_of_process__ && __ILA_DECODER_grant__[1] ) begin
           mem_act <= bv_3_7_n119;
       end else if ( __ILA_DECODER_decode_of_step_0__ && __ILA_DECODER_grant__[2] ) begin
           mem_act <= n132;
       end else if ( __ILA_DECODER_decode_of_step_1__ && __ILA_DECODER_grant__[3] ) begin
           mem_act <= bv_3_7_n119;
       end else if ( __ILA_DECODER_decode_of_step_2__ && __ILA_DECODER_grant__[4] ) begin
           mem_act <= bv_3_7_n119;
       end
       if ( __ILA_DECODER_decode_of_stall__ && __ILA_DECODER_grant__[0] ) begin
           ram_wr_sel <= n133;
       end else if ( __ILA_DECODER_decode_of_process__ && __ILA_DECODER_grant__[1] ) begin
           ram_wr_sel <= bv_3_0_n124;
       end else if ( __ILA_DECODER_decode_of_step_0__ && __ILA_DECODER_grant__[2] ) begin
           ram_wr_sel <= n235;
       end else if ( __ILA_DECODER_decode_of_step_1__ && __ILA_DECODER_grant__[3] ) begin
           ram_wr_sel <= n239;
       end else if ( __ILA_DECODER_decode_of_step_2__ && __ILA_DECODER_grant__[4] ) begin
           ram_wr_sel <= n246;
       end
       if ( __ILA_DECODER_decode_of_stall__ && __ILA_DECODER_grant__[0] ) begin
           ram_rd_sel_r <= n441;
       end else if ( __ILA_DECODER_decode_of_process__ && __ILA_DECODER_grant__[1] ) begin
           ram_rd_sel_r <= n461;
       end else if ( __ILA_DECODER_decode_of_step_0__ && __ILA_DECODER_grant__[2] ) begin
           ram_rd_sel_r <= n441;
       end else if ( __ILA_DECODER_decode_of_step_1__ && __ILA_DECODER_grant__[3] ) begin
           ram_rd_sel_r <= n465;
       end else if ( __ILA_DECODER_decode_of_step_2__ && __ILA_DECODER_grant__[4] ) begin
           ram_rd_sel_r <= n504;
       end
       if ( __ILA_DECODER_decode_of_stall__ && __ILA_DECODER_grant__[0] ) begin
           src_sel1 <= n505;
       end else if ( __ILA_DECODER_decode_of_process__ && __ILA_DECODER_grant__[1] ) begin
           src_sel1 <= n513;
       end else if ( __ILA_DECODER_decode_of_step_0__ && __ILA_DECODER_grant__[2] ) begin
           src_sel1 <= n698;
       end else if ( __ILA_DECODER_decode_of_step_1__ && __ILA_DECODER_grant__[3] ) begin
           src_sel1 <= n710;
       end else if ( __ILA_DECODER_decode_of_step_2__ && __ILA_DECODER_grant__[4] ) begin
           src_sel1 <= n720;
       end
       if ( __ILA_DECODER_decode_of_stall__ && __ILA_DECODER_grant__[0] ) begin
           src_sel2 <= n721;
       end else if ( __ILA_DECODER_decode_of_process__ && __ILA_DECODER_grant__[1] ) begin
           src_sel2 <= bv_2_0_n9;
       end else if ( __ILA_DECODER_decode_of_step_0__ && __ILA_DECODER_grant__[2] ) begin
           src_sel2 <= n791;
       end else if ( __ILA_DECODER_decode_of_step_1__ && __ILA_DECODER_grant__[3] ) begin
           src_sel2 <= bv_2_0_n9;
       end else if ( __ILA_DECODER_decode_of_step_2__ && __ILA_DECODER_grant__[4] ) begin
           src_sel2 <= bv_2_0_n9;
       end
       if ( __ILA_DECODER_decode_of_stall__ && __ILA_DECODER_grant__[0] ) begin
           src_sel3 <= n792;
       end else if ( __ILA_DECODER_decode_of_process__ && __ILA_DECODER_grant__[1] ) begin
           src_sel3 <= 1'b0;
       end else if ( __ILA_DECODER_decode_of_step_0__ && __ILA_DECODER_grant__[2] ) begin
           src_sel3 <= n822;
       end else if ( __ILA_DECODER_decode_of_step_1__ && __ILA_DECODER_grant__[3] ) begin
           src_sel3 <= 1'b0;
       end else if ( __ILA_DECODER_decode_of_step_2__ && __ILA_DECODER_grant__[4] ) begin
           src_sel3 <= 1'b0;
       end
       if ( __ILA_DECODER_decode_of_stall__ && __ILA_DECODER_grant__[0] ) begin
           alu_op <= n824;
       end else if ( __ILA_DECODER_decode_of_process__ && __ILA_DECODER_grant__[1] ) begin
           alu_op <= n830;
       end else if ( __ILA_DECODER_decode_of_step_0__ && __ILA_DECODER_grant__[2] ) begin
           alu_op <= n980;
       end else if ( __ILA_DECODER_decode_of_step_1__ && __ILA_DECODER_grant__[3] ) begin
           alu_op <= n984;
       end else if ( __ILA_DECODER_decode_of_step_2__ && __ILA_DECODER_grant__[4] ) begin
           alu_op <= n988;
       end
       if ( __ILA_DECODER_decode_of_stall__ && __ILA_DECODER_grant__[0] ) begin
           cy_sel <= n989;
       end else if ( __ILA_DECODER_decode_of_process__ && __ILA_DECODER_grant__[1] ) begin
           cy_sel <= bv_2_0_n9;
       end else if ( __ILA_DECODER_decode_of_step_0__ && __ILA_DECODER_grant__[2] ) begin
           cy_sel <= n1051;
       end else if ( __ILA_DECODER_decode_of_step_1__ && __ILA_DECODER_grant__[3] ) begin
           cy_sel <= bv_2_0_n9;
       end else if ( __ILA_DECODER_decode_of_step_2__ && __ILA_DECODER_grant__[4] ) begin
           cy_sel <= bv_2_0_n9;
       end
       if ( __ILA_DECODER_decode_of_stall__ && __ILA_DECODER_grant__[0] ) begin
           psw <= n1052;
       end else if ( __ILA_DECODER_decode_of_process__ && __ILA_DECODER_grant__[1] ) begin
           psw <= n1056;
       end else if ( __ILA_DECODER_decode_of_step_0__ && __ILA_DECODER_grant__[2] ) begin
           psw <= n1114;
       end else if ( __ILA_DECODER_decode_of_step_1__ && __ILA_DECODER_grant__[3] ) begin
           psw <= n1118;
       end else if ( __ILA_DECODER_decode_of_step_2__ && __ILA_DECODER_grant__[4] ) begin
           psw <= n1122;
       end
       if ( __ILA_DECODER_decode_of_stall__ && __ILA_DECODER_grant__[0] ) begin
           wr <= n1123;
       end else if ( __ILA_DECODER_decode_of_process__ && __ILA_DECODER_grant__[1] ) begin
           wr <= 1'b0;
       end else if ( __ILA_DECODER_decode_of_step_0__ && __ILA_DECODER_grant__[2] ) begin
           wr <= n1160;
       end else if ( __ILA_DECODER_decode_of_step_1__ && __ILA_DECODER_grant__[3] ) begin
           wr <= n1162;
       end else if ( __ILA_DECODER_decode_of_step_2__ && __ILA_DECODER_grant__[4] ) begin
           wr <= n1165;
       end
       if ( __ILA_DECODER_decode_of_stall__ && __ILA_DECODER_grant__[0] ) begin
           wr_sfr <= n1166;
       end else if ( __ILA_DECODER_decode_of_process__ && __ILA_DECODER_grant__[1] ) begin
           wr_sfr <= bv_2_0_n9;
       end else if ( __ILA_DECODER_decode_of_step_0__ && __ILA_DECODER_grant__[2] ) begin
           wr_sfr <= n1254;
       end else if ( __ILA_DECODER_decode_of_step_1__ && __ILA_DECODER_grant__[3] ) begin
           wr_sfr <= n1266;
       end else if ( __ILA_DECODER_decode_of_step_2__ && __ILA_DECODER_grant__[4] ) begin
           wr_sfr <= bv_2_0_n9;
       end
   end
end
endmodule
