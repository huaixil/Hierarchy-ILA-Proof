/* PREHEADER */
module fun_Adptfloat2Fixed (
    input [7:0] arg0,
    input [2:0] arg1,
    output [19:0] result
);
//TODO: Add the specific function HERE.
endmodule
module fun_Fixed2Adaptfloat (
    input [19:0] arg0,
    input [2:0] arg1,
    output [7:0] result
);
//TODO: Add the specific function HERE.
endmodule
module fun_PEActEadd (
    input [19:0] arg0,
    input [19:0] arg1,
    output [19:0] result
);
//TODO: Add the specific function HERE.
endmodule
module fun_PEActEmul (
    input [19:0] arg0,
    input [19:0] arg1,
    output [19:0] result
);
//TODO: Add the specific function HERE.
endmodule
module fun_PEActSigmoid (
    input [19:0] arg0,
    output [19:0] result
);
//TODO: Add the specific function HERE.
endmodule
module fun_PEActTanh (
    input [19:0] arg0,
    output [19:0] result
);
//TODO: Add the specific function HERE.
endmodule
module fun_PEActRelu (
    input [19:0] arg0,
    output [19:0] result
);
//TODO: Add the specific function HERE.
endmodule
module fun_PEActOnex (
    input [19:0] arg0,
    output [19:0] result
);
//TODO: Add the specific function HERE.
endmodule

/* END OF PREHEADER */
module pe_act(
PE0_core_act_vector_0,
PE0_core_act_vector_1,
PE0_core_act_vector_10,
PE0_core_act_vector_11,
PE0_core_act_vector_12,
PE0_core_act_vector_13,
PE0_core_act_vector_14,
PE0_core_act_vector_15,
PE0_core_act_vector_2,
PE0_core_act_vector_3,
PE0_core_act_vector_4,
PE0_core_act_vector_5,
PE0_core_act_vector_6,
PE0_core_act_vector_7,
PE0_core_act_vector_8,
PE0_core_act_vector_9,
__ILA_pe_act_grant__,
act_start,
act_start_valid,
addr,
axi_rw,
clk,
data_in_0,
data_in_1,
data_in_10,
data_in_11,
data_in_12,
data_in_13,
data_in_14,
data_in_15,
data_in_2,
data_in_3,
data_in_4,
data_in_5,
data_in_6,
data_in_7,
data_in_8,
data_in_9,
done_ready,
output_port_ready,
pe0_act_reg_port_valid,
rst,
rva_in_valid,
wstrb,
__ILA_pe_act_acc_decode__,
__ILA_pe_act_decode_of_PE0_ACT_STORE_BUFFER__,
__ILA_pe_act_decode_of_PE0_CONFIG_ACT_MNGR__,
__ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_0_15__,
__ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_16_31__,
__ILA_pe_act_decode_of_PE0_act_child_done_sent__,
__ILA_pe_act_decode_of_PE0_act_child_initiate__,
__ILA_pe_act_decode_of_PE0_act_child_op_copy__,
__ILA_pe_act_decode_of_PE0_act_child_op_eadd__,
__ILA_pe_act_decode_of_PE0_act_child_op_emul__,
__ILA_pe_act_decode_of_PE0_act_child_op_inpe__,
__ILA_pe_act_decode_of_PE0_act_child_op_load__,
__ILA_pe_act_decode_of_PE0_act_child_op_load_zero__,
__ILA_pe_act_decode_of_PE0_act_child_op_onex__,
__ILA_pe_act_decode_of_PE0_act_child_op_outgb__,
__ILA_pe_act_decode_of_PE0_act_child_op_relu__,
__ILA_pe_act_decode_of_PE0_act_child_op_sigm__,
__ILA_pe_act_decode_of_PE0_act_child_op_store__,
__ILA_pe_act_decode_of_PE0_act_child_op_tanh__,
__ILA_pe_act_decode_of_PE0_act_child_out_sent__,
__ILA_pe_act_decode_of_PE0_act_child_reg_store__,
__ILA_pe_act_valid__,
PE0_act_regs_3_data_n405,
PE0_act_regs_2_data_n409,
PE0_act_regs_1_data_n413,
PE0_act_regs_0_data_n417,
PE0_act_regs_3_data_n432,
PE0_act_regs_2_data_n436,
PE0_act_regs_1_data_n440,
PE0_act_regs_0_data_n444,
PE0_act_regs_3_data_n457,
PE0_act_regs_2_data_n461,
PE0_act_regs_1_data_n465,
PE0_act_regs_0_data_n469,
PE0_act_regs_3_data_n482,
PE0_act_regs_2_data_n486,
PE0_act_regs_1_data_n490,
PE0_act_regs_0_data_n494,
PE0_act_regs_3_data_n507,
PE0_act_regs_2_data_n511,
PE0_act_regs_1_data_n515,
PE0_act_regs_0_data_n519,
PE0_act_regs_3_data_n532,
PE0_act_regs_2_data_n536,
PE0_act_regs_1_data_n540,
PE0_act_regs_0_data_n544,
PE0_act_regs_3_data_n557,
PE0_act_regs_2_data_n561,
PE0_act_regs_1_data_n565,
PE0_act_regs_0_data_n569,
PE0_act_regs_3_data_n582,
PE0_act_regs_2_data_n586,
PE0_act_regs_1_data_n590,
PE0_act_regs_0_data_n594,
PE0_act_regs_3_data_n607,
PE0_act_regs_2_data_n611,
PE0_act_regs_1_data_n615,
PE0_act_regs_0_data_n619,
PE0_act_regs_3_data_n633,
PE0_act_regs_2_data_n637,
PE0_act_regs_1_data_n641,
PE0_act_regs_0_data_n645,
PE0_act_regs_3_data_n659,
PE0_act_regs_2_data_n663,
PE0_act_regs_1_data_n667,
PE0_act_regs_0_data_n671,
PE0_act_regs_3_data_n684,
PE0_act_regs_2_data_n688,
PE0_act_regs_1_data_n692,
PE0_act_regs_0_data_n696,
PE0_act_regs_3_data_n709,
PE0_act_regs_2_data_n713,
PE0_act_regs_1_data_n717,
PE0_act_regs_0_data_n721,
PE0_act_regs_3_data_n734,
PE0_act_regs_2_data_n738,
PE0_act_regs_1_data_n742,
PE0_act_regs_0_data_n746,
PE0_act_regs_3_data_n759,
PE0_act_regs_2_data_n763,
PE0_act_regs_1_data_n767,
PE0_act_regs_0_data_n771,
PE0_act_regs_3_data_n784,
PE0_act_regs_2_data_n788,
PE0_act_regs_1_data_n792,
PE0_act_regs_0_data_n796,
pe0_act_buffer_data_n1036,
PE0_act_regs_3_data_n1045,
PE0_act_regs_2_data_n1049,
PE0_act_regs_1_data_n1053,
PE0_act_regs_0_data_n1057,
PE0_act_regs_3_data_n1066,
PE0_act_regs_2_data_n1070,
PE0_act_regs_1_data_n1074,
PE0_act_regs_0_data_n1078,
PE0_act_regs_3_data_n1086,
PE0_act_regs_2_data_n1090,
PE0_act_regs_1_data_n1094,
PE0_act_regs_0_data_n1098,
PE0_act_regs_3_data_n1110,
PE0_act_regs_2_data_n1114,
PE0_act_regs_1_data_n1118,
PE0_act_regs_0_data_n1122,
PE0_act_regs_3_data_n1130,
PE0_act_regs_2_data_n1134,
PE0_act_regs_1_data_n1138,
PE0_act_regs_0_data_n1142,
PE0_act_regs_3_data_n1154,
PE0_act_regs_2_data_n1158,
PE0_act_regs_1_data_n1162,
PE0_act_regs_0_data_n1166,
PE0_act_regs_3_data_n1178,
PE0_act_regs_2_data_n1182,
PE0_act_regs_1_data_n1186,
PE0_act_regs_0_data_n1190,
PE0_act_regs_3_data_n1202,
PE0_act_regs_2_data_n1206,
PE0_act_regs_1_data_n1210,
PE0_act_regs_0_data_n1214,
PE0_act_regs_3_data_n1226,
PE0_act_regs_2_data_n1230,
PE0_act_regs_1_data_n1234,
PE0_act_regs_0_data_n1238,
pe0_act_buffer_data_n1250,
PE0_act_regs_3_data_n1258,
PE0_act_regs_2_data_n1262,
PE0_act_regs_1_data_n1266,
PE0_act_regs_0_data_n1270,
PE0_act_regs_3_data_n1279,
PE0_act_regs_2_data_n1283,
PE0_act_regs_1_data_n1287,
PE0_act_regs_0_data_n1291,
PE0_act_regs_3_data_n1299,
PE0_act_regs_2_data_n1303,
PE0_act_regs_1_data_n1307,
PE0_act_regs_0_data_n1311,
PE0_act_regs_3_data_n1323,
PE0_act_regs_2_data_n1327,
PE0_act_regs_1_data_n1331,
PE0_act_regs_0_data_n1335,
PE0_act_regs_3_data_n1343,
PE0_act_regs_2_data_n1347,
PE0_act_regs_1_data_n1351,
PE0_act_regs_0_data_n1355,
PE0_act_regs_3_data_n1367,
PE0_act_regs_2_data_n1371,
PE0_act_regs_1_data_n1375,
PE0_act_regs_0_data_n1379,
PE0_act_regs_3_data_n1391,
PE0_act_regs_2_data_n1395,
PE0_act_regs_1_data_n1399,
PE0_act_regs_0_data_n1403,
PE0_act_regs_3_data_n1415,
PE0_act_regs_2_data_n1419,
PE0_act_regs_1_data_n1423,
PE0_act_regs_0_data_n1427,
PE0_act_regs_3_data_n1439,
PE0_act_regs_2_data_n1443,
PE0_act_regs_1_data_n1447,
PE0_act_regs_0_data_n1451,
pe0_act_buffer_data_n1463,
PE0_act_regs_3_data_n1471,
PE0_act_regs_2_data_n1475,
PE0_act_regs_1_data_n1479,
PE0_act_regs_0_data_n1483,
PE0_act_regs_3_data_n1492,
PE0_act_regs_2_data_n1496,
PE0_act_regs_1_data_n1500,
PE0_act_regs_0_data_n1504,
PE0_act_regs_3_data_n1512,
PE0_act_regs_2_data_n1516,
PE0_act_regs_1_data_n1520,
PE0_act_regs_0_data_n1524,
PE0_act_regs_3_data_n1536,
PE0_act_regs_2_data_n1540,
PE0_act_regs_1_data_n1544,
PE0_act_regs_0_data_n1548,
PE0_act_regs_3_data_n1556,
PE0_act_regs_2_data_n1560,
PE0_act_regs_1_data_n1564,
PE0_act_regs_0_data_n1568,
PE0_act_regs_3_data_n1580,
PE0_act_regs_2_data_n1584,
PE0_act_regs_1_data_n1588,
PE0_act_regs_0_data_n1592,
PE0_act_regs_3_data_n1604,
PE0_act_regs_2_data_n1608,
PE0_act_regs_1_data_n1612,
PE0_act_regs_0_data_n1616,
PE0_act_regs_3_data_n1628,
PE0_act_regs_2_data_n1632,
PE0_act_regs_1_data_n1636,
PE0_act_regs_0_data_n1640,
PE0_act_regs_3_data_n1652,
PE0_act_regs_2_data_n1656,
PE0_act_regs_1_data_n1660,
PE0_act_regs_0_data_n1664,
pe0_act_buffer_data_n1676,
PE0_act_regs_3_data_n1684,
PE0_act_regs_2_data_n1688,
PE0_act_regs_1_data_n1692,
PE0_act_regs_0_data_n1696,
PE0_act_regs_3_data_n1705,
PE0_act_regs_2_data_n1709,
PE0_act_regs_1_data_n1713,
PE0_act_regs_0_data_n1717,
PE0_act_regs_3_data_n1725,
PE0_act_regs_2_data_n1729,
PE0_act_regs_1_data_n1733,
PE0_act_regs_0_data_n1737,
PE0_act_regs_3_data_n1749,
PE0_act_regs_2_data_n1753,
PE0_act_regs_1_data_n1757,
PE0_act_regs_0_data_n1761,
PE0_act_regs_3_data_n1769,
PE0_act_regs_2_data_n1773,
PE0_act_regs_1_data_n1777,
PE0_act_regs_0_data_n1781,
PE0_act_regs_3_data_n1793,
PE0_act_regs_2_data_n1797,
PE0_act_regs_1_data_n1801,
PE0_act_regs_0_data_n1805,
PE0_act_regs_3_data_n1817,
PE0_act_regs_2_data_n1821,
PE0_act_regs_1_data_n1825,
PE0_act_regs_0_data_n1829,
PE0_act_regs_3_data_n1841,
PE0_act_regs_2_data_n1845,
PE0_act_regs_1_data_n1849,
PE0_act_regs_0_data_n1853,
PE0_act_regs_3_data_n1865,
PE0_act_regs_2_data_n1869,
PE0_act_regs_1_data_n1873,
PE0_act_regs_0_data_n1877,
pe0_act_buffer_data_n1889,
PE0_act_regs_3_data_n1897,
PE0_act_regs_2_data_n1901,
PE0_act_regs_1_data_n1905,
PE0_act_regs_0_data_n1909,
PE0_act_regs_3_data_n1918,
PE0_act_regs_2_data_n1922,
PE0_act_regs_1_data_n1926,
PE0_act_regs_0_data_n1930,
PE0_act_regs_3_data_n1938,
PE0_act_regs_2_data_n1942,
PE0_act_regs_1_data_n1946,
PE0_act_regs_0_data_n1950,
PE0_act_regs_3_data_n1962,
PE0_act_regs_2_data_n1966,
PE0_act_regs_1_data_n1970,
PE0_act_regs_0_data_n1974,
PE0_act_regs_3_data_n1982,
PE0_act_regs_2_data_n1986,
PE0_act_regs_1_data_n1990,
PE0_act_regs_0_data_n1994,
PE0_act_regs_3_data_n2006,
PE0_act_regs_2_data_n2010,
PE0_act_regs_1_data_n2014,
PE0_act_regs_0_data_n2018,
PE0_act_regs_3_data_n2030,
PE0_act_regs_2_data_n2034,
PE0_act_regs_1_data_n2038,
PE0_act_regs_0_data_n2042,
PE0_act_regs_3_data_n2054,
PE0_act_regs_2_data_n2058,
PE0_act_regs_1_data_n2062,
PE0_act_regs_0_data_n2066,
PE0_act_regs_3_data_n2078,
PE0_act_regs_2_data_n2082,
PE0_act_regs_1_data_n2086,
PE0_act_regs_0_data_n2090,
pe0_act_buffer_data_n2102,
PE0_act_regs_3_data_n2110,
PE0_act_regs_2_data_n2114,
PE0_act_regs_1_data_n2118,
PE0_act_regs_0_data_n2122,
PE0_act_regs_3_data_n2131,
PE0_act_regs_2_data_n2135,
PE0_act_regs_1_data_n2139,
PE0_act_regs_0_data_n2143,
PE0_act_regs_3_data_n2151,
PE0_act_regs_2_data_n2155,
PE0_act_regs_1_data_n2159,
PE0_act_regs_0_data_n2163,
PE0_act_regs_3_data_n2175,
PE0_act_regs_2_data_n2179,
PE0_act_regs_1_data_n2183,
PE0_act_regs_0_data_n2187,
PE0_act_regs_3_data_n2195,
PE0_act_regs_2_data_n2199,
PE0_act_regs_1_data_n2203,
PE0_act_regs_0_data_n2207,
PE0_act_regs_3_data_n2219,
PE0_act_regs_2_data_n2223,
PE0_act_regs_1_data_n2227,
PE0_act_regs_0_data_n2231,
PE0_act_regs_3_data_n2243,
PE0_act_regs_2_data_n2247,
PE0_act_regs_1_data_n2251,
PE0_act_regs_0_data_n2255,
PE0_act_regs_3_data_n2267,
PE0_act_regs_2_data_n2271,
PE0_act_regs_1_data_n2275,
PE0_act_regs_0_data_n2279,
PE0_act_regs_3_data_n2291,
PE0_act_regs_2_data_n2295,
PE0_act_regs_1_data_n2299,
PE0_act_regs_0_data_n2303,
pe0_act_buffer_data_n2315,
PE0_act_regs_3_data_n2323,
PE0_act_regs_2_data_n2327,
PE0_act_regs_1_data_n2331,
PE0_act_regs_0_data_n2335,
PE0_act_regs_3_data_n2344,
PE0_act_regs_2_data_n2348,
PE0_act_regs_1_data_n2352,
PE0_act_regs_0_data_n2356,
PE0_act_regs_3_data_n2364,
PE0_act_regs_2_data_n2368,
PE0_act_regs_1_data_n2372,
PE0_act_regs_0_data_n2376,
PE0_act_regs_3_data_n2388,
PE0_act_regs_2_data_n2392,
PE0_act_regs_1_data_n2396,
PE0_act_regs_0_data_n2400,
PE0_act_regs_3_data_n2408,
PE0_act_regs_2_data_n2412,
PE0_act_regs_1_data_n2416,
PE0_act_regs_0_data_n2420,
PE0_act_regs_3_data_n2432,
PE0_act_regs_2_data_n2436,
PE0_act_regs_1_data_n2440,
PE0_act_regs_0_data_n2444,
PE0_act_regs_3_data_n2456,
PE0_act_regs_2_data_n2460,
PE0_act_regs_1_data_n2464,
PE0_act_regs_0_data_n2468,
PE0_act_regs_3_data_n2480,
PE0_act_regs_2_data_n2484,
PE0_act_regs_1_data_n2488,
PE0_act_regs_0_data_n2492,
PE0_act_regs_3_data_n2504,
PE0_act_regs_2_data_n2508,
PE0_act_regs_1_data_n2512,
PE0_act_regs_0_data_n2516,
pe0_act_buffer_data_n2528,
PE0_act_regs_3_data_n2536,
PE0_act_regs_2_data_n2540,
PE0_act_regs_1_data_n2544,
PE0_act_regs_0_data_n2548,
PE0_act_regs_3_data_n2557,
PE0_act_regs_2_data_n2561,
PE0_act_regs_1_data_n2565,
PE0_act_regs_0_data_n2569,
PE0_act_regs_3_data_n2577,
PE0_act_regs_2_data_n2581,
PE0_act_regs_1_data_n2585,
PE0_act_regs_0_data_n2589,
PE0_act_regs_3_data_n2601,
PE0_act_regs_2_data_n2605,
PE0_act_regs_1_data_n2609,
PE0_act_regs_0_data_n2613,
PE0_act_regs_3_data_n2621,
PE0_act_regs_2_data_n2625,
PE0_act_regs_1_data_n2629,
PE0_act_regs_0_data_n2633,
PE0_act_regs_3_data_n2645,
PE0_act_regs_2_data_n2649,
PE0_act_regs_1_data_n2653,
PE0_act_regs_0_data_n2657,
PE0_act_regs_3_data_n2669,
PE0_act_regs_2_data_n2673,
PE0_act_regs_1_data_n2677,
PE0_act_regs_0_data_n2681,
PE0_act_regs_3_data_n2693,
PE0_act_regs_2_data_n2697,
PE0_act_regs_1_data_n2701,
PE0_act_regs_0_data_n2705,
PE0_act_regs_3_data_n2717,
PE0_act_regs_2_data_n2721,
PE0_act_regs_1_data_n2725,
PE0_act_regs_0_data_n2729,
pe0_act_buffer_data_n2741,
PE0_act_regs_3_data_n2749,
PE0_act_regs_2_data_n2753,
PE0_act_regs_1_data_n2757,
PE0_act_regs_0_data_n2761,
PE0_act_regs_3_data_n2770,
PE0_act_regs_2_data_n2774,
PE0_act_regs_1_data_n2778,
PE0_act_regs_0_data_n2782,
PE0_act_regs_3_data_n2790,
PE0_act_regs_2_data_n2794,
PE0_act_regs_1_data_n2798,
PE0_act_regs_0_data_n2802,
PE0_act_regs_3_data_n2814,
PE0_act_regs_2_data_n2818,
PE0_act_regs_1_data_n2822,
PE0_act_regs_0_data_n2826,
PE0_act_regs_3_data_n2834,
PE0_act_regs_2_data_n2838,
PE0_act_regs_1_data_n2842,
PE0_act_regs_0_data_n2846,
PE0_act_regs_3_data_n2858,
PE0_act_regs_2_data_n2862,
PE0_act_regs_1_data_n2866,
PE0_act_regs_0_data_n2870,
PE0_act_regs_3_data_n2882,
PE0_act_regs_2_data_n2886,
PE0_act_regs_1_data_n2890,
PE0_act_regs_0_data_n2894,
PE0_act_regs_3_data_n2906,
PE0_act_regs_2_data_n2910,
PE0_act_regs_1_data_n2914,
PE0_act_regs_0_data_n2918,
PE0_act_regs_3_data_n2930,
PE0_act_regs_2_data_n2934,
PE0_act_regs_1_data_n2938,
PE0_act_regs_0_data_n2942,
pe0_act_buffer_data_n2954,
PE0_act_regs_3_data_n2962,
PE0_act_regs_2_data_n2966,
PE0_act_regs_1_data_n2970,
PE0_act_regs_0_data_n2974,
PE0_act_regs_3_data_n2983,
PE0_act_regs_2_data_n2987,
PE0_act_regs_1_data_n2991,
PE0_act_regs_0_data_n2995,
PE0_act_regs_3_data_n3003,
PE0_act_regs_2_data_n3007,
PE0_act_regs_1_data_n3011,
PE0_act_regs_0_data_n3015,
PE0_act_regs_3_data_n3027,
PE0_act_regs_2_data_n3031,
PE0_act_regs_1_data_n3035,
PE0_act_regs_0_data_n3039,
PE0_act_regs_3_data_n3047,
PE0_act_regs_2_data_n3051,
PE0_act_regs_1_data_n3055,
PE0_act_regs_0_data_n3059,
PE0_act_regs_3_data_n3071,
PE0_act_regs_2_data_n3075,
PE0_act_regs_1_data_n3079,
PE0_act_regs_0_data_n3083,
PE0_act_regs_3_data_n3095,
PE0_act_regs_2_data_n3099,
PE0_act_regs_1_data_n3103,
PE0_act_regs_0_data_n3107,
PE0_act_regs_3_data_n3119,
PE0_act_regs_2_data_n3123,
PE0_act_regs_1_data_n3127,
PE0_act_regs_0_data_n3131,
PE0_act_regs_3_data_n3143,
PE0_act_regs_2_data_n3147,
PE0_act_regs_1_data_n3151,
PE0_act_regs_0_data_n3155,
pe0_act_buffer_data_n3167,
PE0_act_regs_3_data_n3175,
PE0_act_regs_2_data_n3179,
PE0_act_regs_1_data_n3183,
PE0_act_regs_0_data_n3187,
PE0_act_regs_3_data_n3196,
PE0_act_regs_2_data_n3200,
PE0_act_regs_1_data_n3204,
PE0_act_regs_0_data_n3208,
PE0_act_regs_3_data_n3216,
PE0_act_regs_2_data_n3220,
PE0_act_regs_1_data_n3224,
PE0_act_regs_0_data_n3228,
PE0_act_regs_3_data_n3240,
PE0_act_regs_2_data_n3244,
PE0_act_regs_1_data_n3248,
PE0_act_regs_0_data_n3252,
PE0_act_regs_3_data_n3260,
PE0_act_regs_2_data_n3264,
PE0_act_regs_1_data_n3268,
PE0_act_regs_0_data_n3272,
PE0_act_regs_3_data_n3284,
PE0_act_regs_2_data_n3288,
PE0_act_regs_1_data_n3292,
PE0_act_regs_0_data_n3296,
PE0_act_regs_3_data_n3308,
PE0_act_regs_2_data_n3312,
PE0_act_regs_1_data_n3316,
PE0_act_regs_0_data_n3320,
PE0_act_regs_3_data_n3332,
PE0_act_regs_2_data_n3336,
PE0_act_regs_1_data_n3340,
PE0_act_regs_0_data_n3344,
PE0_act_regs_3_data_n3356,
PE0_act_regs_2_data_n3360,
PE0_act_regs_1_data_n3364,
PE0_act_regs_0_data_n3368,
pe0_act_buffer_data_n3380,
PE0_act_regs_3_data_n3388,
PE0_act_regs_2_data_n3392,
PE0_act_regs_1_data_n3396,
PE0_act_regs_0_data_n3400,
PE0_act_regs_3_data_n3409,
PE0_act_regs_2_data_n3413,
PE0_act_regs_1_data_n3417,
PE0_act_regs_0_data_n3421,
PE0_act_regs_3_data_n3429,
PE0_act_regs_2_data_n3433,
PE0_act_regs_1_data_n3437,
PE0_act_regs_0_data_n3441,
PE0_act_regs_3_data_n3453,
PE0_act_regs_2_data_n3457,
PE0_act_regs_1_data_n3461,
PE0_act_regs_0_data_n3465,
PE0_act_regs_3_data_n3473,
PE0_act_regs_2_data_n3477,
PE0_act_regs_1_data_n3481,
PE0_act_regs_0_data_n3485,
PE0_act_regs_3_data_n3497,
PE0_act_regs_2_data_n3501,
PE0_act_regs_1_data_n3505,
PE0_act_regs_0_data_n3509,
PE0_act_regs_3_data_n3521,
PE0_act_regs_2_data_n3525,
PE0_act_regs_1_data_n3529,
PE0_act_regs_0_data_n3533,
PE0_act_regs_3_data_n3545,
PE0_act_regs_2_data_n3549,
PE0_act_regs_1_data_n3553,
PE0_act_regs_0_data_n3557,
PE0_act_regs_3_data_n3569,
PE0_act_regs_2_data_n3573,
PE0_act_regs_1_data_n3577,
PE0_act_regs_0_data_n3581,
pe0_act_buffer_data_n3593,
PE0_act_regs_3_data_n3601,
PE0_act_regs_2_data_n3605,
PE0_act_regs_1_data_n3609,
PE0_act_regs_0_data_n3613,
PE0_act_regs_3_data_n3622,
PE0_act_regs_2_data_n3626,
PE0_act_regs_1_data_n3630,
PE0_act_regs_0_data_n3634,
PE0_act_regs_3_data_n3642,
PE0_act_regs_2_data_n3646,
PE0_act_regs_1_data_n3650,
PE0_act_regs_0_data_n3654,
PE0_act_regs_3_data_n3666,
PE0_act_regs_2_data_n3670,
PE0_act_regs_1_data_n3674,
PE0_act_regs_0_data_n3678,
PE0_act_regs_3_data_n3686,
PE0_act_regs_2_data_n3690,
PE0_act_regs_1_data_n3694,
PE0_act_regs_0_data_n3698,
PE0_act_regs_3_data_n3710,
PE0_act_regs_2_data_n3714,
PE0_act_regs_1_data_n3718,
PE0_act_regs_0_data_n3722,
PE0_act_regs_3_data_n3734,
PE0_act_regs_2_data_n3738,
PE0_act_regs_1_data_n3742,
PE0_act_regs_0_data_n3746,
PE0_act_regs_3_data_n3758,
PE0_act_regs_2_data_n3762,
PE0_act_regs_1_data_n3766,
PE0_act_regs_0_data_n3770,
PE0_act_regs_3_data_n3782,
PE0_act_regs_2_data_n3786,
PE0_act_regs_1_data_n3790,
PE0_act_regs_0_data_n3794,
pe0_act_buffer_data_n3806,
PE0_act_regs_3_data_n3814,
PE0_act_regs_2_data_n3818,
PE0_act_regs_1_data_n3822,
PE0_act_regs_0_data_n3826,
PE0_act_regs_3_data_n3835,
PE0_act_regs_2_data_n3839,
PE0_act_regs_1_data_n3843,
PE0_act_regs_0_data_n3847,
PE0_act_regs_3_data_n3855,
PE0_act_regs_2_data_n3859,
PE0_act_regs_1_data_n3863,
PE0_act_regs_0_data_n3867,
PE0_act_regs_3_data_n3879,
PE0_act_regs_2_data_n3883,
PE0_act_regs_1_data_n3887,
PE0_act_regs_0_data_n3891,
PE0_act_regs_3_data_n3899,
PE0_act_regs_2_data_n3903,
PE0_act_regs_1_data_n3907,
PE0_act_regs_0_data_n3911,
PE0_act_regs_3_data_n3923,
PE0_act_regs_2_data_n3927,
PE0_act_regs_1_data_n3931,
PE0_act_regs_0_data_n3935,
PE0_act_regs_3_data_n3947,
PE0_act_regs_2_data_n3951,
PE0_act_regs_1_data_n3955,
PE0_act_regs_0_data_n3959,
PE0_act_regs_3_data_n3971,
PE0_act_regs_2_data_n3975,
PE0_act_regs_1_data_n3979,
PE0_act_regs_0_data_n3983,
PE0_act_regs_3_data_n3995,
PE0_act_regs_2_data_n3999,
PE0_act_regs_1_data_n4003,
PE0_act_regs_0_data_n4007,
pe0_act_buffer_data_n4019,
PE0_act_regs_3_data_n4027,
PE0_act_regs_2_data_n4031,
PE0_act_regs_1_data_n4035,
PE0_act_regs_0_data_n4039,
PE0_act_regs_3_data_n4048,
PE0_act_regs_2_data_n4052,
PE0_act_regs_1_data_n4056,
PE0_act_regs_0_data_n4060,
PE0_act_regs_3_data_n4068,
PE0_act_regs_2_data_n4072,
PE0_act_regs_1_data_n4076,
PE0_act_regs_0_data_n4080,
PE0_act_regs_3_data_n4092,
PE0_act_regs_2_data_n4096,
PE0_act_regs_1_data_n4100,
PE0_act_regs_0_data_n4104,
PE0_act_regs_3_data_n4112,
PE0_act_regs_2_data_n4116,
PE0_act_regs_1_data_n4120,
PE0_act_regs_0_data_n4124,
PE0_act_regs_3_data_n4136,
PE0_act_regs_2_data_n4140,
PE0_act_regs_1_data_n4144,
PE0_act_regs_0_data_n4148,
PE0_act_regs_3_data_n4160,
PE0_act_regs_2_data_n4164,
PE0_act_regs_1_data_n4168,
PE0_act_regs_0_data_n4172,
PE0_act_regs_3_data_n4184,
PE0_act_regs_2_data_n4188,
PE0_act_regs_1_data_n4192,
PE0_act_regs_0_data_n4196,
PE0_act_regs_3_data_n4208,
PE0_act_regs_2_data_n4212,
PE0_act_regs_1_data_n4216,
PE0_act_regs_0_data_n4220,
pe0_act_buffer_data_n4232,
PE0_act_regs_3_data_n4240,
PE0_act_regs_2_data_n4244,
PE0_act_regs_1_data_n4248,
PE0_act_regs_0_data_n4252,
PE0_act_regs_3_data_n4261,
PE0_act_regs_2_data_n4265,
PE0_act_regs_1_data_n4269,
PE0_act_regs_0_data_n4273,
PE0_act_regs_3_data_n4281,
PE0_act_regs_2_data_n4285,
PE0_act_regs_1_data_n4289,
PE0_act_regs_0_data_n4293,
PE0_act_regs_3_data_n4305,
PE0_act_regs_2_data_n4309,
PE0_act_regs_1_data_n4313,
PE0_act_regs_0_data_n4317,
PE0_act_regs_3_data_n4325,
PE0_act_regs_2_data_n4329,
PE0_act_regs_1_data_n4333,
PE0_act_regs_0_data_n4337,
PE0_act_regs_3_data_n4349,
PE0_act_regs_2_data_n4353,
PE0_act_regs_1_data_n4357,
PE0_act_regs_0_data_n4361,
PE0_act_regs_3_data_n4373,
PE0_act_regs_2_data_n4377,
PE0_act_regs_1_data_n4381,
PE0_act_regs_0_data_n4385,
PE0_act_regs_3_data_n4397,
PE0_act_regs_2_data_n4401,
PE0_act_regs_1_data_n4405,
PE0_act_regs_0_data_n4409,
PE0_act_regs_3_data_n4421,
PE0_act_regs_2_data_n4425,
PE0_act_regs_1_data_n4429,
PE0_act_regs_0_data_n4433,
pe0_act_buffer_addr0,
pe0_act_buffer_data0,
pe0_act_buffer_wen0,
pe0_act_buffer_addr1,
pe0_act_buffer_data1,
pe0_act_buffer_wen1,
pe0_act_buffer_addr2,
pe0_act_buffer_data2,
pe0_act_buffer_wen2,
pe0_act_buffer_addr3,
pe0_act_buffer_data3,
pe0_act_buffer_wen3,
pe0_act_buffer_addr4,
pe0_act_buffer_data4,
pe0_act_buffer_wen4,
pe0_act_buffer_addr5,
pe0_act_buffer_data5,
pe0_act_buffer_wen5,
pe0_act_buffer_addr6,
pe0_act_buffer_data6,
pe0_act_buffer_wen6,
pe0_act_buffer_addr7,
pe0_act_buffer_data7,
pe0_act_buffer_wen7,
pe0_act_buffer_addr8,
pe0_act_buffer_data8,
pe0_act_buffer_wen8,
pe0_act_buffer_addr9,
pe0_act_buffer_data9,
pe0_act_buffer_wen9,
pe0_act_buffer_addr10,
pe0_act_buffer_data10,
pe0_act_buffer_wen10,
pe0_act_buffer_addr11,
pe0_act_buffer_data11,
pe0_act_buffer_wen11,
pe0_act_buffer_addr12,
pe0_act_buffer_data12,
pe0_act_buffer_wen12,
pe0_act_buffer_addr13,
pe0_act_buffer_data13,
pe0_act_buffer_wen13,
pe0_act_buffer_addr14,
pe0_act_buffer_data14,
pe0_act_buffer_wen14,
pe0_act_buffer_addr15,
pe0_act_buffer_data15,
pe0_act_buffer_wen15,
PE0_act_regs_3_addr_n404,
PE0_act_regs_2_addr_n408,
PE0_act_regs_1_addr_n412,
PE0_act_regs_0_addr_n416,
PE0_act_regs_3_addr_n431,
PE0_act_regs_2_addr_n435,
PE0_act_regs_1_addr_n439,
PE0_act_regs_0_addr_n443,
PE0_act_regs_3_addr_n456,
PE0_act_regs_2_addr_n460,
PE0_act_regs_1_addr_n464,
PE0_act_regs_0_addr_n468,
PE0_act_regs_3_addr_n481,
PE0_act_regs_2_addr_n485,
PE0_act_regs_1_addr_n489,
PE0_act_regs_0_addr_n493,
PE0_act_regs_3_addr_n506,
PE0_act_regs_2_addr_n510,
PE0_act_regs_1_addr_n514,
PE0_act_regs_0_addr_n518,
PE0_act_regs_3_addr_n531,
PE0_act_regs_2_addr_n535,
PE0_act_regs_1_addr_n539,
PE0_act_regs_0_addr_n543,
PE0_act_regs_3_addr_n556,
PE0_act_regs_2_addr_n560,
PE0_act_regs_1_addr_n564,
PE0_act_regs_0_addr_n568,
PE0_act_regs_3_addr_n581,
PE0_act_regs_2_addr_n585,
PE0_act_regs_1_addr_n589,
PE0_act_regs_0_addr_n593,
PE0_act_regs_3_addr_n606,
PE0_act_regs_2_addr_n610,
PE0_act_regs_1_addr_n614,
PE0_act_regs_0_addr_n618,
PE0_act_regs_3_addr_n632,
PE0_act_regs_2_addr_n636,
PE0_act_regs_1_addr_n640,
PE0_act_regs_0_addr_n644,
PE0_act_regs_3_addr_n658,
PE0_act_regs_2_addr_n662,
PE0_act_regs_1_addr_n666,
PE0_act_regs_0_addr_n670,
PE0_act_regs_3_addr_n683,
PE0_act_regs_2_addr_n687,
PE0_act_regs_1_addr_n691,
PE0_act_regs_0_addr_n695,
PE0_act_regs_3_addr_n708,
PE0_act_regs_2_addr_n712,
PE0_act_regs_1_addr_n716,
PE0_act_regs_0_addr_n720,
PE0_act_regs_3_addr_n733,
PE0_act_regs_2_addr_n737,
PE0_act_regs_1_addr_n741,
PE0_act_regs_0_addr_n745,
PE0_act_regs_3_addr_n758,
PE0_act_regs_2_addr_n762,
PE0_act_regs_1_addr_n766,
PE0_act_regs_0_addr_n770,
PE0_act_regs_3_addr_n783,
PE0_act_regs_2_addr_n787,
PE0_act_regs_1_addr_n791,
PE0_act_regs_0_addr_n795,
PE0_act_regs_0_addr0,
PE0_act_regs_0_data0,
PE0_act_regs_0_wen0,
PE0_act_regs_0_addr1,
PE0_act_regs_0_data1,
PE0_act_regs_0_wen1,
PE0_act_regs_0_addr2,
PE0_act_regs_0_data2,
PE0_act_regs_0_wen2,
PE0_act_regs_0_addr3,
PE0_act_regs_0_data3,
PE0_act_regs_0_wen3,
PE0_act_regs_0_addr4,
PE0_act_regs_0_data4,
PE0_act_regs_0_wen4,
PE0_act_regs_0_addr5,
PE0_act_regs_0_data5,
PE0_act_regs_0_wen5,
PE0_act_regs_0_addr6,
PE0_act_regs_0_data6,
PE0_act_regs_0_wen6,
PE0_act_regs_0_addr7,
PE0_act_regs_0_data7,
PE0_act_regs_0_wen7,
PE0_act_regs_0_addr8,
PE0_act_regs_0_data8,
PE0_act_regs_0_wen8,
PE0_act_regs_0_addr9,
PE0_act_regs_0_data9,
PE0_act_regs_0_wen9,
PE0_act_regs_0_addr10,
PE0_act_regs_0_data10,
PE0_act_regs_0_wen10,
PE0_act_regs_0_addr11,
PE0_act_regs_0_data11,
PE0_act_regs_0_wen11,
PE0_act_regs_0_addr12,
PE0_act_regs_0_data12,
PE0_act_regs_0_wen12,
PE0_act_regs_0_addr13,
PE0_act_regs_0_data13,
PE0_act_regs_0_wen13,
PE0_act_regs_0_addr14,
PE0_act_regs_0_data14,
PE0_act_regs_0_wen14,
PE0_act_regs_0_addr15,
PE0_act_regs_0_data15,
PE0_act_regs_0_wen15,
PE0_act_regs_1_addr0,
PE0_act_regs_1_data0,
PE0_act_regs_1_wen0,
PE0_act_regs_1_addr1,
PE0_act_regs_1_data1,
PE0_act_regs_1_wen1,
PE0_act_regs_1_addr2,
PE0_act_regs_1_data2,
PE0_act_regs_1_wen2,
PE0_act_regs_1_addr3,
PE0_act_regs_1_data3,
PE0_act_regs_1_wen3,
PE0_act_regs_1_addr4,
PE0_act_regs_1_data4,
PE0_act_regs_1_wen4,
PE0_act_regs_1_addr5,
PE0_act_regs_1_data5,
PE0_act_regs_1_wen5,
PE0_act_regs_1_addr6,
PE0_act_regs_1_data6,
PE0_act_regs_1_wen6,
PE0_act_regs_1_addr7,
PE0_act_regs_1_data7,
PE0_act_regs_1_wen7,
PE0_act_regs_1_addr8,
PE0_act_regs_1_data8,
PE0_act_regs_1_wen8,
PE0_act_regs_1_addr9,
PE0_act_regs_1_data9,
PE0_act_regs_1_wen9,
PE0_act_regs_1_addr10,
PE0_act_regs_1_data10,
PE0_act_regs_1_wen10,
PE0_act_regs_1_addr11,
PE0_act_regs_1_data11,
PE0_act_regs_1_wen11,
PE0_act_regs_1_addr12,
PE0_act_regs_1_data12,
PE0_act_regs_1_wen12,
PE0_act_regs_1_addr13,
PE0_act_regs_1_data13,
PE0_act_regs_1_wen13,
PE0_act_regs_1_addr14,
PE0_act_regs_1_data14,
PE0_act_regs_1_wen14,
PE0_act_regs_1_addr15,
PE0_act_regs_1_data15,
PE0_act_regs_1_wen15,
PE0_act_regs_2_addr0,
PE0_act_regs_2_data0,
PE0_act_regs_2_wen0,
PE0_act_regs_2_addr1,
PE0_act_regs_2_data1,
PE0_act_regs_2_wen1,
PE0_act_regs_2_addr2,
PE0_act_regs_2_data2,
PE0_act_regs_2_wen2,
PE0_act_regs_2_addr3,
PE0_act_regs_2_data3,
PE0_act_regs_2_wen3,
PE0_act_regs_2_addr4,
PE0_act_regs_2_data4,
PE0_act_regs_2_wen4,
PE0_act_regs_2_addr5,
PE0_act_regs_2_data5,
PE0_act_regs_2_wen5,
PE0_act_regs_2_addr6,
PE0_act_regs_2_data6,
PE0_act_regs_2_wen6,
PE0_act_regs_2_addr7,
PE0_act_regs_2_data7,
PE0_act_regs_2_wen7,
PE0_act_regs_2_addr8,
PE0_act_regs_2_data8,
PE0_act_regs_2_wen8,
PE0_act_regs_2_addr9,
PE0_act_regs_2_data9,
PE0_act_regs_2_wen9,
PE0_act_regs_2_addr10,
PE0_act_regs_2_data10,
PE0_act_regs_2_wen10,
PE0_act_regs_2_addr11,
PE0_act_regs_2_data11,
PE0_act_regs_2_wen11,
PE0_act_regs_2_addr12,
PE0_act_regs_2_data12,
PE0_act_regs_2_wen12,
PE0_act_regs_2_addr13,
PE0_act_regs_2_data13,
PE0_act_regs_2_wen13,
PE0_act_regs_2_addr14,
PE0_act_regs_2_data14,
PE0_act_regs_2_wen14,
PE0_act_regs_2_addr15,
PE0_act_regs_2_data15,
PE0_act_regs_2_wen15,
PE0_act_regs_3_addr0,
PE0_act_regs_3_data0,
PE0_act_regs_3_wen0,
PE0_act_regs_3_addr1,
PE0_act_regs_3_data1,
PE0_act_regs_3_wen1,
PE0_act_regs_3_addr2,
PE0_act_regs_3_data2,
PE0_act_regs_3_wen2,
PE0_act_regs_3_addr3,
PE0_act_regs_3_data3,
PE0_act_regs_3_wen3,
PE0_act_regs_3_addr4,
PE0_act_regs_3_data4,
PE0_act_regs_3_wen4,
PE0_act_regs_3_addr5,
PE0_act_regs_3_data5,
PE0_act_regs_3_wen5,
PE0_act_regs_3_addr6,
PE0_act_regs_3_data6,
PE0_act_regs_3_wen6,
PE0_act_regs_3_addr7,
PE0_act_regs_3_data7,
PE0_act_regs_3_wen7,
PE0_act_regs_3_addr8,
PE0_act_regs_3_data8,
PE0_act_regs_3_wen8,
PE0_act_regs_3_addr9,
PE0_act_regs_3_data9,
PE0_act_regs_3_wen9,
PE0_act_regs_3_addr10,
PE0_act_regs_3_data10,
PE0_act_regs_3_wen10,
PE0_act_regs_3_addr11,
PE0_act_regs_3_data11,
PE0_act_regs_3_wen11,
PE0_act_regs_3_addr12,
PE0_act_regs_3_data12,
PE0_act_regs_3_wen12,
PE0_act_regs_3_addr13,
PE0_act_regs_3_data13,
PE0_act_regs_3_wen13,
PE0_act_regs_3_addr14,
PE0_act_regs_3_data14,
PE0_act_regs_3_wen14,
PE0_act_regs_3_addr15,
PE0_act_regs_3_data15,
PE0_act_regs_3_wen15,
pe0_act_buffer_addr_n1035,
PE0_act_regs_3_addr_n1044,
PE0_act_regs_2_addr_n1048,
PE0_act_regs_1_addr_n1052,
PE0_act_regs_0_addr_n1056,
PE0_act_regs_3_addr_n1065,
PE0_act_regs_2_addr_n1069,
PE0_act_regs_1_addr_n1073,
PE0_act_regs_0_addr_n1077,
PE0_act_regs_3_addr_n1085,
PE0_act_regs_2_addr_n1089,
PE0_act_regs_1_addr_n1093,
PE0_act_regs_0_addr_n1097,
PE0_act_regs_3_addr_n1109,
PE0_act_regs_2_addr_n1113,
PE0_act_regs_1_addr_n1117,
PE0_act_regs_0_addr_n1121,
PE0_act_regs_3_addr_n1129,
PE0_act_regs_2_addr_n1133,
PE0_act_regs_1_addr_n1137,
PE0_act_regs_0_addr_n1141,
PE0_act_regs_3_addr_n1153,
PE0_act_regs_2_addr_n1157,
PE0_act_regs_1_addr_n1161,
PE0_act_regs_0_addr_n1165,
PE0_act_regs_3_addr_n1177,
PE0_act_regs_2_addr_n1181,
PE0_act_regs_1_addr_n1185,
PE0_act_regs_0_addr_n1189,
PE0_act_regs_3_addr_n1201,
PE0_act_regs_2_addr_n1205,
PE0_act_regs_1_addr_n1209,
PE0_act_regs_0_addr_n1213,
PE0_act_regs_3_addr_n1225,
PE0_act_regs_2_addr_n1229,
PE0_act_regs_1_addr_n1233,
PE0_act_regs_0_addr_n1237,
pe0_act_buffer_addr_n1249,
PE0_act_regs_3_addr_n1257,
PE0_act_regs_2_addr_n1261,
PE0_act_regs_1_addr_n1265,
PE0_act_regs_0_addr_n1269,
PE0_act_regs_3_addr_n1278,
PE0_act_regs_2_addr_n1282,
PE0_act_regs_1_addr_n1286,
PE0_act_regs_0_addr_n1290,
PE0_act_regs_3_addr_n1298,
PE0_act_regs_2_addr_n1302,
PE0_act_regs_1_addr_n1306,
PE0_act_regs_0_addr_n1310,
PE0_act_regs_3_addr_n1322,
PE0_act_regs_2_addr_n1326,
PE0_act_regs_1_addr_n1330,
PE0_act_regs_0_addr_n1334,
PE0_act_regs_3_addr_n1342,
PE0_act_regs_2_addr_n1346,
PE0_act_regs_1_addr_n1350,
PE0_act_regs_0_addr_n1354,
PE0_act_regs_3_addr_n1366,
PE0_act_regs_2_addr_n1370,
PE0_act_regs_1_addr_n1374,
PE0_act_regs_0_addr_n1378,
PE0_act_regs_3_addr_n1390,
PE0_act_regs_2_addr_n1394,
PE0_act_regs_1_addr_n1398,
PE0_act_regs_0_addr_n1402,
PE0_act_regs_3_addr_n1414,
PE0_act_regs_2_addr_n1418,
PE0_act_regs_1_addr_n1422,
PE0_act_regs_0_addr_n1426,
PE0_act_regs_3_addr_n1438,
PE0_act_regs_2_addr_n1442,
PE0_act_regs_1_addr_n1446,
PE0_act_regs_0_addr_n1450,
pe0_act_buffer_addr_n1462,
PE0_act_regs_3_addr_n1470,
PE0_act_regs_2_addr_n1474,
PE0_act_regs_1_addr_n1478,
PE0_act_regs_0_addr_n1482,
PE0_act_regs_3_addr_n1491,
PE0_act_regs_2_addr_n1495,
PE0_act_regs_1_addr_n1499,
PE0_act_regs_0_addr_n1503,
PE0_act_regs_3_addr_n1511,
PE0_act_regs_2_addr_n1515,
PE0_act_regs_1_addr_n1519,
PE0_act_regs_0_addr_n1523,
PE0_act_regs_3_addr_n1535,
PE0_act_regs_2_addr_n1539,
PE0_act_regs_1_addr_n1543,
PE0_act_regs_0_addr_n1547,
PE0_act_regs_3_addr_n1555,
PE0_act_regs_2_addr_n1559,
PE0_act_regs_1_addr_n1563,
PE0_act_regs_0_addr_n1567,
PE0_act_regs_3_addr_n1579,
PE0_act_regs_2_addr_n1583,
PE0_act_regs_1_addr_n1587,
PE0_act_regs_0_addr_n1591,
PE0_act_regs_3_addr_n1603,
PE0_act_regs_2_addr_n1607,
PE0_act_regs_1_addr_n1611,
PE0_act_regs_0_addr_n1615,
PE0_act_regs_3_addr_n1627,
PE0_act_regs_2_addr_n1631,
PE0_act_regs_1_addr_n1635,
PE0_act_regs_0_addr_n1639,
PE0_act_regs_3_addr_n1651,
PE0_act_regs_2_addr_n1655,
PE0_act_regs_1_addr_n1659,
PE0_act_regs_0_addr_n1663,
pe0_act_buffer_addr_n1675,
PE0_act_regs_3_addr_n1683,
PE0_act_regs_2_addr_n1687,
PE0_act_regs_1_addr_n1691,
PE0_act_regs_0_addr_n1695,
PE0_act_regs_3_addr_n1704,
PE0_act_regs_2_addr_n1708,
PE0_act_regs_1_addr_n1712,
PE0_act_regs_0_addr_n1716,
PE0_act_regs_3_addr_n1724,
PE0_act_regs_2_addr_n1728,
PE0_act_regs_1_addr_n1732,
PE0_act_regs_0_addr_n1736,
PE0_act_regs_3_addr_n1748,
PE0_act_regs_2_addr_n1752,
PE0_act_regs_1_addr_n1756,
PE0_act_regs_0_addr_n1760,
PE0_act_regs_3_addr_n1768,
PE0_act_regs_2_addr_n1772,
PE0_act_regs_1_addr_n1776,
PE0_act_regs_0_addr_n1780,
PE0_act_regs_3_addr_n1792,
PE0_act_regs_2_addr_n1796,
PE0_act_regs_1_addr_n1800,
PE0_act_regs_0_addr_n1804,
PE0_act_regs_3_addr_n1816,
PE0_act_regs_2_addr_n1820,
PE0_act_regs_1_addr_n1824,
PE0_act_regs_0_addr_n1828,
PE0_act_regs_3_addr_n1840,
PE0_act_regs_2_addr_n1844,
PE0_act_regs_1_addr_n1848,
PE0_act_regs_0_addr_n1852,
PE0_act_regs_3_addr_n1864,
PE0_act_regs_2_addr_n1868,
PE0_act_regs_1_addr_n1872,
PE0_act_regs_0_addr_n1876,
pe0_act_buffer_addr_n1888,
PE0_act_regs_3_addr_n1896,
PE0_act_regs_2_addr_n1900,
PE0_act_regs_1_addr_n1904,
PE0_act_regs_0_addr_n1908,
PE0_act_regs_3_addr_n1917,
PE0_act_regs_2_addr_n1921,
PE0_act_regs_1_addr_n1925,
PE0_act_regs_0_addr_n1929,
PE0_act_regs_3_addr_n1937,
PE0_act_regs_2_addr_n1941,
PE0_act_regs_1_addr_n1945,
PE0_act_regs_0_addr_n1949,
PE0_act_regs_3_addr_n1961,
PE0_act_regs_2_addr_n1965,
PE0_act_regs_1_addr_n1969,
PE0_act_regs_0_addr_n1973,
PE0_act_regs_3_addr_n1981,
PE0_act_regs_2_addr_n1985,
PE0_act_regs_1_addr_n1989,
PE0_act_regs_0_addr_n1993,
PE0_act_regs_3_addr_n2005,
PE0_act_regs_2_addr_n2009,
PE0_act_regs_1_addr_n2013,
PE0_act_regs_0_addr_n2017,
PE0_act_regs_3_addr_n2029,
PE0_act_regs_2_addr_n2033,
PE0_act_regs_1_addr_n2037,
PE0_act_regs_0_addr_n2041,
PE0_act_regs_3_addr_n2053,
PE0_act_regs_2_addr_n2057,
PE0_act_regs_1_addr_n2061,
PE0_act_regs_0_addr_n2065,
PE0_act_regs_3_addr_n2077,
PE0_act_regs_2_addr_n2081,
PE0_act_regs_1_addr_n2085,
PE0_act_regs_0_addr_n2089,
pe0_act_buffer_addr_n2101,
PE0_act_regs_3_addr_n2109,
PE0_act_regs_2_addr_n2113,
PE0_act_regs_1_addr_n2117,
PE0_act_regs_0_addr_n2121,
PE0_act_regs_3_addr_n2130,
PE0_act_regs_2_addr_n2134,
PE0_act_regs_1_addr_n2138,
PE0_act_regs_0_addr_n2142,
PE0_act_regs_3_addr_n2150,
PE0_act_regs_2_addr_n2154,
PE0_act_regs_1_addr_n2158,
PE0_act_regs_0_addr_n2162,
PE0_act_regs_3_addr_n2174,
PE0_act_regs_2_addr_n2178,
PE0_act_regs_1_addr_n2182,
PE0_act_regs_0_addr_n2186,
PE0_act_regs_3_addr_n2194,
PE0_act_regs_2_addr_n2198,
PE0_act_regs_1_addr_n2202,
PE0_act_regs_0_addr_n2206,
PE0_act_regs_3_addr_n2218,
PE0_act_regs_2_addr_n2222,
PE0_act_regs_1_addr_n2226,
PE0_act_regs_0_addr_n2230,
PE0_act_regs_3_addr_n2242,
PE0_act_regs_2_addr_n2246,
PE0_act_regs_1_addr_n2250,
PE0_act_regs_0_addr_n2254,
PE0_act_regs_3_addr_n2266,
PE0_act_regs_2_addr_n2270,
PE0_act_regs_1_addr_n2274,
PE0_act_regs_0_addr_n2278,
PE0_act_regs_3_addr_n2290,
PE0_act_regs_2_addr_n2294,
PE0_act_regs_1_addr_n2298,
PE0_act_regs_0_addr_n2302,
pe0_act_buffer_addr_n2314,
PE0_act_regs_3_addr_n2322,
PE0_act_regs_2_addr_n2326,
PE0_act_regs_1_addr_n2330,
PE0_act_regs_0_addr_n2334,
PE0_act_regs_3_addr_n2343,
PE0_act_regs_2_addr_n2347,
PE0_act_regs_1_addr_n2351,
PE0_act_regs_0_addr_n2355,
PE0_act_regs_3_addr_n2363,
PE0_act_regs_2_addr_n2367,
PE0_act_regs_1_addr_n2371,
PE0_act_regs_0_addr_n2375,
PE0_act_regs_3_addr_n2387,
PE0_act_regs_2_addr_n2391,
PE0_act_regs_1_addr_n2395,
PE0_act_regs_0_addr_n2399,
PE0_act_regs_3_addr_n2407,
PE0_act_regs_2_addr_n2411,
PE0_act_regs_1_addr_n2415,
PE0_act_regs_0_addr_n2419,
PE0_act_regs_3_addr_n2431,
PE0_act_regs_2_addr_n2435,
PE0_act_regs_1_addr_n2439,
PE0_act_regs_0_addr_n2443,
PE0_act_regs_3_addr_n2455,
PE0_act_regs_2_addr_n2459,
PE0_act_regs_1_addr_n2463,
PE0_act_regs_0_addr_n2467,
PE0_act_regs_3_addr_n2479,
PE0_act_regs_2_addr_n2483,
PE0_act_regs_1_addr_n2487,
PE0_act_regs_0_addr_n2491,
PE0_act_regs_3_addr_n2503,
PE0_act_regs_2_addr_n2507,
PE0_act_regs_1_addr_n2511,
PE0_act_regs_0_addr_n2515,
pe0_act_buffer_addr_n2527,
PE0_act_regs_3_addr_n2535,
PE0_act_regs_2_addr_n2539,
PE0_act_regs_1_addr_n2543,
PE0_act_regs_0_addr_n2547,
PE0_act_regs_3_addr_n2556,
PE0_act_regs_2_addr_n2560,
PE0_act_regs_1_addr_n2564,
PE0_act_regs_0_addr_n2568,
PE0_act_regs_3_addr_n2576,
PE0_act_regs_2_addr_n2580,
PE0_act_regs_1_addr_n2584,
PE0_act_regs_0_addr_n2588,
PE0_act_regs_3_addr_n2600,
PE0_act_regs_2_addr_n2604,
PE0_act_regs_1_addr_n2608,
PE0_act_regs_0_addr_n2612,
PE0_act_regs_3_addr_n2620,
PE0_act_regs_2_addr_n2624,
PE0_act_regs_1_addr_n2628,
PE0_act_regs_0_addr_n2632,
PE0_act_regs_3_addr_n2644,
PE0_act_regs_2_addr_n2648,
PE0_act_regs_1_addr_n2652,
PE0_act_regs_0_addr_n2656,
PE0_act_regs_3_addr_n2668,
PE0_act_regs_2_addr_n2672,
PE0_act_regs_1_addr_n2676,
PE0_act_regs_0_addr_n2680,
PE0_act_regs_3_addr_n2692,
PE0_act_regs_2_addr_n2696,
PE0_act_regs_1_addr_n2700,
PE0_act_regs_0_addr_n2704,
PE0_act_regs_3_addr_n2716,
PE0_act_regs_2_addr_n2720,
PE0_act_regs_1_addr_n2724,
PE0_act_regs_0_addr_n2728,
pe0_act_buffer_addr_n2740,
PE0_act_regs_3_addr_n2748,
PE0_act_regs_2_addr_n2752,
PE0_act_regs_1_addr_n2756,
PE0_act_regs_0_addr_n2760,
PE0_act_regs_3_addr_n2769,
PE0_act_regs_2_addr_n2773,
PE0_act_regs_1_addr_n2777,
PE0_act_regs_0_addr_n2781,
PE0_act_regs_3_addr_n2789,
PE0_act_regs_2_addr_n2793,
PE0_act_regs_1_addr_n2797,
PE0_act_regs_0_addr_n2801,
PE0_act_regs_3_addr_n2813,
PE0_act_regs_2_addr_n2817,
PE0_act_regs_1_addr_n2821,
PE0_act_regs_0_addr_n2825,
PE0_act_regs_3_addr_n2833,
PE0_act_regs_2_addr_n2837,
PE0_act_regs_1_addr_n2841,
PE0_act_regs_0_addr_n2845,
PE0_act_regs_3_addr_n2857,
PE0_act_regs_2_addr_n2861,
PE0_act_regs_1_addr_n2865,
PE0_act_regs_0_addr_n2869,
PE0_act_regs_3_addr_n2881,
PE0_act_regs_2_addr_n2885,
PE0_act_regs_1_addr_n2889,
PE0_act_regs_0_addr_n2893,
PE0_act_regs_3_addr_n2905,
PE0_act_regs_2_addr_n2909,
PE0_act_regs_1_addr_n2913,
PE0_act_regs_0_addr_n2917,
PE0_act_regs_3_addr_n2929,
PE0_act_regs_2_addr_n2933,
PE0_act_regs_1_addr_n2937,
PE0_act_regs_0_addr_n2941,
pe0_act_buffer_addr_n2953,
PE0_act_regs_3_addr_n2961,
PE0_act_regs_2_addr_n2965,
PE0_act_regs_1_addr_n2969,
PE0_act_regs_0_addr_n2973,
PE0_act_regs_3_addr_n2982,
PE0_act_regs_2_addr_n2986,
PE0_act_regs_1_addr_n2990,
PE0_act_regs_0_addr_n2994,
PE0_act_regs_3_addr_n3002,
PE0_act_regs_2_addr_n3006,
PE0_act_regs_1_addr_n3010,
PE0_act_regs_0_addr_n3014,
PE0_act_regs_3_addr_n3026,
PE0_act_regs_2_addr_n3030,
PE0_act_regs_1_addr_n3034,
PE0_act_regs_0_addr_n3038,
PE0_act_regs_3_addr_n3046,
PE0_act_regs_2_addr_n3050,
PE0_act_regs_1_addr_n3054,
PE0_act_regs_0_addr_n3058,
PE0_act_regs_3_addr_n3070,
PE0_act_regs_2_addr_n3074,
PE0_act_regs_1_addr_n3078,
PE0_act_regs_0_addr_n3082,
PE0_act_regs_3_addr_n3094,
PE0_act_regs_2_addr_n3098,
PE0_act_regs_1_addr_n3102,
PE0_act_regs_0_addr_n3106,
PE0_act_regs_3_addr_n3118,
PE0_act_regs_2_addr_n3122,
PE0_act_regs_1_addr_n3126,
PE0_act_regs_0_addr_n3130,
PE0_act_regs_3_addr_n3142,
PE0_act_regs_2_addr_n3146,
PE0_act_regs_1_addr_n3150,
PE0_act_regs_0_addr_n3154,
pe0_act_buffer_addr_n3166,
PE0_act_regs_3_addr_n3174,
PE0_act_regs_2_addr_n3178,
PE0_act_regs_1_addr_n3182,
PE0_act_regs_0_addr_n3186,
PE0_act_regs_3_addr_n3195,
PE0_act_regs_2_addr_n3199,
PE0_act_regs_1_addr_n3203,
PE0_act_regs_0_addr_n3207,
PE0_act_regs_3_addr_n3215,
PE0_act_regs_2_addr_n3219,
PE0_act_regs_1_addr_n3223,
PE0_act_regs_0_addr_n3227,
PE0_act_regs_3_addr_n3239,
PE0_act_regs_2_addr_n3243,
PE0_act_regs_1_addr_n3247,
PE0_act_regs_0_addr_n3251,
PE0_act_regs_3_addr_n3259,
PE0_act_regs_2_addr_n3263,
PE0_act_regs_1_addr_n3267,
PE0_act_regs_0_addr_n3271,
PE0_act_regs_3_addr_n3283,
PE0_act_regs_2_addr_n3287,
PE0_act_regs_1_addr_n3291,
PE0_act_regs_0_addr_n3295,
PE0_act_regs_3_addr_n3307,
PE0_act_regs_2_addr_n3311,
PE0_act_regs_1_addr_n3315,
PE0_act_regs_0_addr_n3319,
PE0_act_regs_3_addr_n3331,
PE0_act_regs_2_addr_n3335,
PE0_act_regs_1_addr_n3339,
PE0_act_regs_0_addr_n3343,
PE0_act_regs_3_addr_n3355,
PE0_act_regs_2_addr_n3359,
PE0_act_regs_1_addr_n3363,
PE0_act_regs_0_addr_n3367,
pe0_act_buffer_addr_n3379,
PE0_act_regs_3_addr_n3387,
PE0_act_regs_2_addr_n3391,
PE0_act_regs_1_addr_n3395,
PE0_act_regs_0_addr_n3399,
PE0_act_regs_3_addr_n3408,
PE0_act_regs_2_addr_n3412,
PE0_act_regs_1_addr_n3416,
PE0_act_regs_0_addr_n3420,
PE0_act_regs_3_addr_n3428,
PE0_act_regs_2_addr_n3432,
PE0_act_regs_1_addr_n3436,
PE0_act_regs_0_addr_n3440,
PE0_act_regs_3_addr_n3452,
PE0_act_regs_2_addr_n3456,
PE0_act_regs_1_addr_n3460,
PE0_act_regs_0_addr_n3464,
PE0_act_regs_3_addr_n3472,
PE0_act_regs_2_addr_n3476,
PE0_act_regs_1_addr_n3480,
PE0_act_regs_0_addr_n3484,
PE0_act_regs_3_addr_n3496,
PE0_act_regs_2_addr_n3500,
PE0_act_regs_1_addr_n3504,
PE0_act_regs_0_addr_n3508,
PE0_act_regs_3_addr_n3520,
PE0_act_regs_2_addr_n3524,
PE0_act_regs_1_addr_n3528,
PE0_act_regs_0_addr_n3532,
PE0_act_regs_3_addr_n3544,
PE0_act_regs_2_addr_n3548,
PE0_act_regs_1_addr_n3552,
PE0_act_regs_0_addr_n3556,
PE0_act_regs_3_addr_n3568,
PE0_act_regs_2_addr_n3572,
PE0_act_regs_1_addr_n3576,
PE0_act_regs_0_addr_n3580,
pe0_act_buffer_addr_n3592,
PE0_act_regs_3_addr_n3600,
PE0_act_regs_2_addr_n3604,
PE0_act_regs_1_addr_n3608,
PE0_act_regs_0_addr_n3612,
PE0_act_regs_3_addr_n3621,
PE0_act_regs_2_addr_n3625,
PE0_act_regs_1_addr_n3629,
PE0_act_regs_0_addr_n3633,
PE0_act_regs_3_addr_n3641,
PE0_act_regs_2_addr_n3645,
PE0_act_regs_1_addr_n3649,
PE0_act_regs_0_addr_n3653,
PE0_act_regs_3_addr_n3665,
PE0_act_regs_2_addr_n3669,
PE0_act_regs_1_addr_n3673,
PE0_act_regs_0_addr_n3677,
PE0_act_regs_3_addr_n3685,
PE0_act_regs_2_addr_n3689,
PE0_act_regs_1_addr_n3693,
PE0_act_regs_0_addr_n3697,
PE0_act_regs_3_addr_n3709,
PE0_act_regs_2_addr_n3713,
PE0_act_regs_1_addr_n3717,
PE0_act_regs_0_addr_n3721,
PE0_act_regs_3_addr_n3733,
PE0_act_regs_2_addr_n3737,
PE0_act_regs_1_addr_n3741,
PE0_act_regs_0_addr_n3745,
PE0_act_regs_3_addr_n3757,
PE0_act_regs_2_addr_n3761,
PE0_act_regs_1_addr_n3765,
PE0_act_regs_0_addr_n3769,
PE0_act_regs_3_addr_n3781,
PE0_act_regs_2_addr_n3785,
PE0_act_regs_1_addr_n3789,
PE0_act_regs_0_addr_n3793,
pe0_act_buffer_addr_n3805,
PE0_act_regs_3_addr_n3813,
PE0_act_regs_2_addr_n3817,
PE0_act_regs_1_addr_n3821,
PE0_act_regs_0_addr_n3825,
PE0_act_regs_3_addr_n3834,
PE0_act_regs_2_addr_n3838,
PE0_act_regs_1_addr_n3842,
PE0_act_regs_0_addr_n3846,
PE0_act_regs_3_addr_n3854,
PE0_act_regs_2_addr_n3858,
PE0_act_regs_1_addr_n3862,
PE0_act_regs_0_addr_n3866,
PE0_act_regs_3_addr_n3878,
PE0_act_regs_2_addr_n3882,
PE0_act_regs_1_addr_n3886,
PE0_act_regs_0_addr_n3890,
PE0_act_regs_3_addr_n3898,
PE0_act_regs_2_addr_n3902,
PE0_act_regs_1_addr_n3906,
PE0_act_regs_0_addr_n3910,
PE0_act_regs_3_addr_n3922,
PE0_act_regs_2_addr_n3926,
PE0_act_regs_1_addr_n3930,
PE0_act_regs_0_addr_n3934,
PE0_act_regs_3_addr_n3946,
PE0_act_regs_2_addr_n3950,
PE0_act_regs_1_addr_n3954,
PE0_act_regs_0_addr_n3958,
PE0_act_regs_3_addr_n3970,
PE0_act_regs_2_addr_n3974,
PE0_act_regs_1_addr_n3978,
PE0_act_regs_0_addr_n3982,
PE0_act_regs_3_addr_n3994,
PE0_act_regs_2_addr_n3998,
PE0_act_regs_1_addr_n4002,
PE0_act_regs_0_addr_n4006,
pe0_act_buffer_addr_n4018,
PE0_act_regs_3_addr_n4026,
PE0_act_regs_2_addr_n4030,
PE0_act_regs_1_addr_n4034,
PE0_act_regs_0_addr_n4038,
PE0_act_regs_3_addr_n4047,
PE0_act_regs_2_addr_n4051,
PE0_act_regs_1_addr_n4055,
PE0_act_regs_0_addr_n4059,
PE0_act_regs_3_addr_n4067,
PE0_act_regs_2_addr_n4071,
PE0_act_regs_1_addr_n4075,
PE0_act_regs_0_addr_n4079,
PE0_act_regs_3_addr_n4091,
PE0_act_regs_2_addr_n4095,
PE0_act_regs_1_addr_n4099,
PE0_act_regs_0_addr_n4103,
PE0_act_regs_3_addr_n4111,
PE0_act_regs_2_addr_n4115,
PE0_act_regs_1_addr_n4119,
PE0_act_regs_0_addr_n4123,
PE0_act_regs_3_addr_n4135,
PE0_act_regs_2_addr_n4139,
PE0_act_regs_1_addr_n4143,
PE0_act_regs_0_addr_n4147,
PE0_act_regs_3_addr_n4159,
PE0_act_regs_2_addr_n4163,
PE0_act_regs_1_addr_n4167,
PE0_act_regs_0_addr_n4171,
PE0_act_regs_3_addr_n4183,
PE0_act_regs_2_addr_n4187,
PE0_act_regs_1_addr_n4191,
PE0_act_regs_0_addr_n4195,
PE0_act_regs_3_addr_n4207,
PE0_act_regs_2_addr_n4211,
PE0_act_regs_1_addr_n4215,
PE0_act_regs_0_addr_n4219,
pe0_act_buffer_addr_n4231,
PE0_act_regs_3_addr_n4239,
PE0_act_regs_2_addr_n4243,
PE0_act_regs_1_addr_n4247,
PE0_act_regs_0_addr_n4251,
PE0_act_regs_3_addr_n4260,
PE0_act_regs_2_addr_n4264,
PE0_act_regs_1_addr_n4268,
PE0_act_regs_0_addr_n4272,
PE0_act_regs_3_addr_n4280,
PE0_act_regs_2_addr_n4284,
PE0_act_regs_1_addr_n4288,
PE0_act_regs_0_addr_n4292,
PE0_act_regs_3_addr_n4304,
PE0_act_regs_2_addr_n4308,
PE0_act_regs_1_addr_n4312,
PE0_act_regs_0_addr_n4316,
PE0_act_regs_3_addr_n4324,
PE0_act_regs_2_addr_n4328,
PE0_act_regs_1_addr_n4332,
PE0_act_regs_0_addr_n4336,
PE0_act_regs_3_addr_n4348,
PE0_act_regs_2_addr_n4352,
PE0_act_regs_1_addr_n4356,
PE0_act_regs_0_addr_n4360,
PE0_act_regs_3_addr_n4372,
PE0_act_regs_2_addr_n4376,
PE0_act_regs_1_addr_n4380,
PE0_act_regs_0_addr_n4384,
PE0_act_regs_3_addr_n4396,
PE0_act_regs_2_addr_n4400,
PE0_act_regs_1_addr_n4404,
PE0_act_regs_0_addr_n4408,
PE0_act_regs_3_addr_n4420,
PE0_act_regs_2_addr_n4424,
PE0_act_regs_1_addr_n4428,
PE0_act_regs_0_addr_n4432,
rva_in_ready,
act_start_ready,
act_port_ready,
output_port_data,
output_port_addr,
output_port_valid,
done,
done_valid,
pe0_act_mngr_is_valid,
pe0_act_mngr_is_zero_first,
pe0_act_mngr_adpfloat_bias,
pe0_act_mngr_num_inst,
pe0_act_mngr_num_output,
pe0_act_mngr_buffer_addr_base,
pe0_act_mngr_output_addr_base,
act_vector_0_15_Inst_0,
act_vector_0_15_Inst_1,
act_vector_0_15_Inst_2,
act_vector_0_15_Inst_3,
act_vector_0_15_Inst_4,
act_vector_0_15_Inst_5,
act_vector_0_15_Inst_6,
act_vector_0_15_Inst_7,
act_vector_0_15_Inst_8,
act_vector_0_15_Inst_9,
act_vector_0_15_Inst_10,
act_vector_0_15_Inst_11,
act_vector_0_15_Inst_12,
act_vector_0_15_Inst_13,
act_vector_0_15_Inst_14,
act_vector_0_15_Inst_15,
act_vector_16_31_Inst_0,
act_vector_16_31_Inst_1,
act_vector_16_31_Inst_2,
act_vector_16_31_Inst_3,
act_vector_16_31_Inst_4,
act_vector_16_31_Inst_5,
act_vector_16_31_Inst_6,
act_vector_16_31_Inst_7,
act_vector_16_31_Inst_8,
act_vector_16_31_Inst_9,
act_vector_16_31_Inst_10,
act_vector_16_31_Inst_11,
act_vector_16_31_Inst_12,
act_vector_16_31_Inst_13,
act_vector_16_31_Inst_14,
act_vector_16_31_Inst_15,
pe0_act_is_start_reg,
pe0_act_instruction_counter,
pe0_act_output_counter,
pe0_act_state,
PE0_act_reg_temp_0,
PE0_act_reg_temp_1,
PE0_act_reg_temp_2,
PE0_act_reg_temp_3,
PE0_act_reg_temp_4,
PE0_act_reg_temp_5,
PE0_act_reg_temp_6,
PE0_act_reg_temp_7,
PE0_act_reg_temp_8,
PE0_act_reg_temp_9,
PE0_act_reg_temp_10,
PE0_act_reg_temp_11,
PE0_act_reg_temp_12,
PE0_act_reg_temp_13,
PE0_act_reg_temp_14,
PE0_act_reg_temp_15
);
input     [19:0] PE0_core_act_vector_0;
input     [19:0] PE0_core_act_vector_1;
input     [19:0] PE0_core_act_vector_10;
input     [19:0] PE0_core_act_vector_11;
input     [19:0] PE0_core_act_vector_12;
input     [19:0] PE0_core_act_vector_13;
input     [19:0] PE0_core_act_vector_14;
input     [19:0] PE0_core_act_vector_15;
input     [19:0] PE0_core_act_vector_2;
input     [19:0] PE0_core_act_vector_3;
input     [19:0] PE0_core_act_vector_4;
input     [19:0] PE0_core_act_vector_5;
input     [19:0] PE0_core_act_vector_6;
input     [19:0] PE0_core_act_vector_7;
input     [19:0] PE0_core_act_vector_8;
input     [19:0] PE0_core_act_vector_9;
input     [19:0] __ILA_pe_act_grant__;
input            act_start;
input            act_start_valid;
input     [23:0] addr;
input            axi_rw;
input            clk;
input      [7:0] data_in_0;
input      [7:0] data_in_1;
input      [7:0] data_in_10;
input      [7:0] data_in_11;
input      [7:0] data_in_12;
input      [7:0] data_in_13;
input      [7:0] data_in_14;
input      [7:0] data_in_15;
input      [7:0] data_in_2;
input      [7:0] data_in_3;
input      [7:0] data_in_4;
input      [7:0] data_in_5;
input      [7:0] data_in_6;
input      [7:0] data_in_7;
input      [7:0] data_in_8;
input      [7:0] data_in_9;
input            done_ready;
input            output_port_ready;
input            pe0_act_reg_port_valid;
input            rst;
input            rva_in_valid;
input     [15:0] wstrb;
input     [19:0] PE0_act_regs_3_data_n405;
input     [19:0] PE0_act_regs_2_data_n409;
input     [19:0] PE0_act_regs_1_data_n413;
input     [19:0] PE0_act_regs_0_data_n417;
input     [19:0] PE0_act_regs_3_data_n432;
input     [19:0] PE0_act_regs_2_data_n436;
input     [19:0] PE0_act_regs_1_data_n440;
input     [19:0] PE0_act_regs_0_data_n444;
input     [19:0] PE0_act_regs_3_data_n457;
input     [19:0] PE0_act_regs_2_data_n461;
input     [19:0] PE0_act_regs_1_data_n465;
input     [19:0] PE0_act_regs_0_data_n469;
input     [19:0] PE0_act_regs_3_data_n482;
input     [19:0] PE0_act_regs_2_data_n486;
input     [19:0] PE0_act_regs_1_data_n490;
input     [19:0] PE0_act_regs_0_data_n494;
input     [19:0] PE0_act_regs_3_data_n507;
input     [19:0] PE0_act_regs_2_data_n511;
input     [19:0] PE0_act_regs_1_data_n515;
input     [19:0] PE0_act_regs_0_data_n519;
input     [19:0] PE0_act_regs_3_data_n532;
input     [19:0] PE0_act_regs_2_data_n536;
input     [19:0] PE0_act_regs_1_data_n540;
input     [19:0] PE0_act_regs_0_data_n544;
input     [19:0] PE0_act_regs_3_data_n557;
input     [19:0] PE0_act_regs_2_data_n561;
input     [19:0] PE0_act_regs_1_data_n565;
input     [19:0] PE0_act_regs_0_data_n569;
input     [19:0] PE0_act_regs_3_data_n582;
input     [19:0] PE0_act_regs_2_data_n586;
input     [19:0] PE0_act_regs_1_data_n590;
input     [19:0] PE0_act_regs_0_data_n594;
input     [19:0] PE0_act_regs_3_data_n607;
input     [19:0] PE0_act_regs_2_data_n611;
input     [19:0] PE0_act_regs_1_data_n615;
input     [19:0] PE0_act_regs_0_data_n619;
input     [19:0] PE0_act_regs_3_data_n633;
input     [19:0] PE0_act_regs_2_data_n637;
input     [19:0] PE0_act_regs_1_data_n641;
input     [19:0] PE0_act_regs_0_data_n645;
input     [19:0] PE0_act_regs_3_data_n659;
input     [19:0] PE0_act_regs_2_data_n663;
input     [19:0] PE0_act_regs_1_data_n667;
input     [19:0] PE0_act_regs_0_data_n671;
input     [19:0] PE0_act_regs_3_data_n684;
input     [19:0] PE0_act_regs_2_data_n688;
input     [19:0] PE0_act_regs_1_data_n692;
input     [19:0] PE0_act_regs_0_data_n696;
input     [19:0] PE0_act_regs_3_data_n709;
input     [19:0] PE0_act_regs_2_data_n713;
input     [19:0] PE0_act_regs_1_data_n717;
input     [19:0] PE0_act_regs_0_data_n721;
input     [19:0] PE0_act_regs_3_data_n734;
input     [19:0] PE0_act_regs_2_data_n738;
input     [19:0] PE0_act_regs_1_data_n742;
input     [19:0] PE0_act_regs_0_data_n746;
input     [19:0] PE0_act_regs_3_data_n759;
input     [19:0] PE0_act_regs_2_data_n763;
input     [19:0] PE0_act_regs_1_data_n767;
input     [19:0] PE0_act_regs_0_data_n771;
input     [19:0] PE0_act_regs_3_data_n784;
input     [19:0] PE0_act_regs_2_data_n788;
input     [19:0] PE0_act_regs_1_data_n792;
input     [19:0] PE0_act_regs_0_data_n796;
input      [7:0] pe0_act_buffer_data_n1036;
input     [19:0] PE0_act_regs_3_data_n1045;
input     [19:0] PE0_act_regs_2_data_n1049;
input     [19:0] PE0_act_regs_1_data_n1053;
input     [19:0] PE0_act_regs_0_data_n1057;
input     [19:0] PE0_act_regs_3_data_n1066;
input     [19:0] PE0_act_regs_2_data_n1070;
input     [19:0] PE0_act_regs_1_data_n1074;
input     [19:0] PE0_act_regs_0_data_n1078;
input     [19:0] PE0_act_regs_3_data_n1086;
input     [19:0] PE0_act_regs_2_data_n1090;
input     [19:0] PE0_act_regs_1_data_n1094;
input     [19:0] PE0_act_regs_0_data_n1098;
input     [19:0] PE0_act_regs_3_data_n1110;
input     [19:0] PE0_act_regs_2_data_n1114;
input     [19:0] PE0_act_regs_1_data_n1118;
input     [19:0] PE0_act_regs_0_data_n1122;
input     [19:0] PE0_act_regs_3_data_n1130;
input     [19:0] PE0_act_regs_2_data_n1134;
input     [19:0] PE0_act_regs_1_data_n1138;
input     [19:0] PE0_act_regs_0_data_n1142;
input     [19:0] PE0_act_regs_3_data_n1154;
input     [19:0] PE0_act_regs_2_data_n1158;
input     [19:0] PE0_act_regs_1_data_n1162;
input     [19:0] PE0_act_regs_0_data_n1166;
input     [19:0] PE0_act_regs_3_data_n1178;
input     [19:0] PE0_act_regs_2_data_n1182;
input     [19:0] PE0_act_regs_1_data_n1186;
input     [19:0] PE0_act_regs_0_data_n1190;
input     [19:0] PE0_act_regs_3_data_n1202;
input     [19:0] PE0_act_regs_2_data_n1206;
input     [19:0] PE0_act_regs_1_data_n1210;
input     [19:0] PE0_act_regs_0_data_n1214;
input     [19:0] PE0_act_regs_3_data_n1226;
input     [19:0] PE0_act_regs_2_data_n1230;
input     [19:0] PE0_act_regs_1_data_n1234;
input     [19:0] PE0_act_regs_0_data_n1238;
input      [7:0] pe0_act_buffer_data_n1250;
input     [19:0] PE0_act_regs_3_data_n1258;
input     [19:0] PE0_act_regs_2_data_n1262;
input     [19:0] PE0_act_regs_1_data_n1266;
input     [19:0] PE0_act_regs_0_data_n1270;
input     [19:0] PE0_act_regs_3_data_n1279;
input     [19:0] PE0_act_regs_2_data_n1283;
input     [19:0] PE0_act_regs_1_data_n1287;
input     [19:0] PE0_act_regs_0_data_n1291;
input     [19:0] PE0_act_regs_3_data_n1299;
input     [19:0] PE0_act_regs_2_data_n1303;
input     [19:0] PE0_act_regs_1_data_n1307;
input     [19:0] PE0_act_regs_0_data_n1311;
input     [19:0] PE0_act_regs_3_data_n1323;
input     [19:0] PE0_act_regs_2_data_n1327;
input     [19:0] PE0_act_regs_1_data_n1331;
input     [19:0] PE0_act_regs_0_data_n1335;
input     [19:0] PE0_act_regs_3_data_n1343;
input     [19:0] PE0_act_regs_2_data_n1347;
input     [19:0] PE0_act_regs_1_data_n1351;
input     [19:0] PE0_act_regs_0_data_n1355;
input     [19:0] PE0_act_regs_3_data_n1367;
input     [19:0] PE0_act_regs_2_data_n1371;
input     [19:0] PE0_act_regs_1_data_n1375;
input     [19:0] PE0_act_regs_0_data_n1379;
input     [19:0] PE0_act_regs_3_data_n1391;
input     [19:0] PE0_act_regs_2_data_n1395;
input     [19:0] PE0_act_regs_1_data_n1399;
input     [19:0] PE0_act_regs_0_data_n1403;
input     [19:0] PE0_act_regs_3_data_n1415;
input     [19:0] PE0_act_regs_2_data_n1419;
input     [19:0] PE0_act_regs_1_data_n1423;
input     [19:0] PE0_act_regs_0_data_n1427;
input     [19:0] PE0_act_regs_3_data_n1439;
input     [19:0] PE0_act_regs_2_data_n1443;
input     [19:0] PE0_act_regs_1_data_n1447;
input     [19:0] PE0_act_regs_0_data_n1451;
input      [7:0] pe0_act_buffer_data_n1463;
input     [19:0] PE0_act_regs_3_data_n1471;
input     [19:0] PE0_act_regs_2_data_n1475;
input     [19:0] PE0_act_regs_1_data_n1479;
input     [19:0] PE0_act_regs_0_data_n1483;
input     [19:0] PE0_act_regs_3_data_n1492;
input     [19:0] PE0_act_regs_2_data_n1496;
input     [19:0] PE0_act_regs_1_data_n1500;
input     [19:0] PE0_act_regs_0_data_n1504;
input     [19:0] PE0_act_regs_3_data_n1512;
input     [19:0] PE0_act_regs_2_data_n1516;
input     [19:0] PE0_act_regs_1_data_n1520;
input     [19:0] PE0_act_regs_0_data_n1524;
input     [19:0] PE0_act_regs_3_data_n1536;
input     [19:0] PE0_act_regs_2_data_n1540;
input     [19:0] PE0_act_regs_1_data_n1544;
input     [19:0] PE0_act_regs_0_data_n1548;
input     [19:0] PE0_act_regs_3_data_n1556;
input     [19:0] PE0_act_regs_2_data_n1560;
input     [19:0] PE0_act_regs_1_data_n1564;
input     [19:0] PE0_act_regs_0_data_n1568;
input     [19:0] PE0_act_regs_3_data_n1580;
input     [19:0] PE0_act_regs_2_data_n1584;
input     [19:0] PE0_act_regs_1_data_n1588;
input     [19:0] PE0_act_regs_0_data_n1592;
input     [19:0] PE0_act_regs_3_data_n1604;
input     [19:0] PE0_act_regs_2_data_n1608;
input     [19:0] PE0_act_regs_1_data_n1612;
input     [19:0] PE0_act_regs_0_data_n1616;
input     [19:0] PE0_act_regs_3_data_n1628;
input     [19:0] PE0_act_regs_2_data_n1632;
input     [19:0] PE0_act_regs_1_data_n1636;
input     [19:0] PE0_act_regs_0_data_n1640;
input     [19:0] PE0_act_regs_3_data_n1652;
input     [19:0] PE0_act_regs_2_data_n1656;
input     [19:0] PE0_act_regs_1_data_n1660;
input     [19:0] PE0_act_regs_0_data_n1664;
input      [7:0] pe0_act_buffer_data_n1676;
input     [19:0] PE0_act_regs_3_data_n1684;
input     [19:0] PE0_act_regs_2_data_n1688;
input     [19:0] PE0_act_regs_1_data_n1692;
input     [19:0] PE0_act_regs_0_data_n1696;
input     [19:0] PE0_act_regs_3_data_n1705;
input     [19:0] PE0_act_regs_2_data_n1709;
input     [19:0] PE0_act_regs_1_data_n1713;
input     [19:0] PE0_act_regs_0_data_n1717;
input     [19:0] PE0_act_regs_3_data_n1725;
input     [19:0] PE0_act_regs_2_data_n1729;
input     [19:0] PE0_act_regs_1_data_n1733;
input     [19:0] PE0_act_regs_0_data_n1737;
input     [19:0] PE0_act_regs_3_data_n1749;
input     [19:0] PE0_act_regs_2_data_n1753;
input     [19:0] PE0_act_regs_1_data_n1757;
input     [19:0] PE0_act_regs_0_data_n1761;
input     [19:0] PE0_act_regs_3_data_n1769;
input     [19:0] PE0_act_regs_2_data_n1773;
input     [19:0] PE0_act_regs_1_data_n1777;
input     [19:0] PE0_act_regs_0_data_n1781;
input     [19:0] PE0_act_regs_3_data_n1793;
input     [19:0] PE0_act_regs_2_data_n1797;
input     [19:0] PE0_act_regs_1_data_n1801;
input     [19:0] PE0_act_regs_0_data_n1805;
input     [19:0] PE0_act_regs_3_data_n1817;
input     [19:0] PE0_act_regs_2_data_n1821;
input     [19:0] PE0_act_regs_1_data_n1825;
input     [19:0] PE0_act_regs_0_data_n1829;
input     [19:0] PE0_act_regs_3_data_n1841;
input     [19:0] PE0_act_regs_2_data_n1845;
input     [19:0] PE0_act_regs_1_data_n1849;
input     [19:0] PE0_act_regs_0_data_n1853;
input     [19:0] PE0_act_regs_3_data_n1865;
input     [19:0] PE0_act_regs_2_data_n1869;
input     [19:0] PE0_act_regs_1_data_n1873;
input     [19:0] PE0_act_regs_0_data_n1877;
input      [7:0] pe0_act_buffer_data_n1889;
input     [19:0] PE0_act_regs_3_data_n1897;
input     [19:0] PE0_act_regs_2_data_n1901;
input     [19:0] PE0_act_regs_1_data_n1905;
input     [19:0] PE0_act_regs_0_data_n1909;
input     [19:0] PE0_act_regs_3_data_n1918;
input     [19:0] PE0_act_regs_2_data_n1922;
input     [19:0] PE0_act_regs_1_data_n1926;
input     [19:0] PE0_act_regs_0_data_n1930;
input     [19:0] PE0_act_regs_3_data_n1938;
input     [19:0] PE0_act_regs_2_data_n1942;
input     [19:0] PE0_act_regs_1_data_n1946;
input     [19:0] PE0_act_regs_0_data_n1950;
input     [19:0] PE0_act_regs_3_data_n1962;
input     [19:0] PE0_act_regs_2_data_n1966;
input     [19:0] PE0_act_regs_1_data_n1970;
input     [19:0] PE0_act_regs_0_data_n1974;
input     [19:0] PE0_act_regs_3_data_n1982;
input     [19:0] PE0_act_regs_2_data_n1986;
input     [19:0] PE0_act_regs_1_data_n1990;
input     [19:0] PE0_act_regs_0_data_n1994;
input     [19:0] PE0_act_regs_3_data_n2006;
input     [19:0] PE0_act_regs_2_data_n2010;
input     [19:0] PE0_act_regs_1_data_n2014;
input     [19:0] PE0_act_regs_0_data_n2018;
input     [19:0] PE0_act_regs_3_data_n2030;
input     [19:0] PE0_act_regs_2_data_n2034;
input     [19:0] PE0_act_regs_1_data_n2038;
input     [19:0] PE0_act_regs_0_data_n2042;
input     [19:0] PE0_act_regs_3_data_n2054;
input     [19:0] PE0_act_regs_2_data_n2058;
input     [19:0] PE0_act_regs_1_data_n2062;
input     [19:0] PE0_act_regs_0_data_n2066;
input     [19:0] PE0_act_regs_3_data_n2078;
input     [19:0] PE0_act_regs_2_data_n2082;
input     [19:0] PE0_act_regs_1_data_n2086;
input     [19:0] PE0_act_regs_0_data_n2090;
input      [7:0] pe0_act_buffer_data_n2102;
input     [19:0] PE0_act_regs_3_data_n2110;
input     [19:0] PE0_act_regs_2_data_n2114;
input     [19:0] PE0_act_regs_1_data_n2118;
input     [19:0] PE0_act_regs_0_data_n2122;
input     [19:0] PE0_act_regs_3_data_n2131;
input     [19:0] PE0_act_regs_2_data_n2135;
input     [19:0] PE0_act_regs_1_data_n2139;
input     [19:0] PE0_act_regs_0_data_n2143;
input     [19:0] PE0_act_regs_3_data_n2151;
input     [19:0] PE0_act_regs_2_data_n2155;
input     [19:0] PE0_act_regs_1_data_n2159;
input     [19:0] PE0_act_regs_0_data_n2163;
input     [19:0] PE0_act_regs_3_data_n2175;
input     [19:0] PE0_act_regs_2_data_n2179;
input     [19:0] PE0_act_regs_1_data_n2183;
input     [19:0] PE0_act_regs_0_data_n2187;
input     [19:0] PE0_act_regs_3_data_n2195;
input     [19:0] PE0_act_regs_2_data_n2199;
input     [19:0] PE0_act_regs_1_data_n2203;
input     [19:0] PE0_act_regs_0_data_n2207;
input     [19:0] PE0_act_regs_3_data_n2219;
input     [19:0] PE0_act_regs_2_data_n2223;
input     [19:0] PE0_act_regs_1_data_n2227;
input     [19:0] PE0_act_regs_0_data_n2231;
input     [19:0] PE0_act_regs_3_data_n2243;
input     [19:0] PE0_act_regs_2_data_n2247;
input     [19:0] PE0_act_regs_1_data_n2251;
input     [19:0] PE0_act_regs_0_data_n2255;
input     [19:0] PE0_act_regs_3_data_n2267;
input     [19:0] PE0_act_regs_2_data_n2271;
input     [19:0] PE0_act_regs_1_data_n2275;
input     [19:0] PE0_act_regs_0_data_n2279;
input     [19:0] PE0_act_regs_3_data_n2291;
input     [19:0] PE0_act_regs_2_data_n2295;
input     [19:0] PE0_act_regs_1_data_n2299;
input     [19:0] PE0_act_regs_0_data_n2303;
input      [7:0] pe0_act_buffer_data_n2315;
input     [19:0] PE0_act_regs_3_data_n2323;
input     [19:0] PE0_act_regs_2_data_n2327;
input     [19:0] PE0_act_regs_1_data_n2331;
input     [19:0] PE0_act_regs_0_data_n2335;
input     [19:0] PE0_act_regs_3_data_n2344;
input     [19:0] PE0_act_regs_2_data_n2348;
input     [19:0] PE0_act_regs_1_data_n2352;
input     [19:0] PE0_act_regs_0_data_n2356;
input     [19:0] PE0_act_regs_3_data_n2364;
input     [19:0] PE0_act_regs_2_data_n2368;
input     [19:0] PE0_act_regs_1_data_n2372;
input     [19:0] PE0_act_regs_0_data_n2376;
input     [19:0] PE0_act_regs_3_data_n2388;
input     [19:0] PE0_act_regs_2_data_n2392;
input     [19:0] PE0_act_regs_1_data_n2396;
input     [19:0] PE0_act_regs_0_data_n2400;
input     [19:0] PE0_act_regs_3_data_n2408;
input     [19:0] PE0_act_regs_2_data_n2412;
input     [19:0] PE0_act_regs_1_data_n2416;
input     [19:0] PE0_act_regs_0_data_n2420;
input     [19:0] PE0_act_regs_3_data_n2432;
input     [19:0] PE0_act_regs_2_data_n2436;
input     [19:0] PE0_act_regs_1_data_n2440;
input     [19:0] PE0_act_regs_0_data_n2444;
input     [19:0] PE0_act_regs_3_data_n2456;
input     [19:0] PE0_act_regs_2_data_n2460;
input     [19:0] PE0_act_regs_1_data_n2464;
input     [19:0] PE0_act_regs_0_data_n2468;
input     [19:0] PE0_act_regs_3_data_n2480;
input     [19:0] PE0_act_regs_2_data_n2484;
input     [19:0] PE0_act_regs_1_data_n2488;
input     [19:0] PE0_act_regs_0_data_n2492;
input     [19:0] PE0_act_regs_3_data_n2504;
input     [19:0] PE0_act_regs_2_data_n2508;
input     [19:0] PE0_act_regs_1_data_n2512;
input     [19:0] PE0_act_regs_0_data_n2516;
input      [7:0] pe0_act_buffer_data_n2528;
input     [19:0] PE0_act_regs_3_data_n2536;
input     [19:0] PE0_act_regs_2_data_n2540;
input     [19:0] PE0_act_regs_1_data_n2544;
input     [19:0] PE0_act_regs_0_data_n2548;
input     [19:0] PE0_act_regs_3_data_n2557;
input     [19:0] PE0_act_regs_2_data_n2561;
input     [19:0] PE0_act_regs_1_data_n2565;
input     [19:0] PE0_act_regs_0_data_n2569;
input     [19:0] PE0_act_regs_3_data_n2577;
input     [19:0] PE0_act_regs_2_data_n2581;
input     [19:0] PE0_act_regs_1_data_n2585;
input     [19:0] PE0_act_regs_0_data_n2589;
input     [19:0] PE0_act_regs_3_data_n2601;
input     [19:0] PE0_act_regs_2_data_n2605;
input     [19:0] PE0_act_regs_1_data_n2609;
input     [19:0] PE0_act_regs_0_data_n2613;
input     [19:0] PE0_act_regs_3_data_n2621;
input     [19:0] PE0_act_regs_2_data_n2625;
input     [19:0] PE0_act_regs_1_data_n2629;
input     [19:0] PE0_act_regs_0_data_n2633;
input     [19:0] PE0_act_regs_3_data_n2645;
input     [19:0] PE0_act_regs_2_data_n2649;
input     [19:0] PE0_act_regs_1_data_n2653;
input     [19:0] PE0_act_regs_0_data_n2657;
input     [19:0] PE0_act_regs_3_data_n2669;
input     [19:0] PE0_act_regs_2_data_n2673;
input     [19:0] PE0_act_regs_1_data_n2677;
input     [19:0] PE0_act_regs_0_data_n2681;
input     [19:0] PE0_act_regs_3_data_n2693;
input     [19:0] PE0_act_regs_2_data_n2697;
input     [19:0] PE0_act_regs_1_data_n2701;
input     [19:0] PE0_act_regs_0_data_n2705;
input     [19:0] PE0_act_regs_3_data_n2717;
input     [19:0] PE0_act_regs_2_data_n2721;
input     [19:0] PE0_act_regs_1_data_n2725;
input     [19:0] PE0_act_regs_0_data_n2729;
input      [7:0] pe0_act_buffer_data_n2741;
input     [19:0] PE0_act_regs_3_data_n2749;
input     [19:0] PE0_act_regs_2_data_n2753;
input     [19:0] PE0_act_regs_1_data_n2757;
input     [19:0] PE0_act_regs_0_data_n2761;
input     [19:0] PE0_act_regs_3_data_n2770;
input     [19:0] PE0_act_regs_2_data_n2774;
input     [19:0] PE0_act_regs_1_data_n2778;
input     [19:0] PE0_act_regs_0_data_n2782;
input     [19:0] PE0_act_regs_3_data_n2790;
input     [19:0] PE0_act_regs_2_data_n2794;
input     [19:0] PE0_act_regs_1_data_n2798;
input     [19:0] PE0_act_regs_0_data_n2802;
input     [19:0] PE0_act_regs_3_data_n2814;
input     [19:0] PE0_act_regs_2_data_n2818;
input     [19:0] PE0_act_regs_1_data_n2822;
input     [19:0] PE0_act_regs_0_data_n2826;
input     [19:0] PE0_act_regs_3_data_n2834;
input     [19:0] PE0_act_regs_2_data_n2838;
input     [19:0] PE0_act_regs_1_data_n2842;
input     [19:0] PE0_act_regs_0_data_n2846;
input     [19:0] PE0_act_regs_3_data_n2858;
input     [19:0] PE0_act_regs_2_data_n2862;
input     [19:0] PE0_act_regs_1_data_n2866;
input     [19:0] PE0_act_regs_0_data_n2870;
input     [19:0] PE0_act_regs_3_data_n2882;
input     [19:0] PE0_act_regs_2_data_n2886;
input     [19:0] PE0_act_regs_1_data_n2890;
input     [19:0] PE0_act_regs_0_data_n2894;
input     [19:0] PE0_act_regs_3_data_n2906;
input     [19:0] PE0_act_regs_2_data_n2910;
input     [19:0] PE0_act_regs_1_data_n2914;
input     [19:0] PE0_act_regs_0_data_n2918;
input     [19:0] PE0_act_regs_3_data_n2930;
input     [19:0] PE0_act_regs_2_data_n2934;
input     [19:0] PE0_act_regs_1_data_n2938;
input     [19:0] PE0_act_regs_0_data_n2942;
input      [7:0] pe0_act_buffer_data_n2954;
input     [19:0] PE0_act_regs_3_data_n2962;
input     [19:0] PE0_act_regs_2_data_n2966;
input     [19:0] PE0_act_regs_1_data_n2970;
input     [19:0] PE0_act_regs_0_data_n2974;
input     [19:0] PE0_act_regs_3_data_n2983;
input     [19:0] PE0_act_regs_2_data_n2987;
input     [19:0] PE0_act_regs_1_data_n2991;
input     [19:0] PE0_act_regs_0_data_n2995;
input     [19:0] PE0_act_regs_3_data_n3003;
input     [19:0] PE0_act_regs_2_data_n3007;
input     [19:0] PE0_act_regs_1_data_n3011;
input     [19:0] PE0_act_regs_0_data_n3015;
input     [19:0] PE0_act_regs_3_data_n3027;
input     [19:0] PE0_act_regs_2_data_n3031;
input     [19:0] PE0_act_regs_1_data_n3035;
input     [19:0] PE0_act_regs_0_data_n3039;
input     [19:0] PE0_act_regs_3_data_n3047;
input     [19:0] PE0_act_regs_2_data_n3051;
input     [19:0] PE0_act_regs_1_data_n3055;
input     [19:0] PE0_act_regs_0_data_n3059;
input     [19:0] PE0_act_regs_3_data_n3071;
input     [19:0] PE0_act_regs_2_data_n3075;
input     [19:0] PE0_act_regs_1_data_n3079;
input     [19:0] PE0_act_regs_0_data_n3083;
input     [19:0] PE0_act_regs_3_data_n3095;
input     [19:0] PE0_act_regs_2_data_n3099;
input     [19:0] PE0_act_regs_1_data_n3103;
input     [19:0] PE0_act_regs_0_data_n3107;
input     [19:0] PE0_act_regs_3_data_n3119;
input     [19:0] PE0_act_regs_2_data_n3123;
input     [19:0] PE0_act_regs_1_data_n3127;
input     [19:0] PE0_act_regs_0_data_n3131;
input     [19:0] PE0_act_regs_3_data_n3143;
input     [19:0] PE0_act_regs_2_data_n3147;
input     [19:0] PE0_act_regs_1_data_n3151;
input     [19:0] PE0_act_regs_0_data_n3155;
input      [7:0] pe0_act_buffer_data_n3167;
input     [19:0] PE0_act_regs_3_data_n3175;
input     [19:0] PE0_act_regs_2_data_n3179;
input     [19:0] PE0_act_regs_1_data_n3183;
input     [19:0] PE0_act_regs_0_data_n3187;
input     [19:0] PE0_act_regs_3_data_n3196;
input     [19:0] PE0_act_regs_2_data_n3200;
input     [19:0] PE0_act_regs_1_data_n3204;
input     [19:0] PE0_act_regs_0_data_n3208;
input     [19:0] PE0_act_regs_3_data_n3216;
input     [19:0] PE0_act_regs_2_data_n3220;
input     [19:0] PE0_act_regs_1_data_n3224;
input     [19:0] PE0_act_regs_0_data_n3228;
input     [19:0] PE0_act_regs_3_data_n3240;
input     [19:0] PE0_act_regs_2_data_n3244;
input     [19:0] PE0_act_regs_1_data_n3248;
input     [19:0] PE0_act_regs_0_data_n3252;
input     [19:0] PE0_act_regs_3_data_n3260;
input     [19:0] PE0_act_regs_2_data_n3264;
input     [19:0] PE0_act_regs_1_data_n3268;
input     [19:0] PE0_act_regs_0_data_n3272;
input     [19:0] PE0_act_regs_3_data_n3284;
input     [19:0] PE0_act_regs_2_data_n3288;
input     [19:0] PE0_act_regs_1_data_n3292;
input     [19:0] PE0_act_regs_0_data_n3296;
input     [19:0] PE0_act_regs_3_data_n3308;
input     [19:0] PE0_act_regs_2_data_n3312;
input     [19:0] PE0_act_regs_1_data_n3316;
input     [19:0] PE0_act_regs_0_data_n3320;
input     [19:0] PE0_act_regs_3_data_n3332;
input     [19:0] PE0_act_regs_2_data_n3336;
input     [19:0] PE0_act_regs_1_data_n3340;
input     [19:0] PE0_act_regs_0_data_n3344;
input     [19:0] PE0_act_regs_3_data_n3356;
input     [19:0] PE0_act_regs_2_data_n3360;
input     [19:0] PE0_act_regs_1_data_n3364;
input     [19:0] PE0_act_regs_0_data_n3368;
input      [7:0] pe0_act_buffer_data_n3380;
input     [19:0] PE0_act_regs_3_data_n3388;
input     [19:0] PE0_act_regs_2_data_n3392;
input     [19:0] PE0_act_regs_1_data_n3396;
input     [19:0] PE0_act_regs_0_data_n3400;
input     [19:0] PE0_act_regs_3_data_n3409;
input     [19:0] PE0_act_regs_2_data_n3413;
input     [19:0] PE0_act_regs_1_data_n3417;
input     [19:0] PE0_act_regs_0_data_n3421;
input     [19:0] PE0_act_regs_3_data_n3429;
input     [19:0] PE0_act_regs_2_data_n3433;
input     [19:0] PE0_act_regs_1_data_n3437;
input     [19:0] PE0_act_regs_0_data_n3441;
input     [19:0] PE0_act_regs_3_data_n3453;
input     [19:0] PE0_act_regs_2_data_n3457;
input     [19:0] PE0_act_regs_1_data_n3461;
input     [19:0] PE0_act_regs_0_data_n3465;
input     [19:0] PE0_act_regs_3_data_n3473;
input     [19:0] PE0_act_regs_2_data_n3477;
input     [19:0] PE0_act_regs_1_data_n3481;
input     [19:0] PE0_act_regs_0_data_n3485;
input     [19:0] PE0_act_regs_3_data_n3497;
input     [19:0] PE0_act_regs_2_data_n3501;
input     [19:0] PE0_act_regs_1_data_n3505;
input     [19:0] PE0_act_regs_0_data_n3509;
input     [19:0] PE0_act_regs_3_data_n3521;
input     [19:0] PE0_act_regs_2_data_n3525;
input     [19:0] PE0_act_regs_1_data_n3529;
input     [19:0] PE0_act_regs_0_data_n3533;
input     [19:0] PE0_act_regs_3_data_n3545;
input     [19:0] PE0_act_regs_2_data_n3549;
input     [19:0] PE0_act_regs_1_data_n3553;
input     [19:0] PE0_act_regs_0_data_n3557;
input     [19:0] PE0_act_regs_3_data_n3569;
input     [19:0] PE0_act_regs_2_data_n3573;
input     [19:0] PE0_act_regs_1_data_n3577;
input     [19:0] PE0_act_regs_0_data_n3581;
input      [7:0] pe0_act_buffer_data_n3593;
input     [19:0] PE0_act_regs_3_data_n3601;
input     [19:0] PE0_act_regs_2_data_n3605;
input     [19:0] PE0_act_regs_1_data_n3609;
input     [19:0] PE0_act_regs_0_data_n3613;
input     [19:0] PE0_act_regs_3_data_n3622;
input     [19:0] PE0_act_regs_2_data_n3626;
input     [19:0] PE0_act_regs_1_data_n3630;
input     [19:0] PE0_act_regs_0_data_n3634;
input     [19:0] PE0_act_regs_3_data_n3642;
input     [19:0] PE0_act_regs_2_data_n3646;
input     [19:0] PE0_act_regs_1_data_n3650;
input     [19:0] PE0_act_regs_0_data_n3654;
input     [19:0] PE0_act_regs_3_data_n3666;
input     [19:0] PE0_act_regs_2_data_n3670;
input     [19:0] PE0_act_regs_1_data_n3674;
input     [19:0] PE0_act_regs_0_data_n3678;
input     [19:0] PE0_act_regs_3_data_n3686;
input     [19:0] PE0_act_regs_2_data_n3690;
input     [19:0] PE0_act_regs_1_data_n3694;
input     [19:0] PE0_act_regs_0_data_n3698;
input     [19:0] PE0_act_regs_3_data_n3710;
input     [19:0] PE0_act_regs_2_data_n3714;
input     [19:0] PE0_act_regs_1_data_n3718;
input     [19:0] PE0_act_regs_0_data_n3722;
input     [19:0] PE0_act_regs_3_data_n3734;
input     [19:0] PE0_act_regs_2_data_n3738;
input     [19:0] PE0_act_regs_1_data_n3742;
input     [19:0] PE0_act_regs_0_data_n3746;
input     [19:0] PE0_act_regs_3_data_n3758;
input     [19:0] PE0_act_regs_2_data_n3762;
input     [19:0] PE0_act_regs_1_data_n3766;
input     [19:0] PE0_act_regs_0_data_n3770;
input     [19:0] PE0_act_regs_3_data_n3782;
input     [19:0] PE0_act_regs_2_data_n3786;
input     [19:0] PE0_act_regs_1_data_n3790;
input     [19:0] PE0_act_regs_0_data_n3794;
input      [7:0] pe0_act_buffer_data_n3806;
input     [19:0] PE0_act_regs_3_data_n3814;
input     [19:0] PE0_act_regs_2_data_n3818;
input     [19:0] PE0_act_regs_1_data_n3822;
input     [19:0] PE0_act_regs_0_data_n3826;
input     [19:0] PE0_act_regs_3_data_n3835;
input     [19:0] PE0_act_regs_2_data_n3839;
input     [19:0] PE0_act_regs_1_data_n3843;
input     [19:0] PE0_act_regs_0_data_n3847;
input     [19:0] PE0_act_regs_3_data_n3855;
input     [19:0] PE0_act_regs_2_data_n3859;
input     [19:0] PE0_act_regs_1_data_n3863;
input     [19:0] PE0_act_regs_0_data_n3867;
input     [19:0] PE0_act_regs_3_data_n3879;
input     [19:0] PE0_act_regs_2_data_n3883;
input     [19:0] PE0_act_regs_1_data_n3887;
input     [19:0] PE0_act_regs_0_data_n3891;
input     [19:0] PE0_act_regs_3_data_n3899;
input     [19:0] PE0_act_regs_2_data_n3903;
input     [19:0] PE0_act_regs_1_data_n3907;
input     [19:0] PE0_act_regs_0_data_n3911;
input     [19:0] PE0_act_regs_3_data_n3923;
input     [19:0] PE0_act_regs_2_data_n3927;
input     [19:0] PE0_act_regs_1_data_n3931;
input     [19:0] PE0_act_regs_0_data_n3935;
input     [19:0] PE0_act_regs_3_data_n3947;
input     [19:0] PE0_act_regs_2_data_n3951;
input     [19:0] PE0_act_regs_1_data_n3955;
input     [19:0] PE0_act_regs_0_data_n3959;
input     [19:0] PE0_act_regs_3_data_n3971;
input     [19:0] PE0_act_regs_2_data_n3975;
input     [19:0] PE0_act_regs_1_data_n3979;
input     [19:0] PE0_act_regs_0_data_n3983;
input     [19:0] PE0_act_regs_3_data_n3995;
input     [19:0] PE0_act_regs_2_data_n3999;
input     [19:0] PE0_act_regs_1_data_n4003;
input     [19:0] PE0_act_regs_0_data_n4007;
input      [7:0] pe0_act_buffer_data_n4019;
input     [19:0] PE0_act_regs_3_data_n4027;
input     [19:0] PE0_act_regs_2_data_n4031;
input     [19:0] PE0_act_regs_1_data_n4035;
input     [19:0] PE0_act_regs_0_data_n4039;
input     [19:0] PE0_act_regs_3_data_n4048;
input     [19:0] PE0_act_regs_2_data_n4052;
input     [19:0] PE0_act_regs_1_data_n4056;
input     [19:0] PE0_act_regs_0_data_n4060;
input     [19:0] PE0_act_regs_3_data_n4068;
input     [19:0] PE0_act_regs_2_data_n4072;
input     [19:0] PE0_act_regs_1_data_n4076;
input     [19:0] PE0_act_regs_0_data_n4080;
input     [19:0] PE0_act_regs_3_data_n4092;
input     [19:0] PE0_act_regs_2_data_n4096;
input     [19:0] PE0_act_regs_1_data_n4100;
input     [19:0] PE0_act_regs_0_data_n4104;
input     [19:0] PE0_act_regs_3_data_n4112;
input     [19:0] PE0_act_regs_2_data_n4116;
input     [19:0] PE0_act_regs_1_data_n4120;
input     [19:0] PE0_act_regs_0_data_n4124;
input     [19:0] PE0_act_regs_3_data_n4136;
input     [19:0] PE0_act_regs_2_data_n4140;
input     [19:0] PE0_act_regs_1_data_n4144;
input     [19:0] PE0_act_regs_0_data_n4148;
input     [19:0] PE0_act_regs_3_data_n4160;
input     [19:0] PE0_act_regs_2_data_n4164;
input     [19:0] PE0_act_regs_1_data_n4168;
input     [19:0] PE0_act_regs_0_data_n4172;
input     [19:0] PE0_act_regs_3_data_n4184;
input     [19:0] PE0_act_regs_2_data_n4188;
input     [19:0] PE0_act_regs_1_data_n4192;
input     [19:0] PE0_act_regs_0_data_n4196;
input     [19:0] PE0_act_regs_3_data_n4208;
input     [19:0] PE0_act_regs_2_data_n4212;
input     [19:0] PE0_act_regs_1_data_n4216;
input     [19:0] PE0_act_regs_0_data_n4220;
input      [7:0] pe0_act_buffer_data_n4232;
input     [19:0] PE0_act_regs_3_data_n4240;
input     [19:0] PE0_act_regs_2_data_n4244;
input     [19:0] PE0_act_regs_1_data_n4248;
input     [19:0] PE0_act_regs_0_data_n4252;
input     [19:0] PE0_act_regs_3_data_n4261;
input     [19:0] PE0_act_regs_2_data_n4265;
input     [19:0] PE0_act_regs_1_data_n4269;
input     [19:0] PE0_act_regs_0_data_n4273;
input     [19:0] PE0_act_regs_3_data_n4281;
input     [19:0] PE0_act_regs_2_data_n4285;
input     [19:0] PE0_act_regs_1_data_n4289;
input     [19:0] PE0_act_regs_0_data_n4293;
input     [19:0] PE0_act_regs_3_data_n4305;
input     [19:0] PE0_act_regs_2_data_n4309;
input     [19:0] PE0_act_regs_1_data_n4313;
input     [19:0] PE0_act_regs_0_data_n4317;
input     [19:0] PE0_act_regs_3_data_n4325;
input     [19:0] PE0_act_regs_2_data_n4329;
input     [19:0] PE0_act_regs_1_data_n4333;
input     [19:0] PE0_act_regs_0_data_n4337;
input     [19:0] PE0_act_regs_3_data_n4349;
input     [19:0] PE0_act_regs_2_data_n4353;
input     [19:0] PE0_act_regs_1_data_n4357;
input     [19:0] PE0_act_regs_0_data_n4361;
input     [19:0] PE0_act_regs_3_data_n4373;
input     [19:0] PE0_act_regs_2_data_n4377;
input     [19:0] PE0_act_regs_1_data_n4381;
input     [19:0] PE0_act_regs_0_data_n4385;
input     [19:0] PE0_act_regs_3_data_n4397;
input     [19:0] PE0_act_regs_2_data_n4401;
input     [19:0] PE0_act_regs_1_data_n4405;
input     [19:0] PE0_act_regs_0_data_n4409;
input     [19:0] PE0_act_regs_3_data_n4421;
input     [19:0] PE0_act_regs_2_data_n4425;
input     [19:0] PE0_act_regs_1_data_n4429;
input     [19:0] PE0_act_regs_0_data_n4433;
output     [19:0] __ILA_pe_act_acc_decode__;
output            __ILA_pe_act_decode_of_PE0_ACT_STORE_BUFFER__;
output            __ILA_pe_act_decode_of_PE0_CONFIG_ACT_MNGR__;
output            __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_0_15__;
output            __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_16_31__;
output            __ILA_pe_act_decode_of_PE0_act_child_done_sent__;
output            __ILA_pe_act_decode_of_PE0_act_child_initiate__;
output            __ILA_pe_act_decode_of_PE0_act_child_op_copy__;
output            __ILA_pe_act_decode_of_PE0_act_child_op_eadd__;
output            __ILA_pe_act_decode_of_PE0_act_child_op_emul__;
output            __ILA_pe_act_decode_of_PE0_act_child_op_inpe__;
output            __ILA_pe_act_decode_of_PE0_act_child_op_load__;
output            __ILA_pe_act_decode_of_PE0_act_child_op_load_zero__;
output            __ILA_pe_act_decode_of_PE0_act_child_op_onex__;
output            __ILA_pe_act_decode_of_PE0_act_child_op_outgb__;
output            __ILA_pe_act_decode_of_PE0_act_child_op_relu__;
output            __ILA_pe_act_decode_of_PE0_act_child_op_sigm__;
output            __ILA_pe_act_decode_of_PE0_act_child_op_store__;
output            __ILA_pe_act_decode_of_PE0_act_child_op_tanh__;
output            __ILA_pe_act_decode_of_PE0_act_child_out_sent__;
output            __ILA_pe_act_decode_of_PE0_act_child_reg_store__;
output            __ILA_pe_act_valid__;
output     [31:0] pe0_act_buffer_addr0;
output      [7:0] pe0_act_buffer_data0;
output            pe0_act_buffer_wen0;
output     [31:0] pe0_act_buffer_addr1;
output      [7:0] pe0_act_buffer_data1;
output            pe0_act_buffer_wen1;
output     [31:0] pe0_act_buffer_addr2;
output      [7:0] pe0_act_buffer_data2;
output            pe0_act_buffer_wen2;
output     [31:0] pe0_act_buffer_addr3;
output      [7:0] pe0_act_buffer_data3;
output            pe0_act_buffer_wen3;
output     [31:0] pe0_act_buffer_addr4;
output      [7:0] pe0_act_buffer_data4;
output            pe0_act_buffer_wen4;
output     [31:0] pe0_act_buffer_addr5;
output      [7:0] pe0_act_buffer_data5;
output            pe0_act_buffer_wen5;
output     [31:0] pe0_act_buffer_addr6;
output      [7:0] pe0_act_buffer_data6;
output            pe0_act_buffer_wen6;
output     [31:0] pe0_act_buffer_addr7;
output      [7:0] pe0_act_buffer_data7;
output            pe0_act_buffer_wen7;
output     [31:0] pe0_act_buffer_addr8;
output      [7:0] pe0_act_buffer_data8;
output            pe0_act_buffer_wen8;
output     [31:0] pe0_act_buffer_addr9;
output      [7:0] pe0_act_buffer_data9;
output            pe0_act_buffer_wen9;
output     [31:0] pe0_act_buffer_addr10;
output      [7:0] pe0_act_buffer_data10;
output            pe0_act_buffer_wen10;
output     [31:0] pe0_act_buffer_addr11;
output      [7:0] pe0_act_buffer_data11;
output            pe0_act_buffer_wen11;
output     [31:0] pe0_act_buffer_addr12;
output      [7:0] pe0_act_buffer_data12;
output            pe0_act_buffer_wen12;
output     [31:0] pe0_act_buffer_addr13;
output      [7:0] pe0_act_buffer_data13;
output            pe0_act_buffer_wen13;
output     [31:0] pe0_act_buffer_addr14;
output      [7:0] pe0_act_buffer_data14;
output            pe0_act_buffer_wen14;
output     [31:0] pe0_act_buffer_addr15;
output      [7:0] pe0_act_buffer_data15;
output            pe0_act_buffer_wen15;
output      [3:0] PE0_act_regs_3_addr_n404;
output      [3:0] PE0_act_regs_2_addr_n408;
output      [3:0] PE0_act_regs_1_addr_n412;
output      [3:0] PE0_act_regs_0_addr_n416;
output      [3:0] PE0_act_regs_3_addr_n431;
output      [3:0] PE0_act_regs_2_addr_n435;
output      [3:0] PE0_act_regs_1_addr_n439;
output      [3:0] PE0_act_regs_0_addr_n443;
output      [3:0] PE0_act_regs_3_addr_n456;
output      [3:0] PE0_act_regs_2_addr_n460;
output      [3:0] PE0_act_regs_1_addr_n464;
output      [3:0] PE0_act_regs_0_addr_n468;
output      [3:0] PE0_act_regs_3_addr_n481;
output      [3:0] PE0_act_regs_2_addr_n485;
output      [3:0] PE0_act_regs_1_addr_n489;
output      [3:0] PE0_act_regs_0_addr_n493;
output      [3:0] PE0_act_regs_3_addr_n506;
output      [3:0] PE0_act_regs_2_addr_n510;
output      [3:0] PE0_act_regs_1_addr_n514;
output      [3:0] PE0_act_regs_0_addr_n518;
output      [3:0] PE0_act_regs_3_addr_n531;
output      [3:0] PE0_act_regs_2_addr_n535;
output      [3:0] PE0_act_regs_1_addr_n539;
output      [3:0] PE0_act_regs_0_addr_n543;
output      [3:0] PE0_act_regs_3_addr_n556;
output      [3:0] PE0_act_regs_2_addr_n560;
output      [3:0] PE0_act_regs_1_addr_n564;
output      [3:0] PE0_act_regs_0_addr_n568;
output      [3:0] PE0_act_regs_3_addr_n581;
output      [3:0] PE0_act_regs_2_addr_n585;
output      [3:0] PE0_act_regs_1_addr_n589;
output      [3:0] PE0_act_regs_0_addr_n593;
output      [3:0] PE0_act_regs_3_addr_n606;
output      [3:0] PE0_act_regs_2_addr_n610;
output      [3:0] PE0_act_regs_1_addr_n614;
output      [3:0] PE0_act_regs_0_addr_n618;
output      [3:0] PE0_act_regs_3_addr_n632;
output      [3:0] PE0_act_regs_2_addr_n636;
output      [3:0] PE0_act_regs_1_addr_n640;
output      [3:0] PE0_act_regs_0_addr_n644;
output      [3:0] PE0_act_regs_3_addr_n658;
output      [3:0] PE0_act_regs_2_addr_n662;
output      [3:0] PE0_act_regs_1_addr_n666;
output      [3:0] PE0_act_regs_0_addr_n670;
output      [3:0] PE0_act_regs_3_addr_n683;
output      [3:0] PE0_act_regs_2_addr_n687;
output      [3:0] PE0_act_regs_1_addr_n691;
output      [3:0] PE0_act_regs_0_addr_n695;
output      [3:0] PE0_act_regs_3_addr_n708;
output      [3:0] PE0_act_regs_2_addr_n712;
output      [3:0] PE0_act_regs_1_addr_n716;
output      [3:0] PE0_act_regs_0_addr_n720;
output      [3:0] PE0_act_regs_3_addr_n733;
output      [3:0] PE0_act_regs_2_addr_n737;
output      [3:0] PE0_act_regs_1_addr_n741;
output      [3:0] PE0_act_regs_0_addr_n745;
output      [3:0] PE0_act_regs_3_addr_n758;
output      [3:0] PE0_act_regs_2_addr_n762;
output      [3:0] PE0_act_regs_1_addr_n766;
output      [3:0] PE0_act_regs_0_addr_n770;
output      [3:0] PE0_act_regs_3_addr_n783;
output      [3:0] PE0_act_regs_2_addr_n787;
output      [3:0] PE0_act_regs_1_addr_n791;
output      [3:0] PE0_act_regs_0_addr_n795;
output      [3:0] PE0_act_regs_0_addr0;
output     [19:0] PE0_act_regs_0_data0;
output            PE0_act_regs_0_wen0;
output      [3:0] PE0_act_regs_0_addr1;
output     [19:0] PE0_act_regs_0_data1;
output            PE0_act_regs_0_wen1;
output      [3:0] PE0_act_regs_0_addr2;
output     [19:0] PE0_act_regs_0_data2;
output            PE0_act_regs_0_wen2;
output      [3:0] PE0_act_regs_0_addr3;
output     [19:0] PE0_act_regs_0_data3;
output            PE0_act_regs_0_wen3;
output      [3:0] PE0_act_regs_0_addr4;
output     [19:0] PE0_act_regs_0_data4;
output            PE0_act_regs_0_wen4;
output      [3:0] PE0_act_regs_0_addr5;
output     [19:0] PE0_act_regs_0_data5;
output            PE0_act_regs_0_wen5;
output      [3:0] PE0_act_regs_0_addr6;
output     [19:0] PE0_act_regs_0_data6;
output            PE0_act_regs_0_wen6;
output      [3:0] PE0_act_regs_0_addr7;
output     [19:0] PE0_act_regs_0_data7;
output            PE0_act_regs_0_wen7;
output      [3:0] PE0_act_regs_0_addr8;
output     [19:0] PE0_act_regs_0_data8;
output            PE0_act_regs_0_wen8;
output      [3:0] PE0_act_regs_0_addr9;
output     [19:0] PE0_act_regs_0_data9;
output            PE0_act_regs_0_wen9;
output      [3:0] PE0_act_regs_0_addr10;
output     [19:0] PE0_act_regs_0_data10;
output            PE0_act_regs_0_wen10;
output      [3:0] PE0_act_regs_0_addr11;
output     [19:0] PE0_act_regs_0_data11;
output            PE0_act_regs_0_wen11;
output      [3:0] PE0_act_regs_0_addr12;
output     [19:0] PE0_act_regs_0_data12;
output            PE0_act_regs_0_wen12;
output      [3:0] PE0_act_regs_0_addr13;
output     [19:0] PE0_act_regs_0_data13;
output            PE0_act_regs_0_wen13;
output      [3:0] PE0_act_regs_0_addr14;
output     [19:0] PE0_act_regs_0_data14;
output            PE0_act_regs_0_wen14;
output      [3:0] PE0_act_regs_0_addr15;
output     [19:0] PE0_act_regs_0_data15;
output            PE0_act_regs_0_wen15;
output      [3:0] PE0_act_regs_1_addr0;
output     [19:0] PE0_act_regs_1_data0;
output            PE0_act_regs_1_wen0;
output      [3:0] PE0_act_regs_1_addr1;
output     [19:0] PE0_act_regs_1_data1;
output            PE0_act_regs_1_wen1;
output      [3:0] PE0_act_regs_1_addr2;
output     [19:0] PE0_act_regs_1_data2;
output            PE0_act_regs_1_wen2;
output      [3:0] PE0_act_regs_1_addr3;
output     [19:0] PE0_act_regs_1_data3;
output            PE0_act_regs_1_wen3;
output      [3:0] PE0_act_regs_1_addr4;
output     [19:0] PE0_act_regs_1_data4;
output            PE0_act_regs_1_wen4;
output      [3:0] PE0_act_regs_1_addr5;
output     [19:0] PE0_act_regs_1_data5;
output            PE0_act_regs_1_wen5;
output      [3:0] PE0_act_regs_1_addr6;
output     [19:0] PE0_act_regs_1_data6;
output            PE0_act_regs_1_wen6;
output      [3:0] PE0_act_regs_1_addr7;
output     [19:0] PE0_act_regs_1_data7;
output            PE0_act_regs_1_wen7;
output      [3:0] PE0_act_regs_1_addr8;
output     [19:0] PE0_act_regs_1_data8;
output            PE0_act_regs_1_wen8;
output      [3:0] PE0_act_regs_1_addr9;
output     [19:0] PE0_act_regs_1_data9;
output            PE0_act_regs_1_wen9;
output      [3:0] PE0_act_regs_1_addr10;
output     [19:0] PE0_act_regs_1_data10;
output            PE0_act_regs_1_wen10;
output      [3:0] PE0_act_regs_1_addr11;
output     [19:0] PE0_act_regs_1_data11;
output            PE0_act_regs_1_wen11;
output      [3:0] PE0_act_regs_1_addr12;
output     [19:0] PE0_act_regs_1_data12;
output            PE0_act_regs_1_wen12;
output      [3:0] PE0_act_regs_1_addr13;
output     [19:0] PE0_act_regs_1_data13;
output            PE0_act_regs_1_wen13;
output      [3:0] PE0_act_regs_1_addr14;
output     [19:0] PE0_act_regs_1_data14;
output            PE0_act_regs_1_wen14;
output      [3:0] PE0_act_regs_1_addr15;
output     [19:0] PE0_act_regs_1_data15;
output            PE0_act_regs_1_wen15;
output      [3:0] PE0_act_regs_2_addr0;
output     [19:0] PE0_act_regs_2_data0;
output            PE0_act_regs_2_wen0;
output      [3:0] PE0_act_regs_2_addr1;
output     [19:0] PE0_act_regs_2_data1;
output            PE0_act_regs_2_wen1;
output      [3:0] PE0_act_regs_2_addr2;
output     [19:0] PE0_act_regs_2_data2;
output            PE0_act_regs_2_wen2;
output      [3:0] PE0_act_regs_2_addr3;
output     [19:0] PE0_act_regs_2_data3;
output            PE0_act_regs_2_wen3;
output      [3:0] PE0_act_regs_2_addr4;
output     [19:0] PE0_act_regs_2_data4;
output            PE0_act_regs_2_wen4;
output      [3:0] PE0_act_regs_2_addr5;
output     [19:0] PE0_act_regs_2_data5;
output            PE0_act_regs_2_wen5;
output      [3:0] PE0_act_regs_2_addr6;
output     [19:0] PE0_act_regs_2_data6;
output            PE0_act_regs_2_wen6;
output      [3:0] PE0_act_regs_2_addr7;
output     [19:0] PE0_act_regs_2_data7;
output            PE0_act_regs_2_wen7;
output      [3:0] PE0_act_regs_2_addr8;
output     [19:0] PE0_act_regs_2_data8;
output            PE0_act_regs_2_wen8;
output      [3:0] PE0_act_regs_2_addr9;
output     [19:0] PE0_act_regs_2_data9;
output            PE0_act_regs_2_wen9;
output      [3:0] PE0_act_regs_2_addr10;
output     [19:0] PE0_act_regs_2_data10;
output            PE0_act_regs_2_wen10;
output      [3:0] PE0_act_regs_2_addr11;
output     [19:0] PE0_act_regs_2_data11;
output            PE0_act_regs_2_wen11;
output      [3:0] PE0_act_regs_2_addr12;
output     [19:0] PE0_act_regs_2_data12;
output            PE0_act_regs_2_wen12;
output      [3:0] PE0_act_regs_2_addr13;
output     [19:0] PE0_act_regs_2_data13;
output            PE0_act_regs_2_wen13;
output      [3:0] PE0_act_regs_2_addr14;
output     [19:0] PE0_act_regs_2_data14;
output            PE0_act_regs_2_wen14;
output      [3:0] PE0_act_regs_2_addr15;
output     [19:0] PE0_act_regs_2_data15;
output            PE0_act_regs_2_wen15;
output      [3:0] PE0_act_regs_3_addr0;
output     [19:0] PE0_act_regs_3_data0;
output            PE0_act_regs_3_wen0;
output      [3:0] PE0_act_regs_3_addr1;
output     [19:0] PE0_act_regs_3_data1;
output            PE0_act_regs_3_wen1;
output      [3:0] PE0_act_regs_3_addr2;
output     [19:0] PE0_act_regs_3_data2;
output            PE0_act_regs_3_wen2;
output      [3:0] PE0_act_regs_3_addr3;
output     [19:0] PE0_act_regs_3_data3;
output            PE0_act_regs_3_wen3;
output      [3:0] PE0_act_regs_3_addr4;
output     [19:0] PE0_act_regs_3_data4;
output            PE0_act_regs_3_wen4;
output      [3:0] PE0_act_regs_3_addr5;
output     [19:0] PE0_act_regs_3_data5;
output            PE0_act_regs_3_wen5;
output      [3:0] PE0_act_regs_3_addr6;
output     [19:0] PE0_act_regs_3_data6;
output            PE0_act_regs_3_wen6;
output      [3:0] PE0_act_regs_3_addr7;
output     [19:0] PE0_act_regs_3_data7;
output            PE0_act_regs_3_wen7;
output      [3:0] PE0_act_regs_3_addr8;
output     [19:0] PE0_act_regs_3_data8;
output            PE0_act_regs_3_wen8;
output      [3:0] PE0_act_regs_3_addr9;
output     [19:0] PE0_act_regs_3_data9;
output            PE0_act_regs_3_wen9;
output      [3:0] PE0_act_regs_3_addr10;
output     [19:0] PE0_act_regs_3_data10;
output            PE0_act_regs_3_wen10;
output      [3:0] PE0_act_regs_3_addr11;
output     [19:0] PE0_act_regs_3_data11;
output            PE0_act_regs_3_wen11;
output      [3:0] PE0_act_regs_3_addr12;
output     [19:0] PE0_act_regs_3_data12;
output            PE0_act_regs_3_wen12;
output      [3:0] PE0_act_regs_3_addr13;
output     [19:0] PE0_act_regs_3_data13;
output            PE0_act_regs_3_wen13;
output      [3:0] PE0_act_regs_3_addr14;
output     [19:0] PE0_act_regs_3_data14;
output            PE0_act_regs_3_wen14;
output      [3:0] PE0_act_regs_3_addr15;
output     [19:0] PE0_act_regs_3_data15;
output            PE0_act_regs_3_wen15;
output     [31:0] pe0_act_buffer_addr_n1035;
output      [3:0] PE0_act_regs_3_addr_n1044;
output      [3:0] PE0_act_regs_2_addr_n1048;
output      [3:0] PE0_act_regs_1_addr_n1052;
output      [3:0] PE0_act_regs_0_addr_n1056;
output      [3:0] PE0_act_regs_3_addr_n1065;
output      [3:0] PE0_act_regs_2_addr_n1069;
output      [3:0] PE0_act_regs_1_addr_n1073;
output      [3:0] PE0_act_regs_0_addr_n1077;
output      [3:0] PE0_act_regs_3_addr_n1085;
output      [3:0] PE0_act_regs_2_addr_n1089;
output      [3:0] PE0_act_regs_1_addr_n1093;
output      [3:0] PE0_act_regs_0_addr_n1097;
output      [3:0] PE0_act_regs_3_addr_n1109;
output      [3:0] PE0_act_regs_2_addr_n1113;
output      [3:0] PE0_act_regs_1_addr_n1117;
output      [3:0] PE0_act_regs_0_addr_n1121;
output      [3:0] PE0_act_regs_3_addr_n1129;
output      [3:0] PE0_act_regs_2_addr_n1133;
output      [3:0] PE0_act_regs_1_addr_n1137;
output      [3:0] PE0_act_regs_0_addr_n1141;
output      [3:0] PE0_act_regs_3_addr_n1153;
output      [3:0] PE0_act_regs_2_addr_n1157;
output      [3:0] PE0_act_regs_1_addr_n1161;
output      [3:0] PE0_act_regs_0_addr_n1165;
output      [3:0] PE0_act_regs_3_addr_n1177;
output      [3:0] PE0_act_regs_2_addr_n1181;
output      [3:0] PE0_act_regs_1_addr_n1185;
output      [3:0] PE0_act_regs_0_addr_n1189;
output      [3:0] PE0_act_regs_3_addr_n1201;
output      [3:0] PE0_act_regs_2_addr_n1205;
output      [3:0] PE0_act_regs_1_addr_n1209;
output      [3:0] PE0_act_regs_0_addr_n1213;
output      [3:0] PE0_act_regs_3_addr_n1225;
output      [3:0] PE0_act_regs_2_addr_n1229;
output      [3:0] PE0_act_regs_1_addr_n1233;
output      [3:0] PE0_act_regs_0_addr_n1237;
output     [31:0] pe0_act_buffer_addr_n1249;
output      [3:0] PE0_act_regs_3_addr_n1257;
output      [3:0] PE0_act_regs_2_addr_n1261;
output      [3:0] PE0_act_regs_1_addr_n1265;
output      [3:0] PE0_act_regs_0_addr_n1269;
output      [3:0] PE0_act_regs_3_addr_n1278;
output      [3:0] PE0_act_regs_2_addr_n1282;
output      [3:0] PE0_act_regs_1_addr_n1286;
output      [3:0] PE0_act_regs_0_addr_n1290;
output      [3:0] PE0_act_regs_3_addr_n1298;
output      [3:0] PE0_act_regs_2_addr_n1302;
output      [3:0] PE0_act_regs_1_addr_n1306;
output      [3:0] PE0_act_regs_0_addr_n1310;
output      [3:0] PE0_act_regs_3_addr_n1322;
output      [3:0] PE0_act_regs_2_addr_n1326;
output      [3:0] PE0_act_regs_1_addr_n1330;
output      [3:0] PE0_act_regs_0_addr_n1334;
output      [3:0] PE0_act_regs_3_addr_n1342;
output      [3:0] PE0_act_regs_2_addr_n1346;
output      [3:0] PE0_act_regs_1_addr_n1350;
output      [3:0] PE0_act_regs_0_addr_n1354;
output      [3:0] PE0_act_regs_3_addr_n1366;
output      [3:0] PE0_act_regs_2_addr_n1370;
output      [3:0] PE0_act_regs_1_addr_n1374;
output      [3:0] PE0_act_regs_0_addr_n1378;
output      [3:0] PE0_act_regs_3_addr_n1390;
output      [3:0] PE0_act_regs_2_addr_n1394;
output      [3:0] PE0_act_regs_1_addr_n1398;
output      [3:0] PE0_act_regs_0_addr_n1402;
output      [3:0] PE0_act_regs_3_addr_n1414;
output      [3:0] PE0_act_regs_2_addr_n1418;
output      [3:0] PE0_act_regs_1_addr_n1422;
output      [3:0] PE0_act_regs_0_addr_n1426;
output      [3:0] PE0_act_regs_3_addr_n1438;
output      [3:0] PE0_act_regs_2_addr_n1442;
output      [3:0] PE0_act_regs_1_addr_n1446;
output      [3:0] PE0_act_regs_0_addr_n1450;
output     [31:0] pe0_act_buffer_addr_n1462;
output      [3:0] PE0_act_regs_3_addr_n1470;
output      [3:0] PE0_act_regs_2_addr_n1474;
output      [3:0] PE0_act_regs_1_addr_n1478;
output      [3:0] PE0_act_regs_0_addr_n1482;
output      [3:0] PE0_act_regs_3_addr_n1491;
output      [3:0] PE0_act_regs_2_addr_n1495;
output      [3:0] PE0_act_regs_1_addr_n1499;
output      [3:0] PE0_act_regs_0_addr_n1503;
output      [3:0] PE0_act_regs_3_addr_n1511;
output      [3:0] PE0_act_regs_2_addr_n1515;
output      [3:0] PE0_act_regs_1_addr_n1519;
output      [3:0] PE0_act_regs_0_addr_n1523;
output      [3:0] PE0_act_regs_3_addr_n1535;
output      [3:0] PE0_act_regs_2_addr_n1539;
output      [3:0] PE0_act_regs_1_addr_n1543;
output      [3:0] PE0_act_regs_0_addr_n1547;
output      [3:0] PE0_act_regs_3_addr_n1555;
output      [3:0] PE0_act_regs_2_addr_n1559;
output      [3:0] PE0_act_regs_1_addr_n1563;
output      [3:0] PE0_act_regs_0_addr_n1567;
output      [3:0] PE0_act_regs_3_addr_n1579;
output      [3:0] PE0_act_regs_2_addr_n1583;
output      [3:0] PE0_act_regs_1_addr_n1587;
output      [3:0] PE0_act_regs_0_addr_n1591;
output      [3:0] PE0_act_regs_3_addr_n1603;
output      [3:0] PE0_act_regs_2_addr_n1607;
output      [3:0] PE0_act_regs_1_addr_n1611;
output      [3:0] PE0_act_regs_0_addr_n1615;
output      [3:0] PE0_act_regs_3_addr_n1627;
output      [3:0] PE0_act_regs_2_addr_n1631;
output      [3:0] PE0_act_regs_1_addr_n1635;
output      [3:0] PE0_act_regs_0_addr_n1639;
output      [3:0] PE0_act_regs_3_addr_n1651;
output      [3:0] PE0_act_regs_2_addr_n1655;
output      [3:0] PE0_act_regs_1_addr_n1659;
output      [3:0] PE0_act_regs_0_addr_n1663;
output     [31:0] pe0_act_buffer_addr_n1675;
output      [3:0] PE0_act_regs_3_addr_n1683;
output      [3:0] PE0_act_regs_2_addr_n1687;
output      [3:0] PE0_act_regs_1_addr_n1691;
output      [3:0] PE0_act_regs_0_addr_n1695;
output      [3:0] PE0_act_regs_3_addr_n1704;
output      [3:0] PE0_act_regs_2_addr_n1708;
output      [3:0] PE0_act_regs_1_addr_n1712;
output      [3:0] PE0_act_regs_0_addr_n1716;
output      [3:0] PE0_act_regs_3_addr_n1724;
output      [3:0] PE0_act_regs_2_addr_n1728;
output      [3:0] PE0_act_regs_1_addr_n1732;
output      [3:0] PE0_act_regs_0_addr_n1736;
output      [3:0] PE0_act_regs_3_addr_n1748;
output      [3:0] PE0_act_regs_2_addr_n1752;
output      [3:0] PE0_act_regs_1_addr_n1756;
output      [3:0] PE0_act_regs_0_addr_n1760;
output      [3:0] PE0_act_regs_3_addr_n1768;
output      [3:0] PE0_act_regs_2_addr_n1772;
output      [3:0] PE0_act_regs_1_addr_n1776;
output      [3:0] PE0_act_regs_0_addr_n1780;
output      [3:0] PE0_act_regs_3_addr_n1792;
output      [3:0] PE0_act_regs_2_addr_n1796;
output      [3:0] PE0_act_regs_1_addr_n1800;
output      [3:0] PE0_act_regs_0_addr_n1804;
output      [3:0] PE0_act_regs_3_addr_n1816;
output      [3:0] PE0_act_regs_2_addr_n1820;
output      [3:0] PE0_act_regs_1_addr_n1824;
output      [3:0] PE0_act_regs_0_addr_n1828;
output      [3:0] PE0_act_regs_3_addr_n1840;
output      [3:0] PE0_act_regs_2_addr_n1844;
output      [3:0] PE0_act_regs_1_addr_n1848;
output      [3:0] PE0_act_regs_0_addr_n1852;
output      [3:0] PE0_act_regs_3_addr_n1864;
output      [3:0] PE0_act_regs_2_addr_n1868;
output      [3:0] PE0_act_regs_1_addr_n1872;
output      [3:0] PE0_act_regs_0_addr_n1876;
output     [31:0] pe0_act_buffer_addr_n1888;
output      [3:0] PE0_act_regs_3_addr_n1896;
output      [3:0] PE0_act_regs_2_addr_n1900;
output      [3:0] PE0_act_regs_1_addr_n1904;
output      [3:0] PE0_act_regs_0_addr_n1908;
output      [3:0] PE0_act_regs_3_addr_n1917;
output      [3:0] PE0_act_regs_2_addr_n1921;
output      [3:0] PE0_act_regs_1_addr_n1925;
output      [3:0] PE0_act_regs_0_addr_n1929;
output      [3:0] PE0_act_regs_3_addr_n1937;
output      [3:0] PE0_act_regs_2_addr_n1941;
output      [3:0] PE0_act_regs_1_addr_n1945;
output      [3:0] PE0_act_regs_0_addr_n1949;
output      [3:0] PE0_act_regs_3_addr_n1961;
output      [3:0] PE0_act_regs_2_addr_n1965;
output      [3:0] PE0_act_regs_1_addr_n1969;
output      [3:0] PE0_act_regs_0_addr_n1973;
output      [3:0] PE0_act_regs_3_addr_n1981;
output      [3:0] PE0_act_regs_2_addr_n1985;
output      [3:0] PE0_act_regs_1_addr_n1989;
output      [3:0] PE0_act_regs_0_addr_n1993;
output      [3:0] PE0_act_regs_3_addr_n2005;
output      [3:0] PE0_act_regs_2_addr_n2009;
output      [3:0] PE0_act_regs_1_addr_n2013;
output      [3:0] PE0_act_regs_0_addr_n2017;
output      [3:0] PE0_act_regs_3_addr_n2029;
output      [3:0] PE0_act_regs_2_addr_n2033;
output      [3:0] PE0_act_regs_1_addr_n2037;
output      [3:0] PE0_act_regs_0_addr_n2041;
output      [3:0] PE0_act_regs_3_addr_n2053;
output      [3:0] PE0_act_regs_2_addr_n2057;
output      [3:0] PE0_act_regs_1_addr_n2061;
output      [3:0] PE0_act_regs_0_addr_n2065;
output      [3:0] PE0_act_regs_3_addr_n2077;
output      [3:0] PE0_act_regs_2_addr_n2081;
output      [3:0] PE0_act_regs_1_addr_n2085;
output      [3:0] PE0_act_regs_0_addr_n2089;
output     [31:0] pe0_act_buffer_addr_n2101;
output      [3:0] PE0_act_regs_3_addr_n2109;
output      [3:0] PE0_act_regs_2_addr_n2113;
output      [3:0] PE0_act_regs_1_addr_n2117;
output      [3:0] PE0_act_regs_0_addr_n2121;
output      [3:0] PE0_act_regs_3_addr_n2130;
output      [3:0] PE0_act_regs_2_addr_n2134;
output      [3:0] PE0_act_regs_1_addr_n2138;
output      [3:0] PE0_act_regs_0_addr_n2142;
output      [3:0] PE0_act_regs_3_addr_n2150;
output      [3:0] PE0_act_regs_2_addr_n2154;
output      [3:0] PE0_act_regs_1_addr_n2158;
output      [3:0] PE0_act_regs_0_addr_n2162;
output      [3:0] PE0_act_regs_3_addr_n2174;
output      [3:0] PE0_act_regs_2_addr_n2178;
output      [3:0] PE0_act_regs_1_addr_n2182;
output      [3:0] PE0_act_regs_0_addr_n2186;
output      [3:0] PE0_act_regs_3_addr_n2194;
output      [3:0] PE0_act_regs_2_addr_n2198;
output      [3:0] PE0_act_regs_1_addr_n2202;
output      [3:0] PE0_act_regs_0_addr_n2206;
output      [3:0] PE0_act_regs_3_addr_n2218;
output      [3:0] PE0_act_regs_2_addr_n2222;
output      [3:0] PE0_act_regs_1_addr_n2226;
output      [3:0] PE0_act_regs_0_addr_n2230;
output      [3:0] PE0_act_regs_3_addr_n2242;
output      [3:0] PE0_act_regs_2_addr_n2246;
output      [3:0] PE0_act_regs_1_addr_n2250;
output      [3:0] PE0_act_regs_0_addr_n2254;
output      [3:0] PE0_act_regs_3_addr_n2266;
output      [3:0] PE0_act_regs_2_addr_n2270;
output      [3:0] PE0_act_regs_1_addr_n2274;
output      [3:0] PE0_act_regs_0_addr_n2278;
output      [3:0] PE0_act_regs_3_addr_n2290;
output      [3:0] PE0_act_regs_2_addr_n2294;
output      [3:0] PE0_act_regs_1_addr_n2298;
output      [3:0] PE0_act_regs_0_addr_n2302;
output     [31:0] pe0_act_buffer_addr_n2314;
output      [3:0] PE0_act_regs_3_addr_n2322;
output      [3:0] PE0_act_regs_2_addr_n2326;
output      [3:0] PE0_act_regs_1_addr_n2330;
output      [3:0] PE0_act_regs_0_addr_n2334;
output      [3:0] PE0_act_regs_3_addr_n2343;
output      [3:0] PE0_act_regs_2_addr_n2347;
output      [3:0] PE0_act_regs_1_addr_n2351;
output      [3:0] PE0_act_regs_0_addr_n2355;
output      [3:0] PE0_act_regs_3_addr_n2363;
output      [3:0] PE0_act_regs_2_addr_n2367;
output      [3:0] PE0_act_regs_1_addr_n2371;
output      [3:0] PE0_act_regs_0_addr_n2375;
output      [3:0] PE0_act_regs_3_addr_n2387;
output      [3:0] PE0_act_regs_2_addr_n2391;
output      [3:0] PE0_act_regs_1_addr_n2395;
output      [3:0] PE0_act_regs_0_addr_n2399;
output      [3:0] PE0_act_regs_3_addr_n2407;
output      [3:0] PE0_act_regs_2_addr_n2411;
output      [3:0] PE0_act_regs_1_addr_n2415;
output      [3:0] PE0_act_regs_0_addr_n2419;
output      [3:0] PE0_act_regs_3_addr_n2431;
output      [3:0] PE0_act_regs_2_addr_n2435;
output      [3:0] PE0_act_regs_1_addr_n2439;
output      [3:0] PE0_act_regs_0_addr_n2443;
output      [3:0] PE0_act_regs_3_addr_n2455;
output      [3:0] PE0_act_regs_2_addr_n2459;
output      [3:0] PE0_act_regs_1_addr_n2463;
output      [3:0] PE0_act_regs_0_addr_n2467;
output      [3:0] PE0_act_regs_3_addr_n2479;
output      [3:0] PE0_act_regs_2_addr_n2483;
output      [3:0] PE0_act_regs_1_addr_n2487;
output      [3:0] PE0_act_regs_0_addr_n2491;
output      [3:0] PE0_act_regs_3_addr_n2503;
output      [3:0] PE0_act_regs_2_addr_n2507;
output      [3:0] PE0_act_regs_1_addr_n2511;
output      [3:0] PE0_act_regs_0_addr_n2515;
output     [31:0] pe0_act_buffer_addr_n2527;
output      [3:0] PE0_act_regs_3_addr_n2535;
output      [3:0] PE0_act_regs_2_addr_n2539;
output      [3:0] PE0_act_regs_1_addr_n2543;
output      [3:0] PE0_act_regs_0_addr_n2547;
output      [3:0] PE0_act_regs_3_addr_n2556;
output      [3:0] PE0_act_regs_2_addr_n2560;
output      [3:0] PE0_act_regs_1_addr_n2564;
output      [3:0] PE0_act_regs_0_addr_n2568;
output      [3:0] PE0_act_regs_3_addr_n2576;
output      [3:0] PE0_act_regs_2_addr_n2580;
output      [3:0] PE0_act_regs_1_addr_n2584;
output      [3:0] PE0_act_regs_0_addr_n2588;
output      [3:0] PE0_act_regs_3_addr_n2600;
output      [3:0] PE0_act_regs_2_addr_n2604;
output      [3:0] PE0_act_regs_1_addr_n2608;
output      [3:0] PE0_act_regs_0_addr_n2612;
output      [3:0] PE0_act_regs_3_addr_n2620;
output      [3:0] PE0_act_regs_2_addr_n2624;
output      [3:0] PE0_act_regs_1_addr_n2628;
output      [3:0] PE0_act_regs_0_addr_n2632;
output      [3:0] PE0_act_regs_3_addr_n2644;
output      [3:0] PE0_act_regs_2_addr_n2648;
output      [3:0] PE0_act_regs_1_addr_n2652;
output      [3:0] PE0_act_regs_0_addr_n2656;
output      [3:0] PE0_act_regs_3_addr_n2668;
output      [3:0] PE0_act_regs_2_addr_n2672;
output      [3:0] PE0_act_regs_1_addr_n2676;
output      [3:0] PE0_act_regs_0_addr_n2680;
output      [3:0] PE0_act_regs_3_addr_n2692;
output      [3:0] PE0_act_regs_2_addr_n2696;
output      [3:0] PE0_act_regs_1_addr_n2700;
output      [3:0] PE0_act_regs_0_addr_n2704;
output      [3:0] PE0_act_regs_3_addr_n2716;
output      [3:0] PE0_act_regs_2_addr_n2720;
output      [3:0] PE0_act_regs_1_addr_n2724;
output      [3:0] PE0_act_regs_0_addr_n2728;
output     [31:0] pe0_act_buffer_addr_n2740;
output      [3:0] PE0_act_regs_3_addr_n2748;
output      [3:0] PE0_act_regs_2_addr_n2752;
output      [3:0] PE0_act_regs_1_addr_n2756;
output      [3:0] PE0_act_regs_0_addr_n2760;
output      [3:0] PE0_act_regs_3_addr_n2769;
output      [3:0] PE0_act_regs_2_addr_n2773;
output      [3:0] PE0_act_regs_1_addr_n2777;
output      [3:0] PE0_act_regs_0_addr_n2781;
output      [3:0] PE0_act_regs_3_addr_n2789;
output      [3:0] PE0_act_regs_2_addr_n2793;
output      [3:0] PE0_act_regs_1_addr_n2797;
output      [3:0] PE0_act_regs_0_addr_n2801;
output      [3:0] PE0_act_regs_3_addr_n2813;
output      [3:0] PE0_act_regs_2_addr_n2817;
output      [3:0] PE0_act_regs_1_addr_n2821;
output      [3:0] PE0_act_regs_0_addr_n2825;
output      [3:0] PE0_act_regs_3_addr_n2833;
output      [3:0] PE0_act_regs_2_addr_n2837;
output      [3:0] PE0_act_regs_1_addr_n2841;
output      [3:0] PE0_act_regs_0_addr_n2845;
output      [3:0] PE0_act_regs_3_addr_n2857;
output      [3:0] PE0_act_regs_2_addr_n2861;
output      [3:0] PE0_act_regs_1_addr_n2865;
output      [3:0] PE0_act_regs_0_addr_n2869;
output      [3:0] PE0_act_regs_3_addr_n2881;
output      [3:0] PE0_act_regs_2_addr_n2885;
output      [3:0] PE0_act_regs_1_addr_n2889;
output      [3:0] PE0_act_regs_0_addr_n2893;
output      [3:0] PE0_act_regs_3_addr_n2905;
output      [3:0] PE0_act_regs_2_addr_n2909;
output      [3:0] PE0_act_regs_1_addr_n2913;
output      [3:0] PE0_act_regs_0_addr_n2917;
output      [3:0] PE0_act_regs_3_addr_n2929;
output      [3:0] PE0_act_regs_2_addr_n2933;
output      [3:0] PE0_act_regs_1_addr_n2937;
output      [3:0] PE0_act_regs_0_addr_n2941;
output     [31:0] pe0_act_buffer_addr_n2953;
output      [3:0] PE0_act_regs_3_addr_n2961;
output      [3:0] PE0_act_regs_2_addr_n2965;
output      [3:0] PE0_act_regs_1_addr_n2969;
output      [3:0] PE0_act_regs_0_addr_n2973;
output      [3:0] PE0_act_regs_3_addr_n2982;
output      [3:0] PE0_act_regs_2_addr_n2986;
output      [3:0] PE0_act_regs_1_addr_n2990;
output      [3:0] PE0_act_regs_0_addr_n2994;
output      [3:0] PE0_act_regs_3_addr_n3002;
output      [3:0] PE0_act_regs_2_addr_n3006;
output      [3:0] PE0_act_regs_1_addr_n3010;
output      [3:0] PE0_act_regs_0_addr_n3014;
output      [3:0] PE0_act_regs_3_addr_n3026;
output      [3:0] PE0_act_regs_2_addr_n3030;
output      [3:0] PE0_act_regs_1_addr_n3034;
output      [3:0] PE0_act_regs_0_addr_n3038;
output      [3:0] PE0_act_regs_3_addr_n3046;
output      [3:0] PE0_act_regs_2_addr_n3050;
output      [3:0] PE0_act_regs_1_addr_n3054;
output      [3:0] PE0_act_regs_0_addr_n3058;
output      [3:0] PE0_act_regs_3_addr_n3070;
output      [3:0] PE0_act_regs_2_addr_n3074;
output      [3:0] PE0_act_regs_1_addr_n3078;
output      [3:0] PE0_act_regs_0_addr_n3082;
output      [3:0] PE0_act_regs_3_addr_n3094;
output      [3:0] PE0_act_regs_2_addr_n3098;
output      [3:0] PE0_act_regs_1_addr_n3102;
output      [3:0] PE0_act_regs_0_addr_n3106;
output      [3:0] PE0_act_regs_3_addr_n3118;
output      [3:0] PE0_act_regs_2_addr_n3122;
output      [3:0] PE0_act_regs_1_addr_n3126;
output      [3:0] PE0_act_regs_0_addr_n3130;
output      [3:0] PE0_act_regs_3_addr_n3142;
output      [3:0] PE0_act_regs_2_addr_n3146;
output      [3:0] PE0_act_regs_1_addr_n3150;
output      [3:0] PE0_act_regs_0_addr_n3154;
output     [31:0] pe0_act_buffer_addr_n3166;
output      [3:0] PE0_act_regs_3_addr_n3174;
output      [3:0] PE0_act_regs_2_addr_n3178;
output      [3:0] PE0_act_regs_1_addr_n3182;
output      [3:0] PE0_act_regs_0_addr_n3186;
output      [3:0] PE0_act_regs_3_addr_n3195;
output      [3:0] PE0_act_regs_2_addr_n3199;
output      [3:0] PE0_act_regs_1_addr_n3203;
output      [3:0] PE0_act_regs_0_addr_n3207;
output      [3:0] PE0_act_regs_3_addr_n3215;
output      [3:0] PE0_act_regs_2_addr_n3219;
output      [3:0] PE0_act_regs_1_addr_n3223;
output      [3:0] PE0_act_regs_0_addr_n3227;
output      [3:0] PE0_act_regs_3_addr_n3239;
output      [3:0] PE0_act_regs_2_addr_n3243;
output      [3:0] PE0_act_regs_1_addr_n3247;
output      [3:0] PE0_act_regs_0_addr_n3251;
output      [3:0] PE0_act_regs_3_addr_n3259;
output      [3:0] PE0_act_regs_2_addr_n3263;
output      [3:0] PE0_act_regs_1_addr_n3267;
output      [3:0] PE0_act_regs_0_addr_n3271;
output      [3:0] PE0_act_regs_3_addr_n3283;
output      [3:0] PE0_act_regs_2_addr_n3287;
output      [3:0] PE0_act_regs_1_addr_n3291;
output      [3:0] PE0_act_regs_0_addr_n3295;
output      [3:0] PE0_act_regs_3_addr_n3307;
output      [3:0] PE0_act_regs_2_addr_n3311;
output      [3:0] PE0_act_regs_1_addr_n3315;
output      [3:0] PE0_act_regs_0_addr_n3319;
output      [3:0] PE0_act_regs_3_addr_n3331;
output      [3:0] PE0_act_regs_2_addr_n3335;
output      [3:0] PE0_act_regs_1_addr_n3339;
output      [3:0] PE0_act_regs_0_addr_n3343;
output      [3:0] PE0_act_regs_3_addr_n3355;
output      [3:0] PE0_act_regs_2_addr_n3359;
output      [3:0] PE0_act_regs_1_addr_n3363;
output      [3:0] PE0_act_regs_0_addr_n3367;
output     [31:0] pe0_act_buffer_addr_n3379;
output      [3:0] PE0_act_regs_3_addr_n3387;
output      [3:0] PE0_act_regs_2_addr_n3391;
output      [3:0] PE0_act_regs_1_addr_n3395;
output      [3:0] PE0_act_regs_0_addr_n3399;
output      [3:0] PE0_act_regs_3_addr_n3408;
output      [3:0] PE0_act_regs_2_addr_n3412;
output      [3:0] PE0_act_regs_1_addr_n3416;
output      [3:0] PE0_act_regs_0_addr_n3420;
output      [3:0] PE0_act_regs_3_addr_n3428;
output      [3:0] PE0_act_regs_2_addr_n3432;
output      [3:0] PE0_act_regs_1_addr_n3436;
output      [3:0] PE0_act_regs_0_addr_n3440;
output      [3:0] PE0_act_regs_3_addr_n3452;
output      [3:0] PE0_act_regs_2_addr_n3456;
output      [3:0] PE0_act_regs_1_addr_n3460;
output      [3:0] PE0_act_regs_0_addr_n3464;
output      [3:0] PE0_act_regs_3_addr_n3472;
output      [3:0] PE0_act_regs_2_addr_n3476;
output      [3:0] PE0_act_regs_1_addr_n3480;
output      [3:0] PE0_act_regs_0_addr_n3484;
output      [3:0] PE0_act_regs_3_addr_n3496;
output      [3:0] PE0_act_regs_2_addr_n3500;
output      [3:0] PE0_act_regs_1_addr_n3504;
output      [3:0] PE0_act_regs_0_addr_n3508;
output      [3:0] PE0_act_regs_3_addr_n3520;
output      [3:0] PE0_act_regs_2_addr_n3524;
output      [3:0] PE0_act_regs_1_addr_n3528;
output      [3:0] PE0_act_regs_0_addr_n3532;
output      [3:0] PE0_act_regs_3_addr_n3544;
output      [3:0] PE0_act_regs_2_addr_n3548;
output      [3:0] PE0_act_regs_1_addr_n3552;
output      [3:0] PE0_act_regs_0_addr_n3556;
output      [3:0] PE0_act_regs_3_addr_n3568;
output      [3:0] PE0_act_regs_2_addr_n3572;
output      [3:0] PE0_act_regs_1_addr_n3576;
output      [3:0] PE0_act_regs_0_addr_n3580;
output     [31:0] pe0_act_buffer_addr_n3592;
output      [3:0] PE0_act_regs_3_addr_n3600;
output      [3:0] PE0_act_regs_2_addr_n3604;
output      [3:0] PE0_act_regs_1_addr_n3608;
output      [3:0] PE0_act_regs_0_addr_n3612;
output      [3:0] PE0_act_regs_3_addr_n3621;
output      [3:0] PE0_act_regs_2_addr_n3625;
output      [3:0] PE0_act_regs_1_addr_n3629;
output      [3:0] PE0_act_regs_0_addr_n3633;
output      [3:0] PE0_act_regs_3_addr_n3641;
output      [3:0] PE0_act_regs_2_addr_n3645;
output      [3:0] PE0_act_regs_1_addr_n3649;
output      [3:0] PE0_act_regs_0_addr_n3653;
output      [3:0] PE0_act_regs_3_addr_n3665;
output      [3:0] PE0_act_regs_2_addr_n3669;
output      [3:0] PE0_act_regs_1_addr_n3673;
output      [3:0] PE0_act_regs_0_addr_n3677;
output      [3:0] PE0_act_regs_3_addr_n3685;
output      [3:0] PE0_act_regs_2_addr_n3689;
output      [3:0] PE0_act_regs_1_addr_n3693;
output      [3:0] PE0_act_regs_0_addr_n3697;
output      [3:0] PE0_act_regs_3_addr_n3709;
output      [3:0] PE0_act_regs_2_addr_n3713;
output      [3:0] PE0_act_regs_1_addr_n3717;
output      [3:0] PE0_act_regs_0_addr_n3721;
output      [3:0] PE0_act_regs_3_addr_n3733;
output      [3:0] PE0_act_regs_2_addr_n3737;
output      [3:0] PE0_act_regs_1_addr_n3741;
output      [3:0] PE0_act_regs_0_addr_n3745;
output      [3:0] PE0_act_regs_3_addr_n3757;
output      [3:0] PE0_act_regs_2_addr_n3761;
output      [3:0] PE0_act_regs_1_addr_n3765;
output      [3:0] PE0_act_regs_0_addr_n3769;
output      [3:0] PE0_act_regs_3_addr_n3781;
output      [3:0] PE0_act_regs_2_addr_n3785;
output      [3:0] PE0_act_regs_1_addr_n3789;
output      [3:0] PE0_act_regs_0_addr_n3793;
output     [31:0] pe0_act_buffer_addr_n3805;
output      [3:0] PE0_act_regs_3_addr_n3813;
output      [3:0] PE0_act_regs_2_addr_n3817;
output      [3:0] PE0_act_regs_1_addr_n3821;
output      [3:0] PE0_act_regs_0_addr_n3825;
output      [3:0] PE0_act_regs_3_addr_n3834;
output      [3:0] PE0_act_regs_2_addr_n3838;
output      [3:0] PE0_act_regs_1_addr_n3842;
output      [3:0] PE0_act_regs_0_addr_n3846;
output      [3:0] PE0_act_regs_3_addr_n3854;
output      [3:0] PE0_act_regs_2_addr_n3858;
output      [3:0] PE0_act_regs_1_addr_n3862;
output      [3:0] PE0_act_regs_0_addr_n3866;
output      [3:0] PE0_act_regs_3_addr_n3878;
output      [3:0] PE0_act_regs_2_addr_n3882;
output      [3:0] PE0_act_regs_1_addr_n3886;
output      [3:0] PE0_act_regs_0_addr_n3890;
output      [3:0] PE0_act_regs_3_addr_n3898;
output      [3:0] PE0_act_regs_2_addr_n3902;
output      [3:0] PE0_act_regs_1_addr_n3906;
output      [3:0] PE0_act_regs_0_addr_n3910;
output      [3:0] PE0_act_regs_3_addr_n3922;
output      [3:0] PE0_act_regs_2_addr_n3926;
output      [3:0] PE0_act_regs_1_addr_n3930;
output      [3:0] PE0_act_regs_0_addr_n3934;
output      [3:0] PE0_act_regs_3_addr_n3946;
output      [3:0] PE0_act_regs_2_addr_n3950;
output      [3:0] PE0_act_regs_1_addr_n3954;
output      [3:0] PE0_act_regs_0_addr_n3958;
output      [3:0] PE0_act_regs_3_addr_n3970;
output      [3:0] PE0_act_regs_2_addr_n3974;
output      [3:0] PE0_act_regs_1_addr_n3978;
output      [3:0] PE0_act_regs_0_addr_n3982;
output      [3:0] PE0_act_regs_3_addr_n3994;
output      [3:0] PE0_act_regs_2_addr_n3998;
output      [3:0] PE0_act_regs_1_addr_n4002;
output      [3:0] PE0_act_regs_0_addr_n4006;
output     [31:0] pe0_act_buffer_addr_n4018;
output      [3:0] PE0_act_regs_3_addr_n4026;
output      [3:0] PE0_act_regs_2_addr_n4030;
output      [3:0] PE0_act_regs_1_addr_n4034;
output      [3:0] PE0_act_regs_0_addr_n4038;
output      [3:0] PE0_act_regs_3_addr_n4047;
output      [3:0] PE0_act_regs_2_addr_n4051;
output      [3:0] PE0_act_regs_1_addr_n4055;
output      [3:0] PE0_act_regs_0_addr_n4059;
output      [3:0] PE0_act_regs_3_addr_n4067;
output      [3:0] PE0_act_regs_2_addr_n4071;
output      [3:0] PE0_act_regs_1_addr_n4075;
output      [3:0] PE0_act_regs_0_addr_n4079;
output      [3:0] PE0_act_regs_3_addr_n4091;
output      [3:0] PE0_act_regs_2_addr_n4095;
output      [3:0] PE0_act_regs_1_addr_n4099;
output      [3:0] PE0_act_regs_0_addr_n4103;
output      [3:0] PE0_act_regs_3_addr_n4111;
output      [3:0] PE0_act_regs_2_addr_n4115;
output      [3:0] PE0_act_regs_1_addr_n4119;
output      [3:0] PE0_act_regs_0_addr_n4123;
output      [3:0] PE0_act_regs_3_addr_n4135;
output      [3:0] PE0_act_regs_2_addr_n4139;
output      [3:0] PE0_act_regs_1_addr_n4143;
output      [3:0] PE0_act_regs_0_addr_n4147;
output      [3:0] PE0_act_regs_3_addr_n4159;
output      [3:0] PE0_act_regs_2_addr_n4163;
output      [3:0] PE0_act_regs_1_addr_n4167;
output      [3:0] PE0_act_regs_0_addr_n4171;
output      [3:0] PE0_act_regs_3_addr_n4183;
output      [3:0] PE0_act_regs_2_addr_n4187;
output      [3:0] PE0_act_regs_1_addr_n4191;
output      [3:0] PE0_act_regs_0_addr_n4195;
output      [3:0] PE0_act_regs_3_addr_n4207;
output      [3:0] PE0_act_regs_2_addr_n4211;
output      [3:0] PE0_act_regs_1_addr_n4215;
output      [3:0] PE0_act_regs_0_addr_n4219;
output     [31:0] pe0_act_buffer_addr_n4231;
output      [3:0] PE0_act_regs_3_addr_n4239;
output      [3:0] PE0_act_regs_2_addr_n4243;
output      [3:0] PE0_act_regs_1_addr_n4247;
output      [3:0] PE0_act_regs_0_addr_n4251;
output      [3:0] PE0_act_regs_3_addr_n4260;
output      [3:0] PE0_act_regs_2_addr_n4264;
output      [3:0] PE0_act_regs_1_addr_n4268;
output      [3:0] PE0_act_regs_0_addr_n4272;
output      [3:0] PE0_act_regs_3_addr_n4280;
output      [3:0] PE0_act_regs_2_addr_n4284;
output      [3:0] PE0_act_regs_1_addr_n4288;
output      [3:0] PE0_act_regs_0_addr_n4292;
output      [3:0] PE0_act_regs_3_addr_n4304;
output      [3:0] PE0_act_regs_2_addr_n4308;
output      [3:0] PE0_act_regs_1_addr_n4312;
output      [3:0] PE0_act_regs_0_addr_n4316;
output      [3:0] PE0_act_regs_3_addr_n4324;
output      [3:0] PE0_act_regs_2_addr_n4328;
output      [3:0] PE0_act_regs_1_addr_n4332;
output      [3:0] PE0_act_regs_0_addr_n4336;
output      [3:0] PE0_act_regs_3_addr_n4348;
output      [3:0] PE0_act_regs_2_addr_n4352;
output      [3:0] PE0_act_regs_1_addr_n4356;
output      [3:0] PE0_act_regs_0_addr_n4360;
output      [3:0] PE0_act_regs_3_addr_n4372;
output      [3:0] PE0_act_regs_2_addr_n4376;
output      [3:0] PE0_act_regs_1_addr_n4380;
output      [3:0] PE0_act_regs_0_addr_n4384;
output      [3:0] PE0_act_regs_3_addr_n4396;
output      [3:0] PE0_act_regs_2_addr_n4400;
output      [3:0] PE0_act_regs_1_addr_n4404;
output      [3:0] PE0_act_regs_0_addr_n4408;
output      [3:0] PE0_act_regs_3_addr_n4420;
output      [3:0] PE0_act_regs_2_addr_n4424;
output      [3:0] PE0_act_regs_1_addr_n4428;
output      [3:0] PE0_act_regs_0_addr_n4432;
output reg            rva_in_ready;
output reg            act_start_ready;
output reg            act_port_ready;
output reg    [127:0] output_port_data;
output reg      [7:0] output_port_addr;
output reg            output_port_valid;
output reg            done;
output reg            done_valid;
output reg            pe0_act_mngr_is_valid;
output reg            pe0_act_mngr_is_zero_first;
output reg      [2:0] pe0_act_mngr_adpfloat_bias;
output reg      [5:0] pe0_act_mngr_num_inst;
output reg      [7:0] pe0_act_mngr_num_output;
output reg      [4:0] pe0_act_mngr_buffer_addr_base;
output reg      [7:0] pe0_act_mngr_output_addr_base;
output reg      [7:0] act_vector_0_15_Inst_0;
output reg      [7:0] act_vector_0_15_Inst_1;
output reg      [7:0] act_vector_0_15_Inst_2;
output reg      [7:0] act_vector_0_15_Inst_3;
output reg      [7:0] act_vector_0_15_Inst_4;
output reg      [7:0] act_vector_0_15_Inst_5;
output reg      [7:0] act_vector_0_15_Inst_6;
output reg      [7:0] act_vector_0_15_Inst_7;
output reg      [7:0] act_vector_0_15_Inst_8;
output reg      [7:0] act_vector_0_15_Inst_9;
output reg      [7:0] act_vector_0_15_Inst_10;
output reg      [7:0] act_vector_0_15_Inst_11;
output reg      [7:0] act_vector_0_15_Inst_12;
output reg      [7:0] act_vector_0_15_Inst_13;
output reg      [7:0] act_vector_0_15_Inst_14;
output reg      [7:0] act_vector_0_15_Inst_15;
output reg      [7:0] act_vector_16_31_Inst_0;
output reg      [7:0] act_vector_16_31_Inst_1;
output reg      [7:0] act_vector_16_31_Inst_2;
output reg      [7:0] act_vector_16_31_Inst_3;
output reg      [7:0] act_vector_16_31_Inst_4;
output reg      [7:0] act_vector_16_31_Inst_5;
output reg      [7:0] act_vector_16_31_Inst_6;
output reg      [7:0] act_vector_16_31_Inst_7;
output reg      [7:0] act_vector_16_31_Inst_8;
output reg      [7:0] act_vector_16_31_Inst_9;
output reg      [7:0] act_vector_16_31_Inst_10;
output reg      [7:0] act_vector_16_31_Inst_11;
output reg      [7:0] act_vector_16_31_Inst_12;
output reg      [7:0] act_vector_16_31_Inst_13;
output reg      [7:0] act_vector_16_31_Inst_14;
output reg      [7:0] act_vector_16_31_Inst_15;
output reg            pe0_act_is_start_reg;
output reg      [5:0] pe0_act_instruction_counter;
output reg      [7:0] pe0_act_output_counter;
output reg      [1:0] pe0_act_state;
output reg     [19:0] PE0_act_reg_temp_0;
output reg     [19:0] PE0_act_reg_temp_1;
output reg     [19:0] PE0_act_reg_temp_2;
output reg     [19:0] PE0_act_reg_temp_3;
output reg     [19:0] PE0_act_reg_temp_4;
output reg     [19:0] PE0_act_reg_temp_5;
output reg     [19:0] PE0_act_reg_temp_6;
output reg     [19:0] PE0_act_reg_temp_7;
output reg     [19:0] PE0_act_reg_temp_8;
output reg     [19:0] PE0_act_reg_temp_9;
output reg     [19:0] PE0_act_reg_temp_10;
output reg     [19:0] PE0_act_reg_temp_11;
output reg     [19:0] PE0_act_reg_temp_12;
output reg     [19:0] PE0_act_reg_temp_13;
output reg     [19:0] PE0_act_reg_temp_14;
output reg     [19:0] PE0_act_reg_temp_15;
wire      [3:0] PE0_act_regs_0_addr0;
wire      [3:0] PE0_act_regs_0_addr1;
wire      [3:0] PE0_act_regs_0_addr10;
wire      [3:0] PE0_act_regs_0_addr11;
wire      [3:0] PE0_act_regs_0_addr12;
wire      [3:0] PE0_act_regs_0_addr13;
wire      [3:0] PE0_act_regs_0_addr14;
wire      [3:0] PE0_act_regs_0_addr15;
wire      [3:0] PE0_act_regs_0_addr2;
wire      [3:0] PE0_act_regs_0_addr3;
wire      [3:0] PE0_act_regs_0_addr4;
wire      [3:0] PE0_act_regs_0_addr5;
wire      [3:0] PE0_act_regs_0_addr6;
wire      [3:0] PE0_act_regs_0_addr7;
wire      [3:0] PE0_act_regs_0_addr8;
wire      [3:0] PE0_act_regs_0_addr9;
wire      [3:0] PE0_act_regs_0_addr_n1056;
wire      [3:0] PE0_act_regs_0_addr_n1077;
wire      [3:0] PE0_act_regs_0_addr_n1097;
wire      [3:0] PE0_act_regs_0_addr_n1121;
wire      [3:0] PE0_act_regs_0_addr_n1141;
wire      [3:0] PE0_act_regs_0_addr_n1165;
wire      [3:0] PE0_act_regs_0_addr_n1189;
wire      [3:0] PE0_act_regs_0_addr_n1213;
wire      [3:0] PE0_act_regs_0_addr_n1237;
wire      [3:0] PE0_act_regs_0_addr_n1269;
wire      [3:0] PE0_act_regs_0_addr_n1290;
wire      [3:0] PE0_act_regs_0_addr_n1310;
wire      [3:0] PE0_act_regs_0_addr_n1334;
wire      [3:0] PE0_act_regs_0_addr_n1354;
wire      [3:0] PE0_act_regs_0_addr_n1378;
wire      [3:0] PE0_act_regs_0_addr_n1402;
wire      [3:0] PE0_act_regs_0_addr_n1426;
wire      [3:0] PE0_act_regs_0_addr_n1450;
wire      [3:0] PE0_act_regs_0_addr_n1482;
wire      [3:0] PE0_act_regs_0_addr_n1503;
wire      [3:0] PE0_act_regs_0_addr_n1523;
wire      [3:0] PE0_act_regs_0_addr_n1547;
wire      [3:0] PE0_act_regs_0_addr_n1567;
wire      [3:0] PE0_act_regs_0_addr_n1591;
wire      [3:0] PE0_act_regs_0_addr_n1615;
wire      [3:0] PE0_act_regs_0_addr_n1639;
wire      [3:0] PE0_act_regs_0_addr_n1663;
wire      [3:0] PE0_act_regs_0_addr_n1695;
wire      [3:0] PE0_act_regs_0_addr_n1716;
wire      [3:0] PE0_act_regs_0_addr_n1736;
wire      [3:0] PE0_act_regs_0_addr_n1760;
wire      [3:0] PE0_act_regs_0_addr_n1780;
wire      [3:0] PE0_act_regs_0_addr_n1804;
wire      [3:0] PE0_act_regs_0_addr_n1828;
wire      [3:0] PE0_act_regs_0_addr_n1852;
wire      [3:0] PE0_act_regs_0_addr_n1876;
wire      [3:0] PE0_act_regs_0_addr_n1908;
wire      [3:0] PE0_act_regs_0_addr_n1929;
wire      [3:0] PE0_act_regs_0_addr_n1949;
wire      [3:0] PE0_act_regs_0_addr_n1973;
wire      [3:0] PE0_act_regs_0_addr_n1993;
wire      [3:0] PE0_act_regs_0_addr_n2017;
wire      [3:0] PE0_act_regs_0_addr_n2041;
wire      [3:0] PE0_act_regs_0_addr_n2065;
wire      [3:0] PE0_act_regs_0_addr_n2089;
wire      [3:0] PE0_act_regs_0_addr_n2121;
wire      [3:0] PE0_act_regs_0_addr_n2142;
wire      [3:0] PE0_act_regs_0_addr_n2162;
wire      [3:0] PE0_act_regs_0_addr_n2186;
wire      [3:0] PE0_act_regs_0_addr_n2206;
wire      [3:0] PE0_act_regs_0_addr_n2230;
wire      [3:0] PE0_act_regs_0_addr_n2254;
wire      [3:0] PE0_act_regs_0_addr_n2278;
wire      [3:0] PE0_act_regs_0_addr_n2302;
wire      [3:0] PE0_act_regs_0_addr_n2334;
wire      [3:0] PE0_act_regs_0_addr_n2355;
wire      [3:0] PE0_act_regs_0_addr_n2375;
wire      [3:0] PE0_act_regs_0_addr_n2399;
wire      [3:0] PE0_act_regs_0_addr_n2419;
wire      [3:0] PE0_act_regs_0_addr_n2443;
wire      [3:0] PE0_act_regs_0_addr_n2467;
wire      [3:0] PE0_act_regs_0_addr_n2491;
wire      [3:0] PE0_act_regs_0_addr_n2515;
wire      [3:0] PE0_act_regs_0_addr_n2547;
wire      [3:0] PE0_act_regs_0_addr_n2568;
wire      [3:0] PE0_act_regs_0_addr_n2588;
wire      [3:0] PE0_act_regs_0_addr_n2612;
wire      [3:0] PE0_act_regs_0_addr_n2632;
wire      [3:0] PE0_act_regs_0_addr_n2656;
wire      [3:0] PE0_act_regs_0_addr_n2680;
wire      [3:0] PE0_act_regs_0_addr_n2704;
wire      [3:0] PE0_act_regs_0_addr_n2728;
wire      [3:0] PE0_act_regs_0_addr_n2760;
wire      [3:0] PE0_act_regs_0_addr_n2781;
wire      [3:0] PE0_act_regs_0_addr_n2801;
wire      [3:0] PE0_act_regs_0_addr_n2825;
wire      [3:0] PE0_act_regs_0_addr_n2845;
wire      [3:0] PE0_act_regs_0_addr_n2869;
wire      [3:0] PE0_act_regs_0_addr_n2893;
wire      [3:0] PE0_act_regs_0_addr_n2917;
wire      [3:0] PE0_act_regs_0_addr_n2941;
wire      [3:0] PE0_act_regs_0_addr_n2973;
wire      [3:0] PE0_act_regs_0_addr_n2994;
wire      [3:0] PE0_act_regs_0_addr_n3014;
wire      [3:0] PE0_act_regs_0_addr_n3038;
wire      [3:0] PE0_act_regs_0_addr_n3058;
wire      [3:0] PE0_act_regs_0_addr_n3082;
wire      [3:0] PE0_act_regs_0_addr_n3106;
wire      [3:0] PE0_act_regs_0_addr_n3130;
wire      [3:0] PE0_act_regs_0_addr_n3154;
wire      [3:0] PE0_act_regs_0_addr_n3186;
wire      [3:0] PE0_act_regs_0_addr_n3207;
wire      [3:0] PE0_act_regs_0_addr_n3227;
wire      [3:0] PE0_act_regs_0_addr_n3251;
wire      [3:0] PE0_act_regs_0_addr_n3271;
wire      [3:0] PE0_act_regs_0_addr_n3295;
wire      [3:0] PE0_act_regs_0_addr_n3319;
wire      [3:0] PE0_act_regs_0_addr_n3343;
wire      [3:0] PE0_act_regs_0_addr_n3367;
wire      [3:0] PE0_act_regs_0_addr_n3399;
wire      [3:0] PE0_act_regs_0_addr_n3420;
wire      [3:0] PE0_act_regs_0_addr_n3440;
wire      [3:0] PE0_act_regs_0_addr_n3464;
wire      [3:0] PE0_act_regs_0_addr_n3484;
wire      [3:0] PE0_act_regs_0_addr_n3508;
wire      [3:0] PE0_act_regs_0_addr_n3532;
wire      [3:0] PE0_act_regs_0_addr_n3556;
wire      [3:0] PE0_act_regs_0_addr_n3580;
wire      [3:0] PE0_act_regs_0_addr_n3612;
wire      [3:0] PE0_act_regs_0_addr_n3633;
wire      [3:0] PE0_act_regs_0_addr_n3653;
wire      [3:0] PE0_act_regs_0_addr_n3677;
wire      [3:0] PE0_act_regs_0_addr_n3697;
wire      [3:0] PE0_act_regs_0_addr_n3721;
wire      [3:0] PE0_act_regs_0_addr_n3745;
wire      [3:0] PE0_act_regs_0_addr_n3769;
wire      [3:0] PE0_act_regs_0_addr_n3793;
wire      [3:0] PE0_act_regs_0_addr_n3825;
wire      [3:0] PE0_act_regs_0_addr_n3846;
wire      [3:0] PE0_act_regs_0_addr_n3866;
wire      [3:0] PE0_act_regs_0_addr_n3890;
wire      [3:0] PE0_act_regs_0_addr_n3910;
wire      [3:0] PE0_act_regs_0_addr_n3934;
wire      [3:0] PE0_act_regs_0_addr_n3958;
wire      [3:0] PE0_act_regs_0_addr_n3982;
wire      [3:0] PE0_act_regs_0_addr_n4006;
wire      [3:0] PE0_act_regs_0_addr_n4038;
wire      [3:0] PE0_act_regs_0_addr_n4059;
wire      [3:0] PE0_act_regs_0_addr_n4079;
wire      [3:0] PE0_act_regs_0_addr_n4103;
wire      [3:0] PE0_act_regs_0_addr_n4123;
wire      [3:0] PE0_act_regs_0_addr_n4147;
wire      [3:0] PE0_act_regs_0_addr_n416;
wire      [3:0] PE0_act_regs_0_addr_n4171;
wire      [3:0] PE0_act_regs_0_addr_n4195;
wire      [3:0] PE0_act_regs_0_addr_n4219;
wire      [3:0] PE0_act_regs_0_addr_n4251;
wire      [3:0] PE0_act_regs_0_addr_n4272;
wire      [3:0] PE0_act_regs_0_addr_n4292;
wire      [3:0] PE0_act_regs_0_addr_n4316;
wire      [3:0] PE0_act_regs_0_addr_n4336;
wire      [3:0] PE0_act_regs_0_addr_n4360;
wire      [3:0] PE0_act_regs_0_addr_n4384;
wire      [3:0] PE0_act_regs_0_addr_n4408;
wire      [3:0] PE0_act_regs_0_addr_n443;
wire      [3:0] PE0_act_regs_0_addr_n4432;
wire      [3:0] PE0_act_regs_0_addr_n468;
wire      [3:0] PE0_act_regs_0_addr_n493;
wire      [3:0] PE0_act_regs_0_addr_n518;
wire      [3:0] PE0_act_regs_0_addr_n543;
wire      [3:0] PE0_act_regs_0_addr_n568;
wire      [3:0] PE0_act_regs_0_addr_n593;
wire      [3:0] PE0_act_regs_0_addr_n618;
wire      [3:0] PE0_act_regs_0_addr_n644;
wire      [3:0] PE0_act_regs_0_addr_n670;
wire      [3:0] PE0_act_regs_0_addr_n695;
wire      [3:0] PE0_act_regs_0_addr_n720;
wire      [3:0] PE0_act_regs_0_addr_n745;
wire      [3:0] PE0_act_regs_0_addr_n770;
wire      [3:0] PE0_act_regs_0_addr_n795;
wire     [19:0] PE0_act_regs_0_data0;
wire     [19:0] PE0_act_regs_0_data1;
wire     [19:0] PE0_act_regs_0_data10;
wire     [19:0] PE0_act_regs_0_data11;
wire     [19:0] PE0_act_regs_0_data12;
wire     [19:0] PE0_act_regs_0_data13;
wire     [19:0] PE0_act_regs_0_data14;
wire     [19:0] PE0_act_regs_0_data15;
wire     [19:0] PE0_act_regs_0_data2;
wire     [19:0] PE0_act_regs_0_data3;
wire     [19:0] PE0_act_regs_0_data4;
wire     [19:0] PE0_act_regs_0_data5;
wire     [19:0] PE0_act_regs_0_data6;
wire     [19:0] PE0_act_regs_0_data7;
wire     [19:0] PE0_act_regs_0_data8;
wire     [19:0] PE0_act_regs_0_data9;
wire     [19:0] PE0_act_regs_0_data_n1057;
wire     [19:0] PE0_act_regs_0_data_n1078;
wire     [19:0] PE0_act_regs_0_data_n1098;
wire     [19:0] PE0_act_regs_0_data_n1122;
wire     [19:0] PE0_act_regs_0_data_n1142;
wire     [19:0] PE0_act_regs_0_data_n1166;
wire     [19:0] PE0_act_regs_0_data_n1190;
wire     [19:0] PE0_act_regs_0_data_n1214;
wire     [19:0] PE0_act_regs_0_data_n1238;
wire     [19:0] PE0_act_regs_0_data_n1270;
wire     [19:0] PE0_act_regs_0_data_n1291;
wire     [19:0] PE0_act_regs_0_data_n1311;
wire     [19:0] PE0_act_regs_0_data_n1335;
wire     [19:0] PE0_act_regs_0_data_n1355;
wire     [19:0] PE0_act_regs_0_data_n1379;
wire     [19:0] PE0_act_regs_0_data_n1403;
wire     [19:0] PE0_act_regs_0_data_n1427;
wire     [19:0] PE0_act_regs_0_data_n1451;
wire     [19:0] PE0_act_regs_0_data_n1483;
wire     [19:0] PE0_act_regs_0_data_n1504;
wire     [19:0] PE0_act_regs_0_data_n1524;
wire     [19:0] PE0_act_regs_0_data_n1548;
wire     [19:0] PE0_act_regs_0_data_n1568;
wire     [19:0] PE0_act_regs_0_data_n1592;
wire     [19:0] PE0_act_regs_0_data_n1616;
wire     [19:0] PE0_act_regs_0_data_n1640;
wire     [19:0] PE0_act_regs_0_data_n1664;
wire     [19:0] PE0_act_regs_0_data_n1696;
wire     [19:0] PE0_act_regs_0_data_n1717;
wire     [19:0] PE0_act_regs_0_data_n1737;
wire     [19:0] PE0_act_regs_0_data_n1761;
wire     [19:0] PE0_act_regs_0_data_n1781;
wire     [19:0] PE0_act_regs_0_data_n1805;
wire     [19:0] PE0_act_regs_0_data_n1829;
wire     [19:0] PE0_act_regs_0_data_n1853;
wire     [19:0] PE0_act_regs_0_data_n1877;
wire     [19:0] PE0_act_regs_0_data_n1909;
wire     [19:0] PE0_act_regs_0_data_n1930;
wire     [19:0] PE0_act_regs_0_data_n1950;
wire     [19:0] PE0_act_regs_0_data_n1974;
wire     [19:0] PE0_act_regs_0_data_n1994;
wire     [19:0] PE0_act_regs_0_data_n2018;
wire     [19:0] PE0_act_regs_0_data_n2042;
wire     [19:0] PE0_act_regs_0_data_n2066;
wire     [19:0] PE0_act_regs_0_data_n2090;
wire     [19:0] PE0_act_regs_0_data_n2122;
wire     [19:0] PE0_act_regs_0_data_n2143;
wire     [19:0] PE0_act_regs_0_data_n2163;
wire     [19:0] PE0_act_regs_0_data_n2187;
wire     [19:0] PE0_act_regs_0_data_n2207;
wire     [19:0] PE0_act_regs_0_data_n2231;
wire     [19:0] PE0_act_regs_0_data_n2255;
wire     [19:0] PE0_act_regs_0_data_n2279;
wire     [19:0] PE0_act_regs_0_data_n2303;
wire     [19:0] PE0_act_regs_0_data_n2335;
wire     [19:0] PE0_act_regs_0_data_n2356;
wire     [19:0] PE0_act_regs_0_data_n2376;
wire     [19:0] PE0_act_regs_0_data_n2400;
wire     [19:0] PE0_act_regs_0_data_n2420;
wire     [19:0] PE0_act_regs_0_data_n2444;
wire     [19:0] PE0_act_regs_0_data_n2468;
wire     [19:0] PE0_act_regs_0_data_n2492;
wire     [19:0] PE0_act_regs_0_data_n2516;
wire     [19:0] PE0_act_regs_0_data_n2548;
wire     [19:0] PE0_act_regs_0_data_n2569;
wire     [19:0] PE0_act_regs_0_data_n2589;
wire     [19:0] PE0_act_regs_0_data_n2613;
wire     [19:0] PE0_act_regs_0_data_n2633;
wire     [19:0] PE0_act_regs_0_data_n2657;
wire     [19:0] PE0_act_regs_0_data_n2681;
wire     [19:0] PE0_act_regs_0_data_n2705;
wire     [19:0] PE0_act_regs_0_data_n2729;
wire     [19:0] PE0_act_regs_0_data_n2761;
wire     [19:0] PE0_act_regs_0_data_n2782;
wire     [19:0] PE0_act_regs_0_data_n2802;
wire     [19:0] PE0_act_regs_0_data_n2826;
wire     [19:0] PE0_act_regs_0_data_n2846;
wire     [19:0] PE0_act_regs_0_data_n2870;
wire     [19:0] PE0_act_regs_0_data_n2894;
wire     [19:0] PE0_act_regs_0_data_n2918;
wire     [19:0] PE0_act_regs_0_data_n2942;
wire     [19:0] PE0_act_regs_0_data_n2974;
wire     [19:0] PE0_act_regs_0_data_n2995;
wire     [19:0] PE0_act_regs_0_data_n3015;
wire     [19:0] PE0_act_regs_0_data_n3039;
wire     [19:0] PE0_act_regs_0_data_n3059;
wire     [19:0] PE0_act_regs_0_data_n3083;
wire     [19:0] PE0_act_regs_0_data_n3107;
wire     [19:0] PE0_act_regs_0_data_n3131;
wire     [19:0] PE0_act_regs_0_data_n3155;
wire     [19:0] PE0_act_regs_0_data_n3187;
wire     [19:0] PE0_act_regs_0_data_n3208;
wire     [19:0] PE0_act_regs_0_data_n3228;
wire     [19:0] PE0_act_regs_0_data_n3252;
wire     [19:0] PE0_act_regs_0_data_n3272;
wire     [19:0] PE0_act_regs_0_data_n3296;
wire     [19:0] PE0_act_regs_0_data_n3320;
wire     [19:0] PE0_act_regs_0_data_n3344;
wire     [19:0] PE0_act_regs_0_data_n3368;
wire     [19:0] PE0_act_regs_0_data_n3400;
wire     [19:0] PE0_act_regs_0_data_n3421;
wire     [19:0] PE0_act_regs_0_data_n3441;
wire     [19:0] PE0_act_regs_0_data_n3465;
wire     [19:0] PE0_act_regs_0_data_n3485;
wire     [19:0] PE0_act_regs_0_data_n3509;
wire     [19:0] PE0_act_regs_0_data_n3533;
wire     [19:0] PE0_act_regs_0_data_n3557;
wire     [19:0] PE0_act_regs_0_data_n3581;
wire     [19:0] PE0_act_regs_0_data_n3613;
wire     [19:0] PE0_act_regs_0_data_n3634;
wire     [19:0] PE0_act_regs_0_data_n3654;
wire     [19:0] PE0_act_regs_0_data_n3678;
wire     [19:0] PE0_act_regs_0_data_n3698;
wire     [19:0] PE0_act_regs_0_data_n3722;
wire     [19:0] PE0_act_regs_0_data_n3746;
wire     [19:0] PE0_act_regs_0_data_n3770;
wire     [19:0] PE0_act_regs_0_data_n3794;
wire     [19:0] PE0_act_regs_0_data_n3826;
wire     [19:0] PE0_act_regs_0_data_n3847;
wire     [19:0] PE0_act_regs_0_data_n3867;
wire     [19:0] PE0_act_regs_0_data_n3891;
wire     [19:0] PE0_act_regs_0_data_n3911;
wire     [19:0] PE0_act_regs_0_data_n3935;
wire     [19:0] PE0_act_regs_0_data_n3959;
wire     [19:0] PE0_act_regs_0_data_n3983;
wire     [19:0] PE0_act_regs_0_data_n4007;
wire     [19:0] PE0_act_regs_0_data_n4039;
wire     [19:0] PE0_act_regs_0_data_n4060;
wire     [19:0] PE0_act_regs_0_data_n4080;
wire     [19:0] PE0_act_regs_0_data_n4104;
wire     [19:0] PE0_act_regs_0_data_n4124;
wire     [19:0] PE0_act_regs_0_data_n4148;
wire     [19:0] PE0_act_regs_0_data_n417;
wire     [19:0] PE0_act_regs_0_data_n4172;
wire     [19:0] PE0_act_regs_0_data_n4196;
wire     [19:0] PE0_act_regs_0_data_n4220;
wire     [19:0] PE0_act_regs_0_data_n4252;
wire     [19:0] PE0_act_regs_0_data_n4273;
wire     [19:0] PE0_act_regs_0_data_n4293;
wire     [19:0] PE0_act_regs_0_data_n4317;
wire     [19:0] PE0_act_regs_0_data_n4337;
wire     [19:0] PE0_act_regs_0_data_n4361;
wire     [19:0] PE0_act_regs_0_data_n4385;
wire     [19:0] PE0_act_regs_0_data_n4409;
wire     [19:0] PE0_act_regs_0_data_n4433;
wire     [19:0] PE0_act_regs_0_data_n444;
wire     [19:0] PE0_act_regs_0_data_n469;
wire     [19:0] PE0_act_regs_0_data_n494;
wire     [19:0] PE0_act_regs_0_data_n519;
wire     [19:0] PE0_act_regs_0_data_n544;
wire     [19:0] PE0_act_regs_0_data_n569;
wire     [19:0] PE0_act_regs_0_data_n594;
wire     [19:0] PE0_act_regs_0_data_n619;
wire     [19:0] PE0_act_regs_0_data_n645;
wire     [19:0] PE0_act_regs_0_data_n671;
wire     [19:0] PE0_act_regs_0_data_n696;
wire     [19:0] PE0_act_regs_0_data_n721;
wire     [19:0] PE0_act_regs_0_data_n746;
wire     [19:0] PE0_act_regs_0_data_n771;
wire     [19:0] PE0_act_regs_0_data_n796;
wire            PE0_act_regs_0_wen0;
wire            PE0_act_regs_0_wen1;
wire            PE0_act_regs_0_wen10;
wire            PE0_act_regs_0_wen11;
wire            PE0_act_regs_0_wen12;
wire            PE0_act_regs_0_wen13;
wire            PE0_act_regs_0_wen14;
wire            PE0_act_regs_0_wen15;
wire            PE0_act_regs_0_wen2;
wire            PE0_act_regs_0_wen3;
wire            PE0_act_regs_0_wen4;
wire            PE0_act_regs_0_wen5;
wire            PE0_act_regs_0_wen6;
wire            PE0_act_regs_0_wen7;
wire            PE0_act_regs_0_wen8;
wire            PE0_act_regs_0_wen9;
wire      [3:0] PE0_act_regs_1_addr0;
wire      [3:0] PE0_act_regs_1_addr1;
wire      [3:0] PE0_act_regs_1_addr10;
wire      [3:0] PE0_act_regs_1_addr11;
wire      [3:0] PE0_act_regs_1_addr12;
wire      [3:0] PE0_act_regs_1_addr13;
wire      [3:0] PE0_act_regs_1_addr14;
wire      [3:0] PE0_act_regs_1_addr15;
wire      [3:0] PE0_act_regs_1_addr2;
wire      [3:0] PE0_act_regs_1_addr3;
wire      [3:0] PE0_act_regs_1_addr4;
wire      [3:0] PE0_act_regs_1_addr5;
wire      [3:0] PE0_act_regs_1_addr6;
wire      [3:0] PE0_act_regs_1_addr7;
wire      [3:0] PE0_act_regs_1_addr8;
wire      [3:0] PE0_act_regs_1_addr9;
wire      [3:0] PE0_act_regs_1_addr_n1052;
wire      [3:0] PE0_act_regs_1_addr_n1073;
wire      [3:0] PE0_act_regs_1_addr_n1093;
wire      [3:0] PE0_act_regs_1_addr_n1117;
wire      [3:0] PE0_act_regs_1_addr_n1137;
wire      [3:0] PE0_act_regs_1_addr_n1161;
wire      [3:0] PE0_act_regs_1_addr_n1185;
wire      [3:0] PE0_act_regs_1_addr_n1209;
wire      [3:0] PE0_act_regs_1_addr_n1233;
wire      [3:0] PE0_act_regs_1_addr_n1265;
wire      [3:0] PE0_act_regs_1_addr_n1286;
wire      [3:0] PE0_act_regs_1_addr_n1306;
wire      [3:0] PE0_act_regs_1_addr_n1330;
wire      [3:0] PE0_act_regs_1_addr_n1350;
wire      [3:0] PE0_act_regs_1_addr_n1374;
wire      [3:0] PE0_act_regs_1_addr_n1398;
wire      [3:0] PE0_act_regs_1_addr_n1422;
wire      [3:0] PE0_act_regs_1_addr_n1446;
wire      [3:0] PE0_act_regs_1_addr_n1478;
wire      [3:0] PE0_act_regs_1_addr_n1499;
wire      [3:0] PE0_act_regs_1_addr_n1519;
wire      [3:0] PE0_act_regs_1_addr_n1543;
wire      [3:0] PE0_act_regs_1_addr_n1563;
wire      [3:0] PE0_act_regs_1_addr_n1587;
wire      [3:0] PE0_act_regs_1_addr_n1611;
wire      [3:0] PE0_act_regs_1_addr_n1635;
wire      [3:0] PE0_act_regs_1_addr_n1659;
wire      [3:0] PE0_act_regs_1_addr_n1691;
wire      [3:0] PE0_act_regs_1_addr_n1712;
wire      [3:0] PE0_act_regs_1_addr_n1732;
wire      [3:0] PE0_act_regs_1_addr_n1756;
wire      [3:0] PE0_act_regs_1_addr_n1776;
wire      [3:0] PE0_act_regs_1_addr_n1800;
wire      [3:0] PE0_act_regs_1_addr_n1824;
wire      [3:0] PE0_act_regs_1_addr_n1848;
wire      [3:0] PE0_act_regs_1_addr_n1872;
wire      [3:0] PE0_act_regs_1_addr_n1904;
wire      [3:0] PE0_act_regs_1_addr_n1925;
wire      [3:0] PE0_act_regs_1_addr_n1945;
wire      [3:0] PE0_act_regs_1_addr_n1969;
wire      [3:0] PE0_act_regs_1_addr_n1989;
wire      [3:0] PE0_act_regs_1_addr_n2013;
wire      [3:0] PE0_act_regs_1_addr_n2037;
wire      [3:0] PE0_act_regs_1_addr_n2061;
wire      [3:0] PE0_act_regs_1_addr_n2085;
wire      [3:0] PE0_act_regs_1_addr_n2117;
wire      [3:0] PE0_act_regs_1_addr_n2138;
wire      [3:0] PE0_act_regs_1_addr_n2158;
wire      [3:0] PE0_act_regs_1_addr_n2182;
wire      [3:0] PE0_act_regs_1_addr_n2202;
wire      [3:0] PE0_act_regs_1_addr_n2226;
wire      [3:0] PE0_act_regs_1_addr_n2250;
wire      [3:0] PE0_act_regs_1_addr_n2274;
wire      [3:0] PE0_act_regs_1_addr_n2298;
wire      [3:0] PE0_act_regs_1_addr_n2330;
wire      [3:0] PE0_act_regs_1_addr_n2351;
wire      [3:0] PE0_act_regs_1_addr_n2371;
wire      [3:0] PE0_act_regs_1_addr_n2395;
wire      [3:0] PE0_act_regs_1_addr_n2415;
wire      [3:0] PE0_act_regs_1_addr_n2439;
wire      [3:0] PE0_act_regs_1_addr_n2463;
wire      [3:0] PE0_act_regs_1_addr_n2487;
wire      [3:0] PE0_act_regs_1_addr_n2511;
wire      [3:0] PE0_act_regs_1_addr_n2543;
wire      [3:0] PE0_act_regs_1_addr_n2564;
wire      [3:0] PE0_act_regs_1_addr_n2584;
wire      [3:0] PE0_act_regs_1_addr_n2608;
wire      [3:0] PE0_act_regs_1_addr_n2628;
wire      [3:0] PE0_act_regs_1_addr_n2652;
wire      [3:0] PE0_act_regs_1_addr_n2676;
wire      [3:0] PE0_act_regs_1_addr_n2700;
wire      [3:0] PE0_act_regs_1_addr_n2724;
wire      [3:0] PE0_act_regs_1_addr_n2756;
wire      [3:0] PE0_act_regs_1_addr_n2777;
wire      [3:0] PE0_act_regs_1_addr_n2797;
wire      [3:0] PE0_act_regs_1_addr_n2821;
wire      [3:0] PE0_act_regs_1_addr_n2841;
wire      [3:0] PE0_act_regs_1_addr_n2865;
wire      [3:0] PE0_act_regs_1_addr_n2889;
wire      [3:0] PE0_act_regs_1_addr_n2913;
wire      [3:0] PE0_act_regs_1_addr_n2937;
wire      [3:0] PE0_act_regs_1_addr_n2969;
wire      [3:0] PE0_act_regs_1_addr_n2990;
wire      [3:0] PE0_act_regs_1_addr_n3010;
wire      [3:0] PE0_act_regs_1_addr_n3034;
wire      [3:0] PE0_act_regs_1_addr_n3054;
wire      [3:0] PE0_act_regs_1_addr_n3078;
wire      [3:0] PE0_act_regs_1_addr_n3102;
wire      [3:0] PE0_act_regs_1_addr_n3126;
wire      [3:0] PE0_act_regs_1_addr_n3150;
wire      [3:0] PE0_act_regs_1_addr_n3182;
wire      [3:0] PE0_act_regs_1_addr_n3203;
wire      [3:0] PE0_act_regs_1_addr_n3223;
wire      [3:0] PE0_act_regs_1_addr_n3247;
wire      [3:0] PE0_act_regs_1_addr_n3267;
wire      [3:0] PE0_act_regs_1_addr_n3291;
wire      [3:0] PE0_act_regs_1_addr_n3315;
wire      [3:0] PE0_act_regs_1_addr_n3339;
wire      [3:0] PE0_act_regs_1_addr_n3363;
wire      [3:0] PE0_act_regs_1_addr_n3395;
wire      [3:0] PE0_act_regs_1_addr_n3416;
wire      [3:0] PE0_act_regs_1_addr_n3436;
wire      [3:0] PE0_act_regs_1_addr_n3460;
wire      [3:0] PE0_act_regs_1_addr_n3480;
wire      [3:0] PE0_act_regs_1_addr_n3504;
wire      [3:0] PE0_act_regs_1_addr_n3528;
wire      [3:0] PE0_act_regs_1_addr_n3552;
wire      [3:0] PE0_act_regs_1_addr_n3576;
wire      [3:0] PE0_act_regs_1_addr_n3608;
wire      [3:0] PE0_act_regs_1_addr_n3629;
wire      [3:0] PE0_act_regs_1_addr_n3649;
wire      [3:0] PE0_act_regs_1_addr_n3673;
wire      [3:0] PE0_act_regs_1_addr_n3693;
wire      [3:0] PE0_act_regs_1_addr_n3717;
wire      [3:0] PE0_act_regs_1_addr_n3741;
wire      [3:0] PE0_act_regs_1_addr_n3765;
wire      [3:0] PE0_act_regs_1_addr_n3789;
wire      [3:0] PE0_act_regs_1_addr_n3821;
wire      [3:0] PE0_act_regs_1_addr_n3842;
wire      [3:0] PE0_act_regs_1_addr_n3862;
wire      [3:0] PE0_act_regs_1_addr_n3886;
wire      [3:0] PE0_act_regs_1_addr_n3906;
wire      [3:0] PE0_act_regs_1_addr_n3930;
wire      [3:0] PE0_act_regs_1_addr_n3954;
wire      [3:0] PE0_act_regs_1_addr_n3978;
wire      [3:0] PE0_act_regs_1_addr_n4002;
wire      [3:0] PE0_act_regs_1_addr_n4034;
wire      [3:0] PE0_act_regs_1_addr_n4055;
wire      [3:0] PE0_act_regs_1_addr_n4075;
wire      [3:0] PE0_act_regs_1_addr_n4099;
wire      [3:0] PE0_act_regs_1_addr_n4119;
wire      [3:0] PE0_act_regs_1_addr_n412;
wire      [3:0] PE0_act_regs_1_addr_n4143;
wire      [3:0] PE0_act_regs_1_addr_n4167;
wire      [3:0] PE0_act_regs_1_addr_n4191;
wire      [3:0] PE0_act_regs_1_addr_n4215;
wire      [3:0] PE0_act_regs_1_addr_n4247;
wire      [3:0] PE0_act_regs_1_addr_n4268;
wire      [3:0] PE0_act_regs_1_addr_n4288;
wire      [3:0] PE0_act_regs_1_addr_n4312;
wire      [3:0] PE0_act_regs_1_addr_n4332;
wire      [3:0] PE0_act_regs_1_addr_n4356;
wire      [3:0] PE0_act_regs_1_addr_n4380;
wire      [3:0] PE0_act_regs_1_addr_n439;
wire      [3:0] PE0_act_regs_1_addr_n4404;
wire      [3:0] PE0_act_regs_1_addr_n4428;
wire      [3:0] PE0_act_regs_1_addr_n464;
wire      [3:0] PE0_act_regs_1_addr_n489;
wire      [3:0] PE0_act_regs_1_addr_n514;
wire      [3:0] PE0_act_regs_1_addr_n539;
wire      [3:0] PE0_act_regs_1_addr_n564;
wire      [3:0] PE0_act_regs_1_addr_n589;
wire      [3:0] PE0_act_regs_1_addr_n614;
wire      [3:0] PE0_act_regs_1_addr_n640;
wire      [3:0] PE0_act_regs_1_addr_n666;
wire      [3:0] PE0_act_regs_1_addr_n691;
wire      [3:0] PE0_act_regs_1_addr_n716;
wire      [3:0] PE0_act_regs_1_addr_n741;
wire      [3:0] PE0_act_regs_1_addr_n766;
wire      [3:0] PE0_act_regs_1_addr_n791;
wire     [19:0] PE0_act_regs_1_data0;
wire     [19:0] PE0_act_regs_1_data1;
wire     [19:0] PE0_act_regs_1_data10;
wire     [19:0] PE0_act_regs_1_data11;
wire     [19:0] PE0_act_regs_1_data12;
wire     [19:0] PE0_act_regs_1_data13;
wire     [19:0] PE0_act_regs_1_data14;
wire     [19:0] PE0_act_regs_1_data15;
wire     [19:0] PE0_act_regs_1_data2;
wire     [19:0] PE0_act_regs_1_data3;
wire     [19:0] PE0_act_regs_1_data4;
wire     [19:0] PE0_act_regs_1_data5;
wire     [19:0] PE0_act_regs_1_data6;
wire     [19:0] PE0_act_regs_1_data7;
wire     [19:0] PE0_act_regs_1_data8;
wire     [19:0] PE0_act_regs_1_data9;
wire     [19:0] PE0_act_regs_1_data_n1053;
wire     [19:0] PE0_act_regs_1_data_n1074;
wire     [19:0] PE0_act_regs_1_data_n1094;
wire     [19:0] PE0_act_regs_1_data_n1118;
wire     [19:0] PE0_act_regs_1_data_n1138;
wire     [19:0] PE0_act_regs_1_data_n1162;
wire     [19:0] PE0_act_regs_1_data_n1186;
wire     [19:0] PE0_act_regs_1_data_n1210;
wire     [19:0] PE0_act_regs_1_data_n1234;
wire     [19:0] PE0_act_regs_1_data_n1266;
wire     [19:0] PE0_act_regs_1_data_n1287;
wire     [19:0] PE0_act_regs_1_data_n1307;
wire     [19:0] PE0_act_regs_1_data_n1331;
wire     [19:0] PE0_act_regs_1_data_n1351;
wire     [19:0] PE0_act_regs_1_data_n1375;
wire     [19:0] PE0_act_regs_1_data_n1399;
wire     [19:0] PE0_act_regs_1_data_n1423;
wire     [19:0] PE0_act_regs_1_data_n1447;
wire     [19:0] PE0_act_regs_1_data_n1479;
wire     [19:0] PE0_act_regs_1_data_n1500;
wire     [19:0] PE0_act_regs_1_data_n1520;
wire     [19:0] PE0_act_regs_1_data_n1544;
wire     [19:0] PE0_act_regs_1_data_n1564;
wire     [19:0] PE0_act_regs_1_data_n1588;
wire     [19:0] PE0_act_regs_1_data_n1612;
wire     [19:0] PE0_act_regs_1_data_n1636;
wire     [19:0] PE0_act_regs_1_data_n1660;
wire     [19:0] PE0_act_regs_1_data_n1692;
wire     [19:0] PE0_act_regs_1_data_n1713;
wire     [19:0] PE0_act_regs_1_data_n1733;
wire     [19:0] PE0_act_regs_1_data_n1757;
wire     [19:0] PE0_act_regs_1_data_n1777;
wire     [19:0] PE0_act_regs_1_data_n1801;
wire     [19:0] PE0_act_regs_1_data_n1825;
wire     [19:0] PE0_act_regs_1_data_n1849;
wire     [19:0] PE0_act_regs_1_data_n1873;
wire     [19:0] PE0_act_regs_1_data_n1905;
wire     [19:0] PE0_act_regs_1_data_n1926;
wire     [19:0] PE0_act_regs_1_data_n1946;
wire     [19:0] PE0_act_regs_1_data_n1970;
wire     [19:0] PE0_act_regs_1_data_n1990;
wire     [19:0] PE0_act_regs_1_data_n2014;
wire     [19:0] PE0_act_regs_1_data_n2038;
wire     [19:0] PE0_act_regs_1_data_n2062;
wire     [19:0] PE0_act_regs_1_data_n2086;
wire     [19:0] PE0_act_regs_1_data_n2118;
wire     [19:0] PE0_act_regs_1_data_n2139;
wire     [19:0] PE0_act_regs_1_data_n2159;
wire     [19:0] PE0_act_regs_1_data_n2183;
wire     [19:0] PE0_act_regs_1_data_n2203;
wire     [19:0] PE0_act_regs_1_data_n2227;
wire     [19:0] PE0_act_regs_1_data_n2251;
wire     [19:0] PE0_act_regs_1_data_n2275;
wire     [19:0] PE0_act_regs_1_data_n2299;
wire     [19:0] PE0_act_regs_1_data_n2331;
wire     [19:0] PE0_act_regs_1_data_n2352;
wire     [19:0] PE0_act_regs_1_data_n2372;
wire     [19:0] PE0_act_regs_1_data_n2396;
wire     [19:0] PE0_act_regs_1_data_n2416;
wire     [19:0] PE0_act_regs_1_data_n2440;
wire     [19:0] PE0_act_regs_1_data_n2464;
wire     [19:0] PE0_act_regs_1_data_n2488;
wire     [19:0] PE0_act_regs_1_data_n2512;
wire     [19:0] PE0_act_regs_1_data_n2544;
wire     [19:0] PE0_act_regs_1_data_n2565;
wire     [19:0] PE0_act_regs_1_data_n2585;
wire     [19:0] PE0_act_regs_1_data_n2609;
wire     [19:0] PE0_act_regs_1_data_n2629;
wire     [19:0] PE0_act_regs_1_data_n2653;
wire     [19:0] PE0_act_regs_1_data_n2677;
wire     [19:0] PE0_act_regs_1_data_n2701;
wire     [19:0] PE0_act_regs_1_data_n2725;
wire     [19:0] PE0_act_regs_1_data_n2757;
wire     [19:0] PE0_act_regs_1_data_n2778;
wire     [19:0] PE0_act_regs_1_data_n2798;
wire     [19:0] PE0_act_regs_1_data_n2822;
wire     [19:0] PE0_act_regs_1_data_n2842;
wire     [19:0] PE0_act_regs_1_data_n2866;
wire     [19:0] PE0_act_regs_1_data_n2890;
wire     [19:0] PE0_act_regs_1_data_n2914;
wire     [19:0] PE0_act_regs_1_data_n2938;
wire     [19:0] PE0_act_regs_1_data_n2970;
wire     [19:0] PE0_act_regs_1_data_n2991;
wire     [19:0] PE0_act_regs_1_data_n3011;
wire     [19:0] PE0_act_regs_1_data_n3035;
wire     [19:0] PE0_act_regs_1_data_n3055;
wire     [19:0] PE0_act_regs_1_data_n3079;
wire     [19:0] PE0_act_regs_1_data_n3103;
wire     [19:0] PE0_act_regs_1_data_n3127;
wire     [19:0] PE0_act_regs_1_data_n3151;
wire     [19:0] PE0_act_regs_1_data_n3183;
wire     [19:0] PE0_act_regs_1_data_n3204;
wire     [19:0] PE0_act_regs_1_data_n3224;
wire     [19:0] PE0_act_regs_1_data_n3248;
wire     [19:0] PE0_act_regs_1_data_n3268;
wire     [19:0] PE0_act_regs_1_data_n3292;
wire     [19:0] PE0_act_regs_1_data_n3316;
wire     [19:0] PE0_act_regs_1_data_n3340;
wire     [19:0] PE0_act_regs_1_data_n3364;
wire     [19:0] PE0_act_regs_1_data_n3396;
wire     [19:0] PE0_act_regs_1_data_n3417;
wire     [19:0] PE0_act_regs_1_data_n3437;
wire     [19:0] PE0_act_regs_1_data_n3461;
wire     [19:0] PE0_act_regs_1_data_n3481;
wire     [19:0] PE0_act_regs_1_data_n3505;
wire     [19:0] PE0_act_regs_1_data_n3529;
wire     [19:0] PE0_act_regs_1_data_n3553;
wire     [19:0] PE0_act_regs_1_data_n3577;
wire     [19:0] PE0_act_regs_1_data_n3609;
wire     [19:0] PE0_act_regs_1_data_n3630;
wire     [19:0] PE0_act_regs_1_data_n3650;
wire     [19:0] PE0_act_regs_1_data_n3674;
wire     [19:0] PE0_act_regs_1_data_n3694;
wire     [19:0] PE0_act_regs_1_data_n3718;
wire     [19:0] PE0_act_regs_1_data_n3742;
wire     [19:0] PE0_act_regs_1_data_n3766;
wire     [19:0] PE0_act_regs_1_data_n3790;
wire     [19:0] PE0_act_regs_1_data_n3822;
wire     [19:0] PE0_act_regs_1_data_n3843;
wire     [19:0] PE0_act_regs_1_data_n3863;
wire     [19:0] PE0_act_regs_1_data_n3887;
wire     [19:0] PE0_act_regs_1_data_n3907;
wire     [19:0] PE0_act_regs_1_data_n3931;
wire     [19:0] PE0_act_regs_1_data_n3955;
wire     [19:0] PE0_act_regs_1_data_n3979;
wire     [19:0] PE0_act_regs_1_data_n4003;
wire     [19:0] PE0_act_regs_1_data_n4035;
wire     [19:0] PE0_act_regs_1_data_n4056;
wire     [19:0] PE0_act_regs_1_data_n4076;
wire     [19:0] PE0_act_regs_1_data_n4100;
wire     [19:0] PE0_act_regs_1_data_n4120;
wire     [19:0] PE0_act_regs_1_data_n413;
wire     [19:0] PE0_act_regs_1_data_n4144;
wire     [19:0] PE0_act_regs_1_data_n4168;
wire     [19:0] PE0_act_regs_1_data_n4192;
wire     [19:0] PE0_act_regs_1_data_n4216;
wire     [19:0] PE0_act_regs_1_data_n4248;
wire     [19:0] PE0_act_regs_1_data_n4269;
wire     [19:0] PE0_act_regs_1_data_n4289;
wire     [19:0] PE0_act_regs_1_data_n4313;
wire     [19:0] PE0_act_regs_1_data_n4333;
wire     [19:0] PE0_act_regs_1_data_n4357;
wire     [19:0] PE0_act_regs_1_data_n4381;
wire     [19:0] PE0_act_regs_1_data_n440;
wire     [19:0] PE0_act_regs_1_data_n4405;
wire     [19:0] PE0_act_regs_1_data_n4429;
wire     [19:0] PE0_act_regs_1_data_n465;
wire     [19:0] PE0_act_regs_1_data_n490;
wire     [19:0] PE0_act_regs_1_data_n515;
wire     [19:0] PE0_act_regs_1_data_n540;
wire     [19:0] PE0_act_regs_1_data_n565;
wire     [19:0] PE0_act_regs_1_data_n590;
wire     [19:0] PE0_act_regs_1_data_n615;
wire     [19:0] PE0_act_regs_1_data_n641;
wire     [19:0] PE0_act_regs_1_data_n667;
wire     [19:0] PE0_act_regs_1_data_n692;
wire     [19:0] PE0_act_regs_1_data_n717;
wire     [19:0] PE0_act_regs_1_data_n742;
wire     [19:0] PE0_act_regs_1_data_n767;
wire     [19:0] PE0_act_regs_1_data_n792;
wire            PE0_act_regs_1_wen0;
wire            PE0_act_regs_1_wen1;
wire            PE0_act_regs_1_wen10;
wire            PE0_act_regs_1_wen11;
wire            PE0_act_regs_1_wen12;
wire            PE0_act_regs_1_wen13;
wire            PE0_act_regs_1_wen14;
wire            PE0_act_regs_1_wen15;
wire            PE0_act_regs_1_wen2;
wire            PE0_act_regs_1_wen3;
wire            PE0_act_regs_1_wen4;
wire            PE0_act_regs_1_wen5;
wire            PE0_act_regs_1_wen6;
wire            PE0_act_regs_1_wen7;
wire            PE0_act_regs_1_wen8;
wire            PE0_act_regs_1_wen9;
wire      [3:0] PE0_act_regs_2_addr0;
wire      [3:0] PE0_act_regs_2_addr1;
wire      [3:0] PE0_act_regs_2_addr10;
wire      [3:0] PE0_act_regs_2_addr11;
wire      [3:0] PE0_act_regs_2_addr12;
wire      [3:0] PE0_act_regs_2_addr13;
wire      [3:0] PE0_act_regs_2_addr14;
wire      [3:0] PE0_act_regs_2_addr15;
wire      [3:0] PE0_act_regs_2_addr2;
wire      [3:0] PE0_act_regs_2_addr3;
wire      [3:0] PE0_act_regs_2_addr4;
wire      [3:0] PE0_act_regs_2_addr5;
wire      [3:0] PE0_act_regs_2_addr6;
wire      [3:0] PE0_act_regs_2_addr7;
wire      [3:0] PE0_act_regs_2_addr8;
wire      [3:0] PE0_act_regs_2_addr9;
wire      [3:0] PE0_act_regs_2_addr_n1048;
wire      [3:0] PE0_act_regs_2_addr_n1069;
wire      [3:0] PE0_act_regs_2_addr_n1089;
wire      [3:0] PE0_act_regs_2_addr_n1113;
wire      [3:0] PE0_act_regs_2_addr_n1133;
wire      [3:0] PE0_act_regs_2_addr_n1157;
wire      [3:0] PE0_act_regs_2_addr_n1181;
wire      [3:0] PE0_act_regs_2_addr_n1205;
wire      [3:0] PE0_act_regs_2_addr_n1229;
wire      [3:0] PE0_act_regs_2_addr_n1261;
wire      [3:0] PE0_act_regs_2_addr_n1282;
wire      [3:0] PE0_act_regs_2_addr_n1302;
wire      [3:0] PE0_act_regs_2_addr_n1326;
wire      [3:0] PE0_act_regs_2_addr_n1346;
wire      [3:0] PE0_act_regs_2_addr_n1370;
wire      [3:0] PE0_act_regs_2_addr_n1394;
wire      [3:0] PE0_act_regs_2_addr_n1418;
wire      [3:0] PE0_act_regs_2_addr_n1442;
wire      [3:0] PE0_act_regs_2_addr_n1474;
wire      [3:0] PE0_act_regs_2_addr_n1495;
wire      [3:0] PE0_act_regs_2_addr_n1515;
wire      [3:0] PE0_act_regs_2_addr_n1539;
wire      [3:0] PE0_act_regs_2_addr_n1559;
wire      [3:0] PE0_act_regs_2_addr_n1583;
wire      [3:0] PE0_act_regs_2_addr_n1607;
wire      [3:0] PE0_act_regs_2_addr_n1631;
wire      [3:0] PE0_act_regs_2_addr_n1655;
wire      [3:0] PE0_act_regs_2_addr_n1687;
wire      [3:0] PE0_act_regs_2_addr_n1708;
wire      [3:0] PE0_act_regs_2_addr_n1728;
wire      [3:0] PE0_act_regs_2_addr_n1752;
wire      [3:0] PE0_act_regs_2_addr_n1772;
wire      [3:0] PE0_act_regs_2_addr_n1796;
wire      [3:0] PE0_act_regs_2_addr_n1820;
wire      [3:0] PE0_act_regs_2_addr_n1844;
wire      [3:0] PE0_act_regs_2_addr_n1868;
wire      [3:0] PE0_act_regs_2_addr_n1900;
wire      [3:0] PE0_act_regs_2_addr_n1921;
wire      [3:0] PE0_act_regs_2_addr_n1941;
wire      [3:0] PE0_act_regs_2_addr_n1965;
wire      [3:0] PE0_act_regs_2_addr_n1985;
wire      [3:0] PE0_act_regs_2_addr_n2009;
wire      [3:0] PE0_act_regs_2_addr_n2033;
wire      [3:0] PE0_act_regs_2_addr_n2057;
wire      [3:0] PE0_act_regs_2_addr_n2081;
wire      [3:0] PE0_act_regs_2_addr_n2113;
wire      [3:0] PE0_act_regs_2_addr_n2134;
wire      [3:0] PE0_act_regs_2_addr_n2154;
wire      [3:0] PE0_act_regs_2_addr_n2178;
wire      [3:0] PE0_act_regs_2_addr_n2198;
wire      [3:0] PE0_act_regs_2_addr_n2222;
wire      [3:0] PE0_act_regs_2_addr_n2246;
wire      [3:0] PE0_act_regs_2_addr_n2270;
wire      [3:0] PE0_act_regs_2_addr_n2294;
wire      [3:0] PE0_act_regs_2_addr_n2326;
wire      [3:0] PE0_act_regs_2_addr_n2347;
wire      [3:0] PE0_act_regs_2_addr_n2367;
wire      [3:0] PE0_act_regs_2_addr_n2391;
wire      [3:0] PE0_act_regs_2_addr_n2411;
wire      [3:0] PE0_act_regs_2_addr_n2435;
wire      [3:0] PE0_act_regs_2_addr_n2459;
wire      [3:0] PE0_act_regs_2_addr_n2483;
wire      [3:0] PE0_act_regs_2_addr_n2507;
wire      [3:0] PE0_act_regs_2_addr_n2539;
wire      [3:0] PE0_act_regs_2_addr_n2560;
wire      [3:0] PE0_act_regs_2_addr_n2580;
wire      [3:0] PE0_act_regs_2_addr_n2604;
wire      [3:0] PE0_act_regs_2_addr_n2624;
wire      [3:0] PE0_act_regs_2_addr_n2648;
wire      [3:0] PE0_act_regs_2_addr_n2672;
wire      [3:0] PE0_act_regs_2_addr_n2696;
wire      [3:0] PE0_act_regs_2_addr_n2720;
wire      [3:0] PE0_act_regs_2_addr_n2752;
wire      [3:0] PE0_act_regs_2_addr_n2773;
wire      [3:0] PE0_act_regs_2_addr_n2793;
wire      [3:0] PE0_act_regs_2_addr_n2817;
wire      [3:0] PE0_act_regs_2_addr_n2837;
wire      [3:0] PE0_act_regs_2_addr_n2861;
wire      [3:0] PE0_act_regs_2_addr_n2885;
wire      [3:0] PE0_act_regs_2_addr_n2909;
wire      [3:0] PE0_act_regs_2_addr_n2933;
wire      [3:0] PE0_act_regs_2_addr_n2965;
wire      [3:0] PE0_act_regs_2_addr_n2986;
wire      [3:0] PE0_act_regs_2_addr_n3006;
wire      [3:0] PE0_act_regs_2_addr_n3030;
wire      [3:0] PE0_act_regs_2_addr_n3050;
wire      [3:0] PE0_act_regs_2_addr_n3074;
wire      [3:0] PE0_act_regs_2_addr_n3098;
wire      [3:0] PE0_act_regs_2_addr_n3122;
wire      [3:0] PE0_act_regs_2_addr_n3146;
wire      [3:0] PE0_act_regs_2_addr_n3178;
wire      [3:0] PE0_act_regs_2_addr_n3199;
wire      [3:0] PE0_act_regs_2_addr_n3219;
wire      [3:0] PE0_act_regs_2_addr_n3243;
wire      [3:0] PE0_act_regs_2_addr_n3263;
wire      [3:0] PE0_act_regs_2_addr_n3287;
wire      [3:0] PE0_act_regs_2_addr_n3311;
wire      [3:0] PE0_act_regs_2_addr_n3335;
wire      [3:0] PE0_act_regs_2_addr_n3359;
wire      [3:0] PE0_act_regs_2_addr_n3391;
wire      [3:0] PE0_act_regs_2_addr_n3412;
wire      [3:0] PE0_act_regs_2_addr_n3432;
wire      [3:0] PE0_act_regs_2_addr_n3456;
wire      [3:0] PE0_act_regs_2_addr_n3476;
wire      [3:0] PE0_act_regs_2_addr_n3500;
wire      [3:0] PE0_act_regs_2_addr_n3524;
wire      [3:0] PE0_act_regs_2_addr_n3548;
wire      [3:0] PE0_act_regs_2_addr_n3572;
wire      [3:0] PE0_act_regs_2_addr_n3604;
wire      [3:0] PE0_act_regs_2_addr_n3625;
wire      [3:0] PE0_act_regs_2_addr_n3645;
wire      [3:0] PE0_act_regs_2_addr_n3669;
wire      [3:0] PE0_act_regs_2_addr_n3689;
wire      [3:0] PE0_act_regs_2_addr_n3713;
wire      [3:0] PE0_act_regs_2_addr_n3737;
wire      [3:0] PE0_act_regs_2_addr_n3761;
wire      [3:0] PE0_act_regs_2_addr_n3785;
wire      [3:0] PE0_act_regs_2_addr_n3817;
wire      [3:0] PE0_act_regs_2_addr_n3838;
wire      [3:0] PE0_act_regs_2_addr_n3858;
wire      [3:0] PE0_act_regs_2_addr_n3882;
wire      [3:0] PE0_act_regs_2_addr_n3902;
wire      [3:0] PE0_act_regs_2_addr_n3926;
wire      [3:0] PE0_act_regs_2_addr_n3950;
wire      [3:0] PE0_act_regs_2_addr_n3974;
wire      [3:0] PE0_act_regs_2_addr_n3998;
wire      [3:0] PE0_act_regs_2_addr_n4030;
wire      [3:0] PE0_act_regs_2_addr_n4051;
wire      [3:0] PE0_act_regs_2_addr_n4071;
wire      [3:0] PE0_act_regs_2_addr_n408;
wire      [3:0] PE0_act_regs_2_addr_n4095;
wire      [3:0] PE0_act_regs_2_addr_n4115;
wire      [3:0] PE0_act_regs_2_addr_n4139;
wire      [3:0] PE0_act_regs_2_addr_n4163;
wire      [3:0] PE0_act_regs_2_addr_n4187;
wire      [3:0] PE0_act_regs_2_addr_n4211;
wire      [3:0] PE0_act_regs_2_addr_n4243;
wire      [3:0] PE0_act_regs_2_addr_n4264;
wire      [3:0] PE0_act_regs_2_addr_n4284;
wire      [3:0] PE0_act_regs_2_addr_n4308;
wire      [3:0] PE0_act_regs_2_addr_n4328;
wire      [3:0] PE0_act_regs_2_addr_n435;
wire      [3:0] PE0_act_regs_2_addr_n4352;
wire      [3:0] PE0_act_regs_2_addr_n4376;
wire      [3:0] PE0_act_regs_2_addr_n4400;
wire      [3:0] PE0_act_regs_2_addr_n4424;
wire      [3:0] PE0_act_regs_2_addr_n460;
wire      [3:0] PE0_act_regs_2_addr_n485;
wire      [3:0] PE0_act_regs_2_addr_n510;
wire      [3:0] PE0_act_regs_2_addr_n535;
wire      [3:0] PE0_act_regs_2_addr_n560;
wire      [3:0] PE0_act_regs_2_addr_n585;
wire      [3:0] PE0_act_regs_2_addr_n610;
wire      [3:0] PE0_act_regs_2_addr_n636;
wire      [3:0] PE0_act_regs_2_addr_n662;
wire      [3:0] PE0_act_regs_2_addr_n687;
wire      [3:0] PE0_act_regs_2_addr_n712;
wire      [3:0] PE0_act_regs_2_addr_n737;
wire      [3:0] PE0_act_regs_2_addr_n762;
wire      [3:0] PE0_act_regs_2_addr_n787;
wire     [19:0] PE0_act_regs_2_data0;
wire     [19:0] PE0_act_regs_2_data1;
wire     [19:0] PE0_act_regs_2_data10;
wire     [19:0] PE0_act_regs_2_data11;
wire     [19:0] PE0_act_regs_2_data12;
wire     [19:0] PE0_act_regs_2_data13;
wire     [19:0] PE0_act_regs_2_data14;
wire     [19:0] PE0_act_regs_2_data15;
wire     [19:0] PE0_act_regs_2_data2;
wire     [19:0] PE0_act_regs_2_data3;
wire     [19:0] PE0_act_regs_2_data4;
wire     [19:0] PE0_act_regs_2_data5;
wire     [19:0] PE0_act_regs_2_data6;
wire     [19:0] PE0_act_regs_2_data7;
wire     [19:0] PE0_act_regs_2_data8;
wire     [19:0] PE0_act_regs_2_data9;
wire     [19:0] PE0_act_regs_2_data_n1049;
wire     [19:0] PE0_act_regs_2_data_n1070;
wire     [19:0] PE0_act_regs_2_data_n1090;
wire     [19:0] PE0_act_regs_2_data_n1114;
wire     [19:0] PE0_act_regs_2_data_n1134;
wire     [19:0] PE0_act_regs_2_data_n1158;
wire     [19:0] PE0_act_regs_2_data_n1182;
wire     [19:0] PE0_act_regs_2_data_n1206;
wire     [19:0] PE0_act_regs_2_data_n1230;
wire     [19:0] PE0_act_regs_2_data_n1262;
wire     [19:0] PE0_act_regs_2_data_n1283;
wire     [19:0] PE0_act_regs_2_data_n1303;
wire     [19:0] PE0_act_regs_2_data_n1327;
wire     [19:0] PE0_act_regs_2_data_n1347;
wire     [19:0] PE0_act_regs_2_data_n1371;
wire     [19:0] PE0_act_regs_2_data_n1395;
wire     [19:0] PE0_act_regs_2_data_n1419;
wire     [19:0] PE0_act_regs_2_data_n1443;
wire     [19:0] PE0_act_regs_2_data_n1475;
wire     [19:0] PE0_act_regs_2_data_n1496;
wire     [19:0] PE0_act_regs_2_data_n1516;
wire     [19:0] PE0_act_regs_2_data_n1540;
wire     [19:0] PE0_act_regs_2_data_n1560;
wire     [19:0] PE0_act_regs_2_data_n1584;
wire     [19:0] PE0_act_regs_2_data_n1608;
wire     [19:0] PE0_act_regs_2_data_n1632;
wire     [19:0] PE0_act_regs_2_data_n1656;
wire     [19:0] PE0_act_regs_2_data_n1688;
wire     [19:0] PE0_act_regs_2_data_n1709;
wire     [19:0] PE0_act_regs_2_data_n1729;
wire     [19:0] PE0_act_regs_2_data_n1753;
wire     [19:0] PE0_act_regs_2_data_n1773;
wire     [19:0] PE0_act_regs_2_data_n1797;
wire     [19:0] PE0_act_regs_2_data_n1821;
wire     [19:0] PE0_act_regs_2_data_n1845;
wire     [19:0] PE0_act_regs_2_data_n1869;
wire     [19:0] PE0_act_regs_2_data_n1901;
wire     [19:0] PE0_act_regs_2_data_n1922;
wire     [19:0] PE0_act_regs_2_data_n1942;
wire     [19:0] PE0_act_regs_2_data_n1966;
wire     [19:0] PE0_act_regs_2_data_n1986;
wire     [19:0] PE0_act_regs_2_data_n2010;
wire     [19:0] PE0_act_regs_2_data_n2034;
wire     [19:0] PE0_act_regs_2_data_n2058;
wire     [19:0] PE0_act_regs_2_data_n2082;
wire     [19:0] PE0_act_regs_2_data_n2114;
wire     [19:0] PE0_act_regs_2_data_n2135;
wire     [19:0] PE0_act_regs_2_data_n2155;
wire     [19:0] PE0_act_regs_2_data_n2179;
wire     [19:0] PE0_act_regs_2_data_n2199;
wire     [19:0] PE0_act_regs_2_data_n2223;
wire     [19:0] PE0_act_regs_2_data_n2247;
wire     [19:0] PE0_act_regs_2_data_n2271;
wire     [19:0] PE0_act_regs_2_data_n2295;
wire     [19:0] PE0_act_regs_2_data_n2327;
wire     [19:0] PE0_act_regs_2_data_n2348;
wire     [19:0] PE0_act_regs_2_data_n2368;
wire     [19:0] PE0_act_regs_2_data_n2392;
wire     [19:0] PE0_act_regs_2_data_n2412;
wire     [19:0] PE0_act_regs_2_data_n2436;
wire     [19:0] PE0_act_regs_2_data_n2460;
wire     [19:0] PE0_act_regs_2_data_n2484;
wire     [19:0] PE0_act_regs_2_data_n2508;
wire     [19:0] PE0_act_regs_2_data_n2540;
wire     [19:0] PE0_act_regs_2_data_n2561;
wire     [19:0] PE0_act_regs_2_data_n2581;
wire     [19:0] PE0_act_regs_2_data_n2605;
wire     [19:0] PE0_act_regs_2_data_n2625;
wire     [19:0] PE0_act_regs_2_data_n2649;
wire     [19:0] PE0_act_regs_2_data_n2673;
wire     [19:0] PE0_act_regs_2_data_n2697;
wire     [19:0] PE0_act_regs_2_data_n2721;
wire     [19:0] PE0_act_regs_2_data_n2753;
wire     [19:0] PE0_act_regs_2_data_n2774;
wire     [19:0] PE0_act_regs_2_data_n2794;
wire     [19:0] PE0_act_regs_2_data_n2818;
wire     [19:0] PE0_act_regs_2_data_n2838;
wire     [19:0] PE0_act_regs_2_data_n2862;
wire     [19:0] PE0_act_regs_2_data_n2886;
wire     [19:0] PE0_act_regs_2_data_n2910;
wire     [19:0] PE0_act_regs_2_data_n2934;
wire     [19:0] PE0_act_regs_2_data_n2966;
wire     [19:0] PE0_act_regs_2_data_n2987;
wire     [19:0] PE0_act_regs_2_data_n3007;
wire     [19:0] PE0_act_regs_2_data_n3031;
wire     [19:0] PE0_act_regs_2_data_n3051;
wire     [19:0] PE0_act_regs_2_data_n3075;
wire     [19:0] PE0_act_regs_2_data_n3099;
wire     [19:0] PE0_act_regs_2_data_n3123;
wire     [19:0] PE0_act_regs_2_data_n3147;
wire     [19:0] PE0_act_regs_2_data_n3179;
wire     [19:0] PE0_act_regs_2_data_n3200;
wire     [19:0] PE0_act_regs_2_data_n3220;
wire     [19:0] PE0_act_regs_2_data_n3244;
wire     [19:0] PE0_act_regs_2_data_n3264;
wire     [19:0] PE0_act_regs_2_data_n3288;
wire     [19:0] PE0_act_regs_2_data_n3312;
wire     [19:0] PE0_act_regs_2_data_n3336;
wire     [19:0] PE0_act_regs_2_data_n3360;
wire     [19:0] PE0_act_regs_2_data_n3392;
wire     [19:0] PE0_act_regs_2_data_n3413;
wire     [19:0] PE0_act_regs_2_data_n3433;
wire     [19:0] PE0_act_regs_2_data_n3457;
wire     [19:0] PE0_act_regs_2_data_n3477;
wire     [19:0] PE0_act_regs_2_data_n3501;
wire     [19:0] PE0_act_regs_2_data_n3525;
wire     [19:0] PE0_act_regs_2_data_n3549;
wire     [19:0] PE0_act_regs_2_data_n3573;
wire     [19:0] PE0_act_regs_2_data_n3605;
wire     [19:0] PE0_act_regs_2_data_n3626;
wire     [19:0] PE0_act_regs_2_data_n3646;
wire     [19:0] PE0_act_regs_2_data_n3670;
wire     [19:0] PE0_act_regs_2_data_n3690;
wire     [19:0] PE0_act_regs_2_data_n3714;
wire     [19:0] PE0_act_regs_2_data_n3738;
wire     [19:0] PE0_act_regs_2_data_n3762;
wire     [19:0] PE0_act_regs_2_data_n3786;
wire     [19:0] PE0_act_regs_2_data_n3818;
wire     [19:0] PE0_act_regs_2_data_n3839;
wire     [19:0] PE0_act_regs_2_data_n3859;
wire     [19:0] PE0_act_regs_2_data_n3883;
wire     [19:0] PE0_act_regs_2_data_n3903;
wire     [19:0] PE0_act_regs_2_data_n3927;
wire     [19:0] PE0_act_regs_2_data_n3951;
wire     [19:0] PE0_act_regs_2_data_n3975;
wire     [19:0] PE0_act_regs_2_data_n3999;
wire     [19:0] PE0_act_regs_2_data_n4031;
wire     [19:0] PE0_act_regs_2_data_n4052;
wire     [19:0] PE0_act_regs_2_data_n4072;
wire     [19:0] PE0_act_regs_2_data_n409;
wire     [19:0] PE0_act_regs_2_data_n4096;
wire     [19:0] PE0_act_regs_2_data_n4116;
wire     [19:0] PE0_act_regs_2_data_n4140;
wire     [19:0] PE0_act_regs_2_data_n4164;
wire     [19:0] PE0_act_regs_2_data_n4188;
wire     [19:0] PE0_act_regs_2_data_n4212;
wire     [19:0] PE0_act_regs_2_data_n4244;
wire     [19:0] PE0_act_regs_2_data_n4265;
wire     [19:0] PE0_act_regs_2_data_n4285;
wire     [19:0] PE0_act_regs_2_data_n4309;
wire     [19:0] PE0_act_regs_2_data_n4329;
wire     [19:0] PE0_act_regs_2_data_n4353;
wire     [19:0] PE0_act_regs_2_data_n436;
wire     [19:0] PE0_act_regs_2_data_n4377;
wire     [19:0] PE0_act_regs_2_data_n4401;
wire     [19:0] PE0_act_regs_2_data_n4425;
wire     [19:0] PE0_act_regs_2_data_n461;
wire     [19:0] PE0_act_regs_2_data_n486;
wire     [19:0] PE0_act_regs_2_data_n511;
wire     [19:0] PE0_act_regs_2_data_n536;
wire     [19:0] PE0_act_regs_2_data_n561;
wire     [19:0] PE0_act_regs_2_data_n586;
wire     [19:0] PE0_act_regs_2_data_n611;
wire     [19:0] PE0_act_regs_2_data_n637;
wire     [19:0] PE0_act_regs_2_data_n663;
wire     [19:0] PE0_act_regs_2_data_n688;
wire     [19:0] PE0_act_regs_2_data_n713;
wire     [19:0] PE0_act_regs_2_data_n738;
wire     [19:0] PE0_act_regs_2_data_n763;
wire     [19:0] PE0_act_regs_2_data_n788;
wire            PE0_act_regs_2_wen0;
wire            PE0_act_regs_2_wen1;
wire            PE0_act_regs_2_wen10;
wire            PE0_act_regs_2_wen11;
wire            PE0_act_regs_2_wen12;
wire            PE0_act_regs_2_wen13;
wire            PE0_act_regs_2_wen14;
wire            PE0_act_regs_2_wen15;
wire            PE0_act_regs_2_wen2;
wire            PE0_act_regs_2_wen3;
wire            PE0_act_regs_2_wen4;
wire            PE0_act_regs_2_wen5;
wire            PE0_act_regs_2_wen6;
wire            PE0_act_regs_2_wen7;
wire            PE0_act_regs_2_wen8;
wire            PE0_act_regs_2_wen9;
wire      [3:0] PE0_act_regs_3_addr0;
wire      [3:0] PE0_act_regs_3_addr1;
wire      [3:0] PE0_act_regs_3_addr10;
wire      [3:0] PE0_act_regs_3_addr11;
wire      [3:0] PE0_act_regs_3_addr12;
wire      [3:0] PE0_act_regs_3_addr13;
wire      [3:0] PE0_act_regs_3_addr14;
wire      [3:0] PE0_act_regs_3_addr15;
wire      [3:0] PE0_act_regs_3_addr2;
wire      [3:0] PE0_act_regs_3_addr3;
wire      [3:0] PE0_act_regs_3_addr4;
wire      [3:0] PE0_act_regs_3_addr5;
wire      [3:0] PE0_act_regs_3_addr6;
wire      [3:0] PE0_act_regs_3_addr7;
wire      [3:0] PE0_act_regs_3_addr8;
wire      [3:0] PE0_act_regs_3_addr9;
wire      [3:0] PE0_act_regs_3_addr_n1044;
wire      [3:0] PE0_act_regs_3_addr_n1065;
wire      [3:0] PE0_act_regs_3_addr_n1085;
wire      [3:0] PE0_act_regs_3_addr_n1109;
wire      [3:0] PE0_act_regs_3_addr_n1129;
wire      [3:0] PE0_act_regs_3_addr_n1153;
wire      [3:0] PE0_act_regs_3_addr_n1177;
wire      [3:0] PE0_act_regs_3_addr_n1201;
wire      [3:0] PE0_act_regs_3_addr_n1225;
wire      [3:0] PE0_act_regs_3_addr_n1257;
wire      [3:0] PE0_act_regs_3_addr_n1278;
wire      [3:0] PE0_act_regs_3_addr_n1298;
wire      [3:0] PE0_act_regs_3_addr_n1322;
wire      [3:0] PE0_act_regs_3_addr_n1342;
wire      [3:0] PE0_act_regs_3_addr_n1366;
wire      [3:0] PE0_act_regs_3_addr_n1390;
wire      [3:0] PE0_act_regs_3_addr_n1414;
wire      [3:0] PE0_act_regs_3_addr_n1438;
wire      [3:0] PE0_act_regs_3_addr_n1470;
wire      [3:0] PE0_act_regs_3_addr_n1491;
wire      [3:0] PE0_act_regs_3_addr_n1511;
wire      [3:0] PE0_act_regs_3_addr_n1535;
wire      [3:0] PE0_act_regs_3_addr_n1555;
wire      [3:0] PE0_act_regs_3_addr_n1579;
wire      [3:0] PE0_act_regs_3_addr_n1603;
wire      [3:0] PE0_act_regs_3_addr_n1627;
wire      [3:0] PE0_act_regs_3_addr_n1651;
wire      [3:0] PE0_act_regs_3_addr_n1683;
wire      [3:0] PE0_act_regs_3_addr_n1704;
wire      [3:0] PE0_act_regs_3_addr_n1724;
wire      [3:0] PE0_act_regs_3_addr_n1748;
wire      [3:0] PE0_act_regs_3_addr_n1768;
wire      [3:0] PE0_act_regs_3_addr_n1792;
wire      [3:0] PE0_act_regs_3_addr_n1816;
wire      [3:0] PE0_act_regs_3_addr_n1840;
wire      [3:0] PE0_act_regs_3_addr_n1864;
wire      [3:0] PE0_act_regs_3_addr_n1896;
wire      [3:0] PE0_act_regs_3_addr_n1917;
wire      [3:0] PE0_act_regs_3_addr_n1937;
wire      [3:0] PE0_act_regs_3_addr_n1961;
wire      [3:0] PE0_act_regs_3_addr_n1981;
wire      [3:0] PE0_act_regs_3_addr_n2005;
wire      [3:0] PE0_act_regs_3_addr_n2029;
wire      [3:0] PE0_act_regs_3_addr_n2053;
wire      [3:0] PE0_act_regs_3_addr_n2077;
wire      [3:0] PE0_act_regs_3_addr_n2109;
wire      [3:0] PE0_act_regs_3_addr_n2130;
wire      [3:0] PE0_act_regs_3_addr_n2150;
wire      [3:0] PE0_act_regs_3_addr_n2174;
wire      [3:0] PE0_act_regs_3_addr_n2194;
wire      [3:0] PE0_act_regs_3_addr_n2218;
wire      [3:0] PE0_act_regs_3_addr_n2242;
wire      [3:0] PE0_act_regs_3_addr_n2266;
wire      [3:0] PE0_act_regs_3_addr_n2290;
wire      [3:0] PE0_act_regs_3_addr_n2322;
wire      [3:0] PE0_act_regs_3_addr_n2343;
wire      [3:0] PE0_act_regs_3_addr_n2363;
wire      [3:0] PE0_act_regs_3_addr_n2387;
wire      [3:0] PE0_act_regs_3_addr_n2407;
wire      [3:0] PE0_act_regs_3_addr_n2431;
wire      [3:0] PE0_act_regs_3_addr_n2455;
wire      [3:0] PE0_act_regs_3_addr_n2479;
wire      [3:0] PE0_act_regs_3_addr_n2503;
wire      [3:0] PE0_act_regs_3_addr_n2535;
wire      [3:0] PE0_act_regs_3_addr_n2556;
wire      [3:0] PE0_act_regs_3_addr_n2576;
wire      [3:0] PE0_act_regs_3_addr_n2600;
wire      [3:0] PE0_act_regs_3_addr_n2620;
wire      [3:0] PE0_act_regs_3_addr_n2644;
wire      [3:0] PE0_act_regs_3_addr_n2668;
wire      [3:0] PE0_act_regs_3_addr_n2692;
wire      [3:0] PE0_act_regs_3_addr_n2716;
wire      [3:0] PE0_act_regs_3_addr_n2748;
wire      [3:0] PE0_act_regs_3_addr_n2769;
wire      [3:0] PE0_act_regs_3_addr_n2789;
wire      [3:0] PE0_act_regs_3_addr_n2813;
wire      [3:0] PE0_act_regs_3_addr_n2833;
wire      [3:0] PE0_act_regs_3_addr_n2857;
wire      [3:0] PE0_act_regs_3_addr_n2881;
wire      [3:0] PE0_act_regs_3_addr_n2905;
wire      [3:0] PE0_act_regs_3_addr_n2929;
wire      [3:0] PE0_act_regs_3_addr_n2961;
wire      [3:0] PE0_act_regs_3_addr_n2982;
wire      [3:0] PE0_act_regs_3_addr_n3002;
wire      [3:0] PE0_act_regs_3_addr_n3026;
wire      [3:0] PE0_act_regs_3_addr_n3046;
wire      [3:0] PE0_act_regs_3_addr_n3070;
wire      [3:0] PE0_act_regs_3_addr_n3094;
wire      [3:0] PE0_act_regs_3_addr_n3118;
wire      [3:0] PE0_act_regs_3_addr_n3142;
wire      [3:0] PE0_act_regs_3_addr_n3174;
wire      [3:0] PE0_act_regs_3_addr_n3195;
wire      [3:0] PE0_act_regs_3_addr_n3215;
wire      [3:0] PE0_act_regs_3_addr_n3239;
wire      [3:0] PE0_act_regs_3_addr_n3259;
wire      [3:0] PE0_act_regs_3_addr_n3283;
wire      [3:0] PE0_act_regs_3_addr_n3307;
wire      [3:0] PE0_act_regs_3_addr_n3331;
wire      [3:0] PE0_act_regs_3_addr_n3355;
wire      [3:0] PE0_act_regs_3_addr_n3387;
wire      [3:0] PE0_act_regs_3_addr_n3408;
wire      [3:0] PE0_act_regs_3_addr_n3428;
wire      [3:0] PE0_act_regs_3_addr_n3452;
wire      [3:0] PE0_act_regs_3_addr_n3472;
wire      [3:0] PE0_act_regs_3_addr_n3496;
wire      [3:0] PE0_act_regs_3_addr_n3520;
wire      [3:0] PE0_act_regs_3_addr_n3544;
wire      [3:0] PE0_act_regs_3_addr_n3568;
wire      [3:0] PE0_act_regs_3_addr_n3600;
wire      [3:0] PE0_act_regs_3_addr_n3621;
wire      [3:0] PE0_act_regs_3_addr_n3641;
wire      [3:0] PE0_act_regs_3_addr_n3665;
wire      [3:0] PE0_act_regs_3_addr_n3685;
wire      [3:0] PE0_act_regs_3_addr_n3709;
wire      [3:0] PE0_act_regs_3_addr_n3733;
wire      [3:0] PE0_act_regs_3_addr_n3757;
wire      [3:0] PE0_act_regs_3_addr_n3781;
wire      [3:0] PE0_act_regs_3_addr_n3813;
wire      [3:0] PE0_act_regs_3_addr_n3834;
wire      [3:0] PE0_act_regs_3_addr_n3854;
wire      [3:0] PE0_act_regs_3_addr_n3878;
wire      [3:0] PE0_act_regs_3_addr_n3898;
wire      [3:0] PE0_act_regs_3_addr_n3922;
wire      [3:0] PE0_act_regs_3_addr_n3946;
wire      [3:0] PE0_act_regs_3_addr_n3970;
wire      [3:0] PE0_act_regs_3_addr_n3994;
wire      [3:0] PE0_act_regs_3_addr_n4026;
wire      [3:0] PE0_act_regs_3_addr_n404;
wire      [3:0] PE0_act_regs_3_addr_n4047;
wire      [3:0] PE0_act_regs_3_addr_n4067;
wire      [3:0] PE0_act_regs_3_addr_n4091;
wire      [3:0] PE0_act_regs_3_addr_n4111;
wire      [3:0] PE0_act_regs_3_addr_n4135;
wire      [3:0] PE0_act_regs_3_addr_n4159;
wire      [3:0] PE0_act_regs_3_addr_n4183;
wire      [3:0] PE0_act_regs_3_addr_n4207;
wire      [3:0] PE0_act_regs_3_addr_n4239;
wire      [3:0] PE0_act_regs_3_addr_n4260;
wire      [3:0] PE0_act_regs_3_addr_n4280;
wire      [3:0] PE0_act_regs_3_addr_n4304;
wire      [3:0] PE0_act_regs_3_addr_n431;
wire      [3:0] PE0_act_regs_3_addr_n4324;
wire      [3:0] PE0_act_regs_3_addr_n4348;
wire      [3:0] PE0_act_regs_3_addr_n4372;
wire      [3:0] PE0_act_regs_3_addr_n4396;
wire      [3:0] PE0_act_regs_3_addr_n4420;
wire      [3:0] PE0_act_regs_3_addr_n456;
wire      [3:0] PE0_act_regs_3_addr_n481;
wire      [3:0] PE0_act_regs_3_addr_n506;
wire      [3:0] PE0_act_regs_3_addr_n531;
wire      [3:0] PE0_act_regs_3_addr_n556;
wire      [3:0] PE0_act_regs_3_addr_n581;
wire      [3:0] PE0_act_regs_3_addr_n606;
wire      [3:0] PE0_act_regs_3_addr_n632;
wire      [3:0] PE0_act_regs_3_addr_n658;
wire      [3:0] PE0_act_regs_3_addr_n683;
wire      [3:0] PE0_act_regs_3_addr_n708;
wire      [3:0] PE0_act_regs_3_addr_n733;
wire      [3:0] PE0_act_regs_3_addr_n758;
wire      [3:0] PE0_act_regs_3_addr_n783;
wire     [19:0] PE0_act_regs_3_data0;
wire     [19:0] PE0_act_regs_3_data1;
wire     [19:0] PE0_act_regs_3_data10;
wire     [19:0] PE0_act_regs_3_data11;
wire     [19:0] PE0_act_regs_3_data12;
wire     [19:0] PE0_act_regs_3_data13;
wire     [19:0] PE0_act_regs_3_data14;
wire     [19:0] PE0_act_regs_3_data15;
wire     [19:0] PE0_act_regs_3_data2;
wire     [19:0] PE0_act_regs_3_data3;
wire     [19:0] PE0_act_regs_3_data4;
wire     [19:0] PE0_act_regs_3_data5;
wire     [19:0] PE0_act_regs_3_data6;
wire     [19:0] PE0_act_regs_3_data7;
wire     [19:0] PE0_act_regs_3_data8;
wire     [19:0] PE0_act_regs_3_data9;
wire     [19:0] PE0_act_regs_3_data_n1045;
wire     [19:0] PE0_act_regs_3_data_n1066;
wire     [19:0] PE0_act_regs_3_data_n1086;
wire     [19:0] PE0_act_regs_3_data_n1110;
wire     [19:0] PE0_act_regs_3_data_n1130;
wire     [19:0] PE0_act_regs_3_data_n1154;
wire     [19:0] PE0_act_regs_3_data_n1178;
wire     [19:0] PE0_act_regs_3_data_n1202;
wire     [19:0] PE0_act_regs_3_data_n1226;
wire     [19:0] PE0_act_regs_3_data_n1258;
wire     [19:0] PE0_act_regs_3_data_n1279;
wire     [19:0] PE0_act_regs_3_data_n1299;
wire     [19:0] PE0_act_regs_3_data_n1323;
wire     [19:0] PE0_act_regs_3_data_n1343;
wire     [19:0] PE0_act_regs_3_data_n1367;
wire     [19:0] PE0_act_regs_3_data_n1391;
wire     [19:0] PE0_act_regs_3_data_n1415;
wire     [19:0] PE0_act_regs_3_data_n1439;
wire     [19:0] PE0_act_regs_3_data_n1471;
wire     [19:0] PE0_act_regs_3_data_n1492;
wire     [19:0] PE0_act_regs_3_data_n1512;
wire     [19:0] PE0_act_regs_3_data_n1536;
wire     [19:0] PE0_act_regs_3_data_n1556;
wire     [19:0] PE0_act_regs_3_data_n1580;
wire     [19:0] PE0_act_regs_3_data_n1604;
wire     [19:0] PE0_act_regs_3_data_n1628;
wire     [19:0] PE0_act_regs_3_data_n1652;
wire     [19:0] PE0_act_regs_3_data_n1684;
wire     [19:0] PE0_act_regs_3_data_n1705;
wire     [19:0] PE0_act_regs_3_data_n1725;
wire     [19:0] PE0_act_regs_3_data_n1749;
wire     [19:0] PE0_act_regs_3_data_n1769;
wire     [19:0] PE0_act_regs_3_data_n1793;
wire     [19:0] PE0_act_regs_3_data_n1817;
wire     [19:0] PE0_act_regs_3_data_n1841;
wire     [19:0] PE0_act_regs_3_data_n1865;
wire     [19:0] PE0_act_regs_3_data_n1897;
wire     [19:0] PE0_act_regs_3_data_n1918;
wire     [19:0] PE0_act_regs_3_data_n1938;
wire     [19:0] PE0_act_regs_3_data_n1962;
wire     [19:0] PE0_act_regs_3_data_n1982;
wire     [19:0] PE0_act_regs_3_data_n2006;
wire     [19:0] PE0_act_regs_3_data_n2030;
wire     [19:0] PE0_act_regs_3_data_n2054;
wire     [19:0] PE0_act_regs_3_data_n2078;
wire     [19:0] PE0_act_regs_3_data_n2110;
wire     [19:0] PE0_act_regs_3_data_n2131;
wire     [19:0] PE0_act_regs_3_data_n2151;
wire     [19:0] PE0_act_regs_3_data_n2175;
wire     [19:0] PE0_act_regs_3_data_n2195;
wire     [19:0] PE0_act_regs_3_data_n2219;
wire     [19:0] PE0_act_regs_3_data_n2243;
wire     [19:0] PE0_act_regs_3_data_n2267;
wire     [19:0] PE0_act_regs_3_data_n2291;
wire     [19:0] PE0_act_regs_3_data_n2323;
wire     [19:0] PE0_act_regs_3_data_n2344;
wire     [19:0] PE0_act_regs_3_data_n2364;
wire     [19:0] PE0_act_regs_3_data_n2388;
wire     [19:0] PE0_act_regs_3_data_n2408;
wire     [19:0] PE0_act_regs_3_data_n2432;
wire     [19:0] PE0_act_regs_3_data_n2456;
wire     [19:0] PE0_act_regs_3_data_n2480;
wire     [19:0] PE0_act_regs_3_data_n2504;
wire     [19:0] PE0_act_regs_3_data_n2536;
wire     [19:0] PE0_act_regs_3_data_n2557;
wire     [19:0] PE0_act_regs_3_data_n2577;
wire     [19:0] PE0_act_regs_3_data_n2601;
wire     [19:0] PE0_act_regs_3_data_n2621;
wire     [19:0] PE0_act_regs_3_data_n2645;
wire     [19:0] PE0_act_regs_3_data_n2669;
wire     [19:0] PE0_act_regs_3_data_n2693;
wire     [19:0] PE0_act_regs_3_data_n2717;
wire     [19:0] PE0_act_regs_3_data_n2749;
wire     [19:0] PE0_act_regs_3_data_n2770;
wire     [19:0] PE0_act_regs_3_data_n2790;
wire     [19:0] PE0_act_regs_3_data_n2814;
wire     [19:0] PE0_act_regs_3_data_n2834;
wire     [19:0] PE0_act_regs_3_data_n2858;
wire     [19:0] PE0_act_regs_3_data_n2882;
wire     [19:0] PE0_act_regs_3_data_n2906;
wire     [19:0] PE0_act_regs_3_data_n2930;
wire     [19:0] PE0_act_regs_3_data_n2962;
wire     [19:0] PE0_act_regs_3_data_n2983;
wire     [19:0] PE0_act_regs_3_data_n3003;
wire     [19:0] PE0_act_regs_3_data_n3027;
wire     [19:0] PE0_act_regs_3_data_n3047;
wire     [19:0] PE0_act_regs_3_data_n3071;
wire     [19:0] PE0_act_regs_3_data_n3095;
wire     [19:0] PE0_act_regs_3_data_n3119;
wire     [19:0] PE0_act_regs_3_data_n3143;
wire     [19:0] PE0_act_regs_3_data_n3175;
wire     [19:0] PE0_act_regs_3_data_n3196;
wire     [19:0] PE0_act_regs_3_data_n3216;
wire     [19:0] PE0_act_regs_3_data_n3240;
wire     [19:0] PE0_act_regs_3_data_n3260;
wire     [19:0] PE0_act_regs_3_data_n3284;
wire     [19:0] PE0_act_regs_3_data_n3308;
wire     [19:0] PE0_act_regs_3_data_n3332;
wire     [19:0] PE0_act_regs_3_data_n3356;
wire     [19:0] PE0_act_regs_3_data_n3388;
wire     [19:0] PE0_act_regs_3_data_n3409;
wire     [19:0] PE0_act_regs_3_data_n3429;
wire     [19:0] PE0_act_regs_3_data_n3453;
wire     [19:0] PE0_act_regs_3_data_n3473;
wire     [19:0] PE0_act_regs_3_data_n3497;
wire     [19:0] PE0_act_regs_3_data_n3521;
wire     [19:0] PE0_act_regs_3_data_n3545;
wire     [19:0] PE0_act_regs_3_data_n3569;
wire     [19:0] PE0_act_regs_3_data_n3601;
wire     [19:0] PE0_act_regs_3_data_n3622;
wire     [19:0] PE0_act_regs_3_data_n3642;
wire     [19:0] PE0_act_regs_3_data_n3666;
wire     [19:0] PE0_act_regs_3_data_n3686;
wire     [19:0] PE0_act_regs_3_data_n3710;
wire     [19:0] PE0_act_regs_3_data_n3734;
wire     [19:0] PE0_act_regs_3_data_n3758;
wire     [19:0] PE0_act_regs_3_data_n3782;
wire     [19:0] PE0_act_regs_3_data_n3814;
wire     [19:0] PE0_act_regs_3_data_n3835;
wire     [19:0] PE0_act_regs_3_data_n3855;
wire     [19:0] PE0_act_regs_3_data_n3879;
wire     [19:0] PE0_act_regs_3_data_n3899;
wire     [19:0] PE0_act_regs_3_data_n3923;
wire     [19:0] PE0_act_regs_3_data_n3947;
wire     [19:0] PE0_act_regs_3_data_n3971;
wire     [19:0] PE0_act_regs_3_data_n3995;
wire     [19:0] PE0_act_regs_3_data_n4027;
wire     [19:0] PE0_act_regs_3_data_n4048;
wire     [19:0] PE0_act_regs_3_data_n405;
wire     [19:0] PE0_act_regs_3_data_n4068;
wire     [19:0] PE0_act_regs_3_data_n4092;
wire     [19:0] PE0_act_regs_3_data_n4112;
wire     [19:0] PE0_act_regs_3_data_n4136;
wire     [19:0] PE0_act_regs_3_data_n4160;
wire     [19:0] PE0_act_regs_3_data_n4184;
wire     [19:0] PE0_act_regs_3_data_n4208;
wire     [19:0] PE0_act_regs_3_data_n4240;
wire     [19:0] PE0_act_regs_3_data_n4261;
wire     [19:0] PE0_act_regs_3_data_n4281;
wire     [19:0] PE0_act_regs_3_data_n4305;
wire     [19:0] PE0_act_regs_3_data_n432;
wire     [19:0] PE0_act_regs_3_data_n4325;
wire     [19:0] PE0_act_regs_3_data_n4349;
wire     [19:0] PE0_act_regs_3_data_n4373;
wire     [19:0] PE0_act_regs_3_data_n4397;
wire     [19:0] PE0_act_regs_3_data_n4421;
wire     [19:0] PE0_act_regs_3_data_n457;
wire     [19:0] PE0_act_regs_3_data_n482;
wire     [19:0] PE0_act_regs_3_data_n507;
wire     [19:0] PE0_act_regs_3_data_n532;
wire     [19:0] PE0_act_regs_3_data_n557;
wire     [19:0] PE0_act_regs_3_data_n582;
wire     [19:0] PE0_act_regs_3_data_n607;
wire     [19:0] PE0_act_regs_3_data_n633;
wire     [19:0] PE0_act_regs_3_data_n659;
wire     [19:0] PE0_act_regs_3_data_n684;
wire     [19:0] PE0_act_regs_3_data_n709;
wire     [19:0] PE0_act_regs_3_data_n734;
wire     [19:0] PE0_act_regs_3_data_n759;
wire     [19:0] PE0_act_regs_3_data_n784;
wire            PE0_act_regs_3_wen0;
wire            PE0_act_regs_3_wen1;
wire            PE0_act_regs_3_wen10;
wire            PE0_act_regs_3_wen11;
wire            PE0_act_regs_3_wen12;
wire            PE0_act_regs_3_wen13;
wire            PE0_act_regs_3_wen14;
wire            PE0_act_regs_3_wen15;
wire            PE0_act_regs_3_wen2;
wire            PE0_act_regs_3_wen3;
wire            PE0_act_regs_3_wen4;
wire            PE0_act_regs_3_wen5;
wire            PE0_act_regs_3_wen6;
wire            PE0_act_regs_3_wen7;
wire            PE0_act_regs_3_wen8;
wire            PE0_act_regs_3_wen9;
wire     [19:0] PE0_core_act_vector_0;
wire     [19:0] PE0_core_act_vector_1;
wire     [19:0] PE0_core_act_vector_10;
wire     [19:0] PE0_core_act_vector_11;
wire     [19:0] PE0_core_act_vector_12;
wire     [19:0] PE0_core_act_vector_13;
wire     [19:0] PE0_core_act_vector_14;
wire     [19:0] PE0_core_act_vector_15;
wire     [19:0] PE0_core_act_vector_2;
wire     [19:0] PE0_core_act_vector_3;
wire     [19:0] PE0_core_act_vector_4;
wire     [19:0] PE0_core_act_vector_5;
wire     [19:0] PE0_core_act_vector_6;
wire     [19:0] PE0_core_act_vector_7;
wire     [19:0] PE0_core_act_vector_8;
wire     [19:0] PE0_core_act_vector_9;
wire     [19:0] __ILA_pe_act_acc_decode__;
wire            __ILA_pe_act_decode_of_PE0_ACT_STORE_BUFFER__;
wire            __ILA_pe_act_decode_of_PE0_CONFIG_ACT_MNGR__;
wire            __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_0_15__;
wire            __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_16_31__;
wire            __ILA_pe_act_decode_of_PE0_act_child_done_sent__;
wire            __ILA_pe_act_decode_of_PE0_act_child_initiate__;
wire            __ILA_pe_act_decode_of_PE0_act_child_op_copy__;
wire            __ILA_pe_act_decode_of_PE0_act_child_op_eadd__;
wire            __ILA_pe_act_decode_of_PE0_act_child_op_emul__;
wire            __ILA_pe_act_decode_of_PE0_act_child_op_inpe__;
wire            __ILA_pe_act_decode_of_PE0_act_child_op_load__;
wire            __ILA_pe_act_decode_of_PE0_act_child_op_load_zero__;
wire            __ILA_pe_act_decode_of_PE0_act_child_op_onex__;
wire            __ILA_pe_act_decode_of_PE0_act_child_op_outgb__;
wire            __ILA_pe_act_decode_of_PE0_act_child_op_relu__;
wire            __ILA_pe_act_decode_of_PE0_act_child_op_sigm__;
wire            __ILA_pe_act_decode_of_PE0_act_child_op_store__;
wire            __ILA_pe_act_decode_of_PE0_act_child_op_tanh__;
wire            __ILA_pe_act_decode_of_PE0_act_child_out_sent__;
wire            __ILA_pe_act_decode_of_PE0_act_child_reg_store__;
wire     [19:0] __ILA_pe_act_grant__;
wire            __ILA_pe_act_valid__;
wire            act_start;
wire            act_start_valid;
wire     [23:0] addr;
wire            axi_rw;
wire            bv_1_0_n32;
wire            bv_1_1_n0;
wire     [19:0] bv_20_0_n419;
wire     [23:0] bv_24_0_n391;
wire     [23:0] bv_24_8388624_n2;
wire     [23:0] bv_24_8388640_n9;
wire     [23:0] bv_24_8388656_n15;
wire     [23:0] bv_24_9437184_n21;
wire     [23:0] bv_24_9437680_n25;
wire     [26:0] bv_27_0_n393;
wire      [1:0] bv_2_0_n41;
wire      [1:0] bv_2_1_n45;
wire      [1:0] bv_2_2_n224;
wire      [1:0] bv_2_3_n399;
wire     [31:0] bv_32_0_n388;
wire     [31:0] bv_32_10_n368;
wire     [31:0] bv_32_11_n366;
wire     [31:0] bv_32_12_n364;
wire     [31:0] bv_32_13_n362;
wire     [31:0] bv_32_14_n360;
wire     [31:0] bv_32_15_n358;
wire     [31:0] bv_32_1_n386;
wire     [31:0] bv_32_2_n384;
wire     [31:0] bv_32_3_n382;
wire     [31:0] bv_32_4_n380;
wire     [31:0] bv_32_5_n378;
wire     [31:0] bv_32_6_n376;
wire     [31:0] bv_32_7_n374;
wire     [31:0] bv_32_8_n372;
wire     [31:0] bv_32_9437184_n356;
wire     [31:0] bv_32_9_n370;
wire      [3:0] bv_4_0_n402;
wire      [3:0] bv_4_10_n202;
wire      [3:0] bv_4_11_n208;
wire      [3:0] bv_4_12_n214;
wire      [3:0] bv_4_13_n220;
wire      [3:0] bv_4_14_n429;
wire      [3:0] bv_4_15_n401;
wire      [3:0] bv_4_1_n145;
wire      [3:0] bv_4_2_n160;
wire      [3:0] bv_4_3_n166;
wire      [3:0] bv_4_4_n176;
wire      [3:0] bv_4_5_n656;
wire      [3:0] bv_4_6_n630;
wire      [3:0] bv_4_7_n184;
wire      [3:0] bv_4_8_n190;
wire      [3:0] bv_4_9_n196;
wire      [5:0] bv_6_0_n110;
wire      [5:0] bv_6_10_n90;
wire      [5:0] bv_6_11_n88;
wire      [5:0] bv_6_12_n86;
wire      [5:0] bv_6_13_n84;
wire      [5:0] bv_6_14_n82;
wire      [5:0] bv_6_15_n80;
wire      [5:0] bv_6_16_n78;
wire      [5:0] bv_6_17_n76;
wire      [5:0] bv_6_18_n74;
wire      [5:0] bv_6_19_n72;
wire      [5:0] bv_6_1_n108;
wire      [5:0] bv_6_20_n70;
wire      [5:0] bv_6_21_n68;
wire      [5:0] bv_6_22_n66;
wire      [5:0] bv_6_23_n64;
wire      [5:0] bv_6_24_n62;
wire      [5:0] bv_6_25_n60;
wire      [5:0] bv_6_26_n58;
wire      [5:0] bv_6_27_n56;
wire      [5:0] bv_6_28_n54;
wire      [5:0] bv_6_29_n52;
wire      [5:0] bv_6_2_n106;
wire      [5:0] bv_6_30_n50;
wire      [5:0] bv_6_31_n48;
wire      [5:0] bv_6_3_n104;
wire      [5:0] bv_6_4_n102;
wire      [5:0] bv_6_5_n100;
wire      [5:0] bv_6_6_n98;
wire      [5:0] bv_6_7_n96;
wire      [5:0] bv_6_8_n94;
wire      [5:0] bv_6_9_n92;
wire      [7:0] bv_8_0_n354;
wire      [7:0] bv_8_1_n248;
wire            clk;
wire      [7:0] data_in_0;
wire      [7:0] data_in_1;
wire      [7:0] data_in_10;
wire      [7:0] data_in_11;
wire      [7:0] data_in_12;
wire      [7:0] data_in_13;
wire      [7:0] data_in_14;
wire      [7:0] data_in_15;
wire      [7:0] data_in_2;
wire      [7:0] data_in_3;
wire      [7:0] data_in_4;
wire      [7:0] data_in_5;
wire      [7:0] data_in_6;
wire      [7:0] data_in_7;
wire      [7:0] data_in_8;
wire      [7:0] data_in_9;
wire            done_ready;
wire            n1;
wire            n10;
wire     [19:0] n1000;
wire      [3:0] n1001;
wire     [19:0] n1002;
wire      [3:0] n1003;
wire     [19:0] n1004;
wire      [3:0] n1005;
wire     [19:0] n1006;
wire      [3:0] n1007;
wire     [19:0] n1008;
wire      [3:0] n1009;
wire            n101;
wire     [19:0] n1010;
wire      [3:0] n1011;
wire     [19:0] n1012;
wire      [3:0] n1013;
wire     [19:0] n1014;
wire      [3:0] n1015;
wire     [19:0] n1016;
wire      [3:0] n1017;
wire     [19:0] n1018;
wire      [3:0] n1019;
wire     [19:0] n1020;
wire      [3:0] n1021;
wire     [19:0] n1022;
wire      [3:0] n1023;
wire     [19:0] n1024;
wire      [3:0] n1025;
wire     [19:0] n1026;
wire      [3:0] n1027;
wire     [19:0] n1028;
wire     [19:0] n1029;
wire            n103;
wire     [31:0] n1030;
wire     [31:0] n1031;
wire     [31:0] n1032;
wire     [31:0] n1033;
wire     [31:0] n1034;
wire      [7:0] n1037;
wire     [19:0] n1038;
wire     [19:0] n1040;
wire      [1:0] n1041;
wire            n1042;
wire      [3:0] n1043;
wire     [19:0] n1046;
wire            n1047;
wire            n105;
wire     [19:0] n1050;
wire            n1051;
wire     [19:0] n1054;
wire            n1055;
wire     [19:0] n1058;
wire     [19:0] n1059;
wire     [19:0] n1060;
wire     [19:0] n1061;
wire     [19:0] n1062;
wire            n1063;
wire      [3:0] n1064;
wire     [19:0] n1067;
wire            n1068;
wire            n107;
wire     [19:0] n1071;
wire            n1072;
wire     [19:0] n1075;
wire            n1076;
wire     [19:0] n1079;
wire     [19:0] n1080;
wire     [19:0] n1081;
wire     [19:0] n1082;
wire     [19:0] n1083;
wire            n1084;
wire     [19:0] n1087;
wire            n1088;
wire            n109;
wire     [19:0] n1091;
wire            n1092;
wire     [19:0] n1095;
wire            n1096;
wire     [19:0] n1099;
wire            n11;
wire     [19:0] n1100;
wire     [19:0] n1101;
wire     [19:0] n1102;
wire     [19:0] n1103;
wire     [19:0] n1104;
wire     [19:0] n1106;
wire            n1107;
wire      [3:0] n1108;
wire            n111;
wire     [19:0] n1111;
wire            n1112;
wire     [19:0] n1115;
wire            n1116;
wire     [19:0] n1119;
wire      [7:0] n112;
wire            n1120;
wire     [19:0] n1123;
wire     [19:0] n1124;
wire     [19:0] n1125;
wire     [19:0] n1126;
wire     [19:0] n1127;
wire            n1128;
wire      [7:0] n113;
wire     [19:0] n1131;
wire            n1132;
wire     [19:0] n1135;
wire            n1136;
wire     [19:0] n1139;
wire      [7:0] n114;
wire            n1140;
wire     [19:0] n1143;
wire     [19:0] n1144;
wire     [19:0] n1145;
wire     [19:0] n1146;
wire     [19:0] n1147;
wire     [19:0] n1148;
wire      [7:0] n115;
wire     [19:0] n1150;
wire            n1151;
wire      [3:0] n1152;
wire     [19:0] n1155;
wire            n1156;
wire     [19:0] n1159;
wire      [7:0] n116;
wire            n1160;
wire     [19:0] n1163;
wire            n1164;
wire     [19:0] n1167;
wire     [19:0] n1168;
wire     [19:0] n1169;
wire      [7:0] n117;
wire     [19:0] n1170;
wire     [19:0] n1171;
wire     [19:0] n1172;
wire     [19:0] n1174;
wire            n1175;
wire      [3:0] n1176;
wire     [19:0] n1179;
wire      [7:0] n118;
wire            n1180;
wire     [19:0] n1183;
wire            n1184;
wire     [19:0] n1187;
wire            n1188;
wire      [7:0] n119;
wire     [19:0] n1191;
wire     [19:0] n1192;
wire     [19:0] n1193;
wire     [19:0] n1194;
wire     [19:0] n1195;
wire     [19:0] n1196;
wire     [19:0] n1198;
wire            n1199;
wire            n12;
wire      [7:0] n120;
wire      [3:0] n1200;
wire     [19:0] n1203;
wire            n1204;
wire     [19:0] n1207;
wire            n1208;
wire      [7:0] n121;
wire     [19:0] n1211;
wire            n1212;
wire     [19:0] n1215;
wire     [19:0] n1216;
wire     [19:0] n1217;
wire     [19:0] n1218;
wire     [19:0] n1219;
wire      [7:0] n122;
wire     [19:0] n1220;
wire     [19:0] n1222;
wire            n1223;
wire      [3:0] n1224;
wire     [19:0] n1227;
wire            n1228;
wire      [7:0] n123;
wire     [19:0] n1231;
wire            n1232;
wire     [19:0] n1235;
wire            n1236;
wire     [19:0] n1239;
wire      [7:0] n124;
wire     [19:0] n1240;
wire     [19:0] n1241;
wire     [19:0] n1242;
wire     [19:0] n1243;
wire     [19:0] n1244;
wire     [19:0] n1246;
wire     [19:0] n1247;
wire     [31:0] n1248;
wire      [7:0] n125;
wire      [7:0] n1251;
wire     [19:0] n1252;
wire     [19:0] n1254;
wire            n1255;
wire      [3:0] n1256;
wire     [19:0] n1259;
wire      [7:0] n126;
wire            n1260;
wire     [19:0] n1263;
wire            n1264;
wire     [19:0] n1267;
wire            n1268;
wire      [7:0] n127;
wire     [19:0] n1271;
wire     [19:0] n1272;
wire     [19:0] n1273;
wire     [19:0] n1274;
wire     [19:0] n1275;
wire            n1276;
wire      [3:0] n1277;
wire      [7:0] n128;
wire     [19:0] n1280;
wire            n1281;
wire     [19:0] n1284;
wire            n1285;
wire     [19:0] n1288;
wire            n1289;
wire      [7:0] n129;
wire     [19:0] n1292;
wire     [19:0] n1293;
wire     [19:0] n1294;
wire     [19:0] n1295;
wire     [19:0] n1296;
wire            n1297;
wire            n13;
wire      [7:0] n130;
wire     [19:0] n1300;
wire            n1301;
wire     [19:0] n1304;
wire            n1305;
wire     [19:0] n1308;
wire            n1309;
wire      [7:0] n131;
wire     [19:0] n1312;
wire     [19:0] n1313;
wire     [19:0] n1314;
wire     [19:0] n1315;
wire     [19:0] n1316;
wire     [19:0] n1317;
wire     [19:0] n1319;
wire      [7:0] n132;
wire            n1320;
wire      [3:0] n1321;
wire     [19:0] n1324;
wire            n1325;
wire     [19:0] n1328;
wire            n1329;
wire      [7:0] n133;
wire     [19:0] n1332;
wire            n1333;
wire     [19:0] n1336;
wire     [19:0] n1337;
wire     [19:0] n1338;
wire     [19:0] n1339;
wire      [7:0] n134;
wire     [19:0] n1340;
wire            n1341;
wire     [19:0] n1344;
wire            n1345;
wire     [19:0] n1348;
wire            n1349;
wire      [7:0] n135;
wire     [19:0] n1352;
wire            n1353;
wire     [19:0] n1356;
wire     [19:0] n1357;
wire     [19:0] n1358;
wire     [19:0] n1359;
wire      [7:0] n136;
wire     [19:0] n1360;
wire     [19:0] n1361;
wire     [19:0] n1363;
wire            n1364;
wire      [3:0] n1365;
wire     [19:0] n1368;
wire            n1369;
wire      [7:0] n137;
wire     [19:0] n1372;
wire            n1373;
wire     [19:0] n1376;
wire            n1377;
wire      [7:0] n138;
wire     [19:0] n1380;
wire     [19:0] n1381;
wire     [19:0] n1382;
wire     [19:0] n1383;
wire     [19:0] n1384;
wire     [19:0] n1385;
wire     [19:0] n1387;
wire            n1388;
wire      [3:0] n1389;
wire      [7:0] n139;
wire     [19:0] n1392;
wire            n1393;
wire     [19:0] n1396;
wire            n1397;
wire            n14;
wire      [7:0] n140;
wire     [19:0] n1400;
wire            n1401;
wire     [19:0] n1404;
wire     [19:0] n1405;
wire     [19:0] n1406;
wire     [19:0] n1407;
wire     [19:0] n1408;
wire     [19:0] n1409;
wire      [7:0] n141;
wire     [19:0] n1411;
wire            n1412;
wire      [3:0] n1413;
wire     [19:0] n1416;
wire            n1417;
wire      [7:0] n142;
wire     [19:0] n1420;
wire            n1421;
wire     [19:0] n1424;
wire            n1425;
wire     [19:0] n1428;
wire     [19:0] n1429;
wire      [7:0] n143;
wire     [19:0] n1430;
wire     [19:0] n1431;
wire     [19:0] n1432;
wire     [19:0] n1433;
wire     [19:0] n1435;
wire            n1436;
wire      [3:0] n1437;
wire      [3:0] n144;
wire     [19:0] n1440;
wire            n1441;
wire     [19:0] n1444;
wire            n1445;
wire     [19:0] n1448;
wire            n1449;
wire     [19:0] n1452;
wire     [19:0] n1453;
wire     [19:0] n1454;
wire     [19:0] n1455;
wire     [19:0] n1456;
wire     [19:0] n1457;
wire     [19:0] n1459;
wire            n146;
wire     [19:0] n1460;
wire     [31:0] n1461;
wire      [7:0] n1464;
wire     [19:0] n1465;
wire     [19:0] n1467;
wire            n1468;
wire      [3:0] n1469;
wire            n147;
wire     [19:0] n1472;
wire            n1473;
wire     [19:0] n1476;
wire            n1477;
wire            n148;
wire     [19:0] n1480;
wire            n1481;
wire     [19:0] n1484;
wire     [19:0] n1485;
wire     [19:0] n1486;
wire     [19:0] n1487;
wire     [19:0] n1488;
wire            n1489;
wire            n149;
wire      [3:0] n1490;
wire     [19:0] n1493;
wire            n1494;
wire     [19:0] n1497;
wire            n1498;
wire            n150;
wire     [19:0] n1501;
wire            n1502;
wire     [19:0] n1505;
wire     [19:0] n1506;
wire     [19:0] n1507;
wire     [19:0] n1508;
wire     [19:0] n1509;
wire            n151;
wire            n1510;
wire     [19:0] n1513;
wire            n1514;
wire     [19:0] n1517;
wire            n1518;
wire            n152;
wire     [19:0] n1521;
wire            n1522;
wire     [19:0] n1525;
wire     [19:0] n1526;
wire     [19:0] n1527;
wire     [19:0] n1528;
wire     [19:0] n1529;
wire            n153;
wire     [19:0] n1530;
wire     [19:0] n1532;
wire            n1533;
wire      [3:0] n1534;
wire     [19:0] n1537;
wire            n1538;
wire            n154;
wire     [19:0] n1541;
wire            n1542;
wire     [19:0] n1545;
wire            n1546;
wire     [19:0] n1549;
wire            n155;
wire     [19:0] n1550;
wire     [19:0] n1551;
wire     [19:0] n1552;
wire     [19:0] n1553;
wire            n1554;
wire     [19:0] n1557;
wire            n1558;
wire            n156;
wire     [19:0] n1561;
wire            n1562;
wire     [19:0] n1565;
wire            n1566;
wire     [19:0] n1569;
wire            n157;
wire     [19:0] n1570;
wire     [19:0] n1571;
wire     [19:0] n1572;
wire     [19:0] n1573;
wire     [19:0] n1574;
wire     [19:0] n1576;
wire            n1577;
wire      [3:0] n1578;
wire            n158;
wire     [19:0] n1581;
wire            n1582;
wire     [19:0] n1585;
wire            n1586;
wire     [19:0] n1589;
wire            n159;
wire            n1590;
wire     [19:0] n1593;
wire     [19:0] n1594;
wire     [19:0] n1595;
wire     [19:0] n1596;
wire     [19:0] n1597;
wire     [19:0] n1598;
wire            n16;
wire     [19:0] n1600;
wire            n1601;
wire      [3:0] n1602;
wire     [19:0] n1605;
wire            n1606;
wire     [19:0] n1609;
wire            n161;
wire            n1610;
wire     [19:0] n1613;
wire            n1614;
wire     [19:0] n1617;
wire     [19:0] n1618;
wire     [19:0] n1619;
wire            n162;
wire     [19:0] n1620;
wire     [19:0] n1621;
wire     [19:0] n1622;
wire     [19:0] n1624;
wire            n1625;
wire      [3:0] n1626;
wire     [19:0] n1629;
wire            n163;
wire            n1630;
wire     [19:0] n1633;
wire            n1634;
wire     [19:0] n1637;
wire            n1638;
wire            n164;
wire     [19:0] n1641;
wire     [19:0] n1642;
wire     [19:0] n1643;
wire     [19:0] n1644;
wire     [19:0] n1645;
wire     [19:0] n1646;
wire     [19:0] n1648;
wire            n1649;
wire            n165;
wire      [3:0] n1650;
wire     [19:0] n1653;
wire            n1654;
wire     [19:0] n1657;
wire            n1658;
wire     [19:0] n1661;
wire            n1662;
wire     [19:0] n1665;
wire     [19:0] n1666;
wire     [19:0] n1667;
wire     [19:0] n1668;
wire     [19:0] n1669;
wire            n167;
wire     [19:0] n1670;
wire     [19:0] n1672;
wire     [19:0] n1673;
wire     [31:0] n1674;
wire      [7:0] n1677;
wire     [19:0] n1678;
wire            n168;
wire     [19:0] n1680;
wire            n1681;
wire      [3:0] n1682;
wire     [19:0] n1685;
wire            n1686;
wire     [19:0] n1689;
wire            n169;
wire            n1690;
wire     [19:0] n1693;
wire            n1694;
wire     [19:0] n1697;
wire     [19:0] n1698;
wire     [19:0] n1699;
wire            n17;
wire            n170;
wire     [19:0] n1700;
wire     [19:0] n1701;
wire            n1702;
wire      [3:0] n1703;
wire     [19:0] n1706;
wire            n1707;
wire            n171;
wire     [19:0] n1710;
wire            n1711;
wire     [19:0] n1714;
wire            n1715;
wire     [19:0] n1718;
wire     [19:0] n1719;
wire            n172;
wire     [19:0] n1720;
wire     [19:0] n1721;
wire     [19:0] n1722;
wire            n1723;
wire     [19:0] n1726;
wire            n1727;
wire            n173;
wire     [19:0] n1730;
wire            n1731;
wire     [19:0] n1734;
wire            n1735;
wire     [19:0] n1738;
wire     [19:0] n1739;
wire            n174;
wire     [19:0] n1740;
wire     [19:0] n1741;
wire     [19:0] n1742;
wire     [19:0] n1743;
wire     [19:0] n1745;
wire            n1746;
wire      [3:0] n1747;
wire            n175;
wire     [19:0] n1750;
wire            n1751;
wire     [19:0] n1754;
wire            n1755;
wire     [19:0] n1758;
wire            n1759;
wire     [19:0] n1762;
wire     [19:0] n1763;
wire     [19:0] n1764;
wire     [19:0] n1765;
wire     [19:0] n1766;
wire            n1767;
wire            n177;
wire     [19:0] n1770;
wire            n1771;
wire     [19:0] n1774;
wire            n1775;
wire     [19:0] n1778;
wire            n1779;
wire            n178;
wire     [19:0] n1782;
wire     [19:0] n1783;
wire     [19:0] n1784;
wire     [19:0] n1785;
wire     [19:0] n1786;
wire     [19:0] n1787;
wire     [19:0] n1789;
wire            n179;
wire            n1790;
wire      [3:0] n1791;
wire     [19:0] n1794;
wire            n1795;
wire     [19:0] n1798;
wire            n1799;
wire            n18;
wire            n180;
wire     [19:0] n1802;
wire            n1803;
wire     [19:0] n1806;
wire     [19:0] n1807;
wire     [19:0] n1808;
wire     [19:0] n1809;
wire            n181;
wire     [19:0] n1810;
wire     [19:0] n1811;
wire     [19:0] n1813;
wire            n1814;
wire      [3:0] n1815;
wire     [19:0] n1818;
wire            n1819;
wire            n182;
wire     [19:0] n1822;
wire            n1823;
wire     [19:0] n1826;
wire            n1827;
wire            n183;
wire     [19:0] n1830;
wire     [19:0] n1831;
wire     [19:0] n1832;
wire     [19:0] n1833;
wire     [19:0] n1834;
wire     [19:0] n1835;
wire     [19:0] n1837;
wire            n1838;
wire      [3:0] n1839;
wire     [19:0] n1842;
wire            n1843;
wire     [19:0] n1846;
wire            n1847;
wire            n185;
wire     [19:0] n1850;
wire            n1851;
wire     [19:0] n1854;
wire     [19:0] n1855;
wire     [19:0] n1856;
wire     [19:0] n1857;
wire     [19:0] n1858;
wire     [19:0] n1859;
wire            n186;
wire     [19:0] n1861;
wire            n1862;
wire      [3:0] n1863;
wire     [19:0] n1866;
wire            n1867;
wire            n187;
wire     [19:0] n1870;
wire            n1871;
wire     [19:0] n1874;
wire            n1875;
wire     [19:0] n1878;
wire     [19:0] n1879;
wire            n188;
wire     [19:0] n1880;
wire     [19:0] n1881;
wire     [19:0] n1882;
wire     [19:0] n1883;
wire     [19:0] n1885;
wire     [19:0] n1886;
wire     [31:0] n1887;
wire            n189;
wire      [7:0] n1890;
wire     [19:0] n1891;
wire     [19:0] n1893;
wire            n1894;
wire      [3:0] n1895;
wire     [19:0] n1898;
wire            n1899;
wire            n19;
wire     [19:0] n1902;
wire            n1903;
wire     [19:0] n1906;
wire            n1907;
wire            n191;
wire     [19:0] n1910;
wire     [19:0] n1911;
wire     [19:0] n1912;
wire     [19:0] n1913;
wire     [19:0] n1914;
wire            n1915;
wire      [3:0] n1916;
wire     [19:0] n1919;
wire            n192;
wire            n1920;
wire     [19:0] n1923;
wire            n1924;
wire     [19:0] n1927;
wire            n1928;
wire            n193;
wire     [19:0] n1931;
wire     [19:0] n1932;
wire     [19:0] n1933;
wire     [19:0] n1934;
wire     [19:0] n1935;
wire            n1936;
wire     [19:0] n1939;
wire            n194;
wire            n1940;
wire     [19:0] n1943;
wire            n1944;
wire     [19:0] n1947;
wire            n1948;
wire            n195;
wire     [19:0] n1951;
wire     [19:0] n1952;
wire     [19:0] n1953;
wire     [19:0] n1954;
wire     [19:0] n1955;
wire     [19:0] n1956;
wire     [19:0] n1958;
wire            n1959;
wire      [3:0] n1960;
wire     [19:0] n1963;
wire            n1964;
wire     [19:0] n1967;
wire            n1968;
wire            n197;
wire     [19:0] n1971;
wire            n1972;
wire     [19:0] n1975;
wire     [19:0] n1976;
wire     [19:0] n1977;
wire     [19:0] n1978;
wire     [19:0] n1979;
wire            n198;
wire            n1980;
wire     [19:0] n1983;
wire            n1984;
wire     [19:0] n1987;
wire            n1988;
wire            n199;
wire     [19:0] n1991;
wire            n1992;
wire     [19:0] n1995;
wire     [19:0] n1996;
wire     [19:0] n1997;
wire     [19:0] n1998;
wire     [19:0] n1999;
wire            n20;
wire            n200;
wire     [19:0] n2000;
wire     [19:0] n2002;
wire            n2003;
wire      [3:0] n2004;
wire     [19:0] n2007;
wire            n2008;
wire            n201;
wire     [19:0] n2011;
wire            n2012;
wire     [19:0] n2015;
wire            n2016;
wire     [19:0] n2019;
wire     [19:0] n2020;
wire     [19:0] n2021;
wire     [19:0] n2022;
wire     [19:0] n2023;
wire     [19:0] n2024;
wire     [19:0] n2026;
wire            n2027;
wire      [3:0] n2028;
wire            n203;
wire     [19:0] n2031;
wire            n2032;
wire     [19:0] n2035;
wire            n2036;
wire     [19:0] n2039;
wire            n204;
wire            n2040;
wire     [19:0] n2043;
wire     [19:0] n2044;
wire     [19:0] n2045;
wire     [19:0] n2046;
wire     [19:0] n2047;
wire     [19:0] n2048;
wire            n205;
wire     [19:0] n2050;
wire            n2051;
wire      [3:0] n2052;
wire     [19:0] n2055;
wire            n2056;
wire     [19:0] n2059;
wire            n206;
wire            n2060;
wire     [19:0] n2063;
wire            n2064;
wire     [19:0] n2067;
wire     [19:0] n2068;
wire     [19:0] n2069;
wire            n207;
wire     [19:0] n2070;
wire     [19:0] n2071;
wire     [19:0] n2072;
wire     [19:0] n2074;
wire            n2075;
wire      [3:0] n2076;
wire     [19:0] n2079;
wire            n2080;
wire     [19:0] n2083;
wire            n2084;
wire     [19:0] n2087;
wire            n2088;
wire            n209;
wire     [19:0] n2091;
wire     [19:0] n2092;
wire     [19:0] n2093;
wire     [19:0] n2094;
wire     [19:0] n2095;
wire     [19:0] n2096;
wire     [19:0] n2098;
wire     [19:0] n2099;
wire            n210;
wire     [31:0] n2100;
wire      [7:0] n2103;
wire     [19:0] n2104;
wire     [19:0] n2106;
wire            n2107;
wire      [3:0] n2108;
wire            n211;
wire     [19:0] n2111;
wire            n2112;
wire     [19:0] n2115;
wire            n2116;
wire     [19:0] n2119;
wire            n212;
wire            n2120;
wire     [19:0] n2123;
wire     [19:0] n2124;
wire     [19:0] n2125;
wire     [19:0] n2126;
wire     [19:0] n2127;
wire            n2128;
wire      [3:0] n2129;
wire            n213;
wire     [19:0] n2132;
wire            n2133;
wire     [19:0] n2136;
wire            n2137;
wire     [19:0] n2140;
wire            n2141;
wire     [19:0] n2144;
wire     [19:0] n2145;
wire     [19:0] n2146;
wire     [19:0] n2147;
wire     [19:0] n2148;
wire            n2149;
wire            n215;
wire     [19:0] n2152;
wire            n2153;
wire     [19:0] n2156;
wire            n2157;
wire            n216;
wire     [19:0] n2160;
wire            n2161;
wire     [19:0] n2164;
wire     [19:0] n2165;
wire     [19:0] n2166;
wire     [19:0] n2167;
wire     [19:0] n2168;
wire     [19:0] n2169;
wire            n217;
wire     [19:0] n2171;
wire            n2172;
wire      [3:0] n2173;
wire     [19:0] n2176;
wire            n2177;
wire            n218;
wire     [19:0] n2180;
wire            n2181;
wire     [19:0] n2184;
wire            n2185;
wire     [19:0] n2188;
wire     [19:0] n2189;
wire            n219;
wire     [19:0] n2190;
wire     [19:0] n2191;
wire     [19:0] n2192;
wire            n2193;
wire     [19:0] n2196;
wire            n2197;
wire            n22;
wire     [19:0] n2200;
wire            n2201;
wire     [19:0] n2204;
wire            n2205;
wire     [19:0] n2208;
wire     [19:0] n2209;
wire            n221;
wire     [19:0] n2210;
wire     [19:0] n2211;
wire     [19:0] n2212;
wire     [19:0] n2213;
wire     [19:0] n2215;
wire            n2216;
wire      [3:0] n2217;
wire            n222;
wire     [19:0] n2220;
wire            n2221;
wire     [19:0] n2224;
wire            n2225;
wire     [19:0] n2228;
wire            n2229;
wire            n223;
wire     [19:0] n2232;
wire     [19:0] n2233;
wire     [19:0] n2234;
wire     [19:0] n2235;
wire     [19:0] n2236;
wire     [19:0] n2237;
wire     [19:0] n2239;
wire            n2240;
wire      [3:0] n2241;
wire     [19:0] n2244;
wire            n2245;
wire     [19:0] n2248;
wire            n2249;
wire            n225;
wire     [19:0] n2252;
wire            n2253;
wire     [19:0] n2256;
wire     [19:0] n2257;
wire     [19:0] n2258;
wire     [19:0] n2259;
wire            n226;
wire     [19:0] n2260;
wire     [19:0] n2261;
wire     [19:0] n2263;
wire            n2264;
wire      [3:0] n2265;
wire     [19:0] n2268;
wire            n2269;
wire            n227;
wire     [19:0] n2272;
wire            n2273;
wire     [19:0] n2276;
wire            n2277;
wire            n228;
wire     [19:0] n2280;
wire     [19:0] n2281;
wire     [19:0] n2282;
wire     [19:0] n2283;
wire     [19:0] n2284;
wire     [19:0] n2285;
wire     [19:0] n2287;
wire            n2288;
wire      [3:0] n2289;
wire            n229;
wire     [19:0] n2292;
wire            n2293;
wire     [19:0] n2296;
wire            n2297;
wire            n23;
wire            n230;
wire     [19:0] n2300;
wire            n2301;
wire     [19:0] n2304;
wire     [19:0] n2305;
wire     [19:0] n2306;
wire     [19:0] n2307;
wire     [19:0] n2308;
wire     [19:0] n2309;
wire            n231;
wire     [19:0] n2311;
wire     [19:0] n2312;
wire     [31:0] n2313;
wire      [7:0] n2316;
wire     [19:0] n2317;
wire     [19:0] n2319;
wire            n232;
wire            n2320;
wire      [3:0] n2321;
wire     [19:0] n2324;
wire            n2325;
wire     [19:0] n2328;
wire            n2329;
wire            n233;
wire     [19:0] n2332;
wire            n2333;
wire     [19:0] n2336;
wire     [19:0] n2337;
wire     [19:0] n2338;
wire     [19:0] n2339;
wire            n234;
wire     [19:0] n2340;
wire            n2341;
wire      [3:0] n2342;
wire     [19:0] n2345;
wire            n2346;
wire     [19:0] n2349;
wire            n235;
wire            n2350;
wire     [19:0] n2353;
wire            n2354;
wire     [19:0] n2357;
wire     [19:0] n2358;
wire     [19:0] n2359;
wire            n236;
wire     [19:0] n2360;
wire     [19:0] n2361;
wire            n2362;
wire     [19:0] n2365;
wire            n2366;
wire     [19:0] n2369;
wire            n237;
wire            n2370;
wire     [19:0] n2373;
wire            n2374;
wire     [19:0] n2377;
wire     [19:0] n2378;
wire     [19:0] n2379;
wire            n238;
wire     [19:0] n2380;
wire     [19:0] n2381;
wire     [19:0] n2382;
wire     [19:0] n2384;
wire            n2385;
wire      [3:0] n2386;
wire     [19:0] n2389;
wire            n239;
wire            n2390;
wire     [19:0] n2393;
wire            n2394;
wire     [19:0] n2397;
wire            n2398;
wire            n24;
wire            n240;
wire     [19:0] n2401;
wire     [19:0] n2402;
wire     [19:0] n2403;
wire     [19:0] n2404;
wire     [19:0] n2405;
wire            n2406;
wire     [19:0] n2409;
wire            n241;
wire            n2410;
wire     [19:0] n2413;
wire            n2414;
wire     [19:0] n2417;
wire            n2418;
wire            n242;
wire     [19:0] n2421;
wire     [19:0] n2422;
wire     [19:0] n2423;
wire     [19:0] n2424;
wire     [19:0] n2425;
wire     [19:0] n2426;
wire     [19:0] n2428;
wire            n2429;
wire            n243;
wire      [3:0] n2430;
wire     [19:0] n2433;
wire            n2434;
wire     [19:0] n2437;
wire            n2438;
wire            n244;
wire     [19:0] n2441;
wire            n2442;
wire     [19:0] n2445;
wire     [19:0] n2446;
wire     [19:0] n2447;
wire     [19:0] n2448;
wire     [19:0] n2449;
wire      [7:0] n245;
wire     [19:0] n2450;
wire     [19:0] n2452;
wire            n2453;
wire      [3:0] n2454;
wire     [19:0] n2457;
wire            n2458;
wire      [5:0] n246;
wire     [19:0] n2461;
wire            n2462;
wire     [19:0] n2465;
wire            n2466;
wire     [19:0] n2469;
wire            n247;
wire     [19:0] n2470;
wire     [19:0] n2471;
wire     [19:0] n2472;
wire     [19:0] n2473;
wire     [19:0] n2474;
wire     [19:0] n2476;
wire            n2477;
wire      [3:0] n2478;
wire     [19:0] n2481;
wire            n2482;
wire     [19:0] n2485;
wire            n2486;
wire     [19:0] n2489;
wire      [7:0] n249;
wire            n2490;
wire     [19:0] n2493;
wire     [19:0] n2494;
wire     [19:0] n2495;
wire     [19:0] n2496;
wire     [19:0] n2497;
wire     [19:0] n2498;
wire            n250;
wire     [19:0] n2500;
wire            n2501;
wire      [3:0] n2502;
wire     [19:0] n2505;
wire            n2506;
wire     [19:0] n2509;
wire            n251;
wire            n2510;
wire     [19:0] n2513;
wire            n2514;
wire     [19:0] n2517;
wire     [19:0] n2518;
wire     [19:0] n2519;
wire            n252;
wire     [19:0] n2520;
wire     [19:0] n2521;
wire     [19:0] n2522;
wire     [19:0] n2524;
wire     [19:0] n2525;
wire     [31:0] n2526;
wire      [7:0] n2529;
wire      [5:0] n253;
wire     [19:0] n2530;
wire     [19:0] n2532;
wire            n2533;
wire      [3:0] n2534;
wire     [19:0] n2537;
wire            n2538;
wire            n254;
wire     [19:0] n2541;
wire            n2542;
wire     [19:0] n2545;
wire            n2546;
wire     [19:0] n2549;
wire      [7:0] n255;
wire     [19:0] n2550;
wire     [19:0] n2551;
wire     [19:0] n2552;
wire     [19:0] n2553;
wire            n2554;
wire      [3:0] n2555;
wire     [19:0] n2558;
wire            n2559;
wire            n256;
wire     [19:0] n2562;
wire            n2563;
wire     [19:0] n2566;
wire            n2567;
wire            n257;
wire     [19:0] n2570;
wire     [19:0] n2571;
wire     [19:0] n2572;
wire     [19:0] n2573;
wire     [19:0] n2574;
wire            n2575;
wire     [19:0] n2578;
wire            n2579;
wire            n258;
wire     [19:0] n2582;
wire            n2583;
wire     [19:0] n2586;
wire            n2587;
wire      [5:0] n259;
wire     [19:0] n2590;
wire     [19:0] n2591;
wire     [19:0] n2592;
wire     [19:0] n2593;
wire     [19:0] n2594;
wire     [19:0] n2595;
wire     [19:0] n2597;
wire            n2598;
wire      [3:0] n2599;
wire            n26;
wire            n260;
wire     [19:0] n2602;
wire            n2603;
wire     [19:0] n2606;
wire            n2607;
wire      [7:0] n261;
wire     [19:0] n2610;
wire            n2611;
wire     [19:0] n2614;
wire     [19:0] n2615;
wire     [19:0] n2616;
wire     [19:0] n2617;
wire     [19:0] n2618;
wire            n2619;
wire            n262;
wire     [19:0] n2622;
wire            n2623;
wire     [19:0] n2626;
wire            n2627;
wire            n263;
wire     [19:0] n2630;
wire            n2631;
wire     [19:0] n2634;
wire     [19:0] n2635;
wire     [19:0] n2636;
wire     [19:0] n2637;
wire     [19:0] n2638;
wire     [19:0] n2639;
wire            n264;
wire     [19:0] n2641;
wire            n2642;
wire      [3:0] n2643;
wire     [19:0] n2646;
wire            n2647;
wire      [5:0] n265;
wire     [19:0] n2650;
wire            n2651;
wire     [19:0] n2654;
wire            n2655;
wire     [19:0] n2658;
wire     [19:0] n2659;
wire            n266;
wire     [19:0] n2660;
wire     [19:0] n2661;
wire     [19:0] n2662;
wire     [19:0] n2663;
wire     [19:0] n2665;
wire            n2666;
wire      [3:0] n2667;
wire      [7:0] n267;
wire     [19:0] n2670;
wire            n2671;
wire     [19:0] n2674;
wire            n2675;
wire     [19:0] n2678;
wire            n2679;
wire            n268;
wire     [19:0] n2682;
wire     [19:0] n2683;
wire     [19:0] n2684;
wire     [19:0] n2685;
wire     [19:0] n2686;
wire     [19:0] n2687;
wire     [19:0] n2689;
wire            n269;
wire            n2690;
wire      [3:0] n2691;
wire     [19:0] n2694;
wire            n2695;
wire     [19:0] n2698;
wire            n2699;
wire            n27;
wire            n270;
wire     [19:0] n2702;
wire            n2703;
wire     [19:0] n2706;
wire     [19:0] n2707;
wire     [19:0] n2708;
wire     [19:0] n2709;
wire      [5:0] n271;
wire     [19:0] n2710;
wire     [19:0] n2711;
wire     [19:0] n2713;
wire            n2714;
wire      [3:0] n2715;
wire     [19:0] n2718;
wire            n2719;
wire            n272;
wire     [19:0] n2722;
wire            n2723;
wire     [19:0] n2726;
wire            n2727;
wire      [7:0] n273;
wire     [19:0] n2730;
wire     [19:0] n2731;
wire     [19:0] n2732;
wire     [19:0] n2733;
wire     [19:0] n2734;
wire     [19:0] n2735;
wire     [19:0] n2737;
wire     [19:0] n2738;
wire     [31:0] n2739;
wire            n274;
wire      [7:0] n2742;
wire     [19:0] n2743;
wire     [19:0] n2745;
wire            n2746;
wire      [3:0] n2747;
wire            n275;
wire     [19:0] n2750;
wire            n2751;
wire     [19:0] n2754;
wire            n2755;
wire     [19:0] n2758;
wire            n2759;
wire            n276;
wire     [19:0] n2762;
wire     [19:0] n2763;
wire     [19:0] n2764;
wire     [19:0] n2765;
wire     [19:0] n2766;
wire            n2767;
wire      [3:0] n2768;
wire      [5:0] n277;
wire     [19:0] n2771;
wire            n2772;
wire     [19:0] n2775;
wire            n2776;
wire     [19:0] n2779;
wire            n278;
wire            n2780;
wire     [19:0] n2783;
wire     [19:0] n2784;
wire     [19:0] n2785;
wire     [19:0] n2786;
wire     [19:0] n2787;
wire            n2788;
wire      [7:0] n279;
wire     [19:0] n2791;
wire            n2792;
wire     [19:0] n2795;
wire            n2796;
wire     [19:0] n2799;
wire            n28;
wire            n280;
wire            n2800;
wire     [19:0] n2803;
wire     [19:0] n2804;
wire     [19:0] n2805;
wire     [19:0] n2806;
wire     [19:0] n2807;
wire     [19:0] n2808;
wire            n281;
wire     [19:0] n2810;
wire            n2811;
wire      [3:0] n2812;
wire     [19:0] n2815;
wire            n2816;
wire     [19:0] n2819;
wire            n282;
wire            n2820;
wire     [19:0] n2823;
wire            n2824;
wire     [19:0] n2827;
wire     [19:0] n2828;
wire     [19:0] n2829;
wire      [5:0] n283;
wire     [19:0] n2830;
wire     [19:0] n2831;
wire            n2832;
wire     [19:0] n2835;
wire            n2836;
wire     [19:0] n2839;
wire            n284;
wire            n2840;
wire     [19:0] n2843;
wire            n2844;
wire     [19:0] n2847;
wire     [19:0] n2848;
wire     [19:0] n2849;
wire      [7:0] n285;
wire     [19:0] n2850;
wire     [19:0] n2851;
wire     [19:0] n2852;
wire     [19:0] n2854;
wire            n2855;
wire      [3:0] n2856;
wire     [19:0] n2859;
wire            n286;
wire            n2860;
wire     [19:0] n2863;
wire            n2864;
wire     [19:0] n2867;
wire            n2868;
wire            n287;
wire     [19:0] n2871;
wire     [19:0] n2872;
wire     [19:0] n2873;
wire     [19:0] n2874;
wire     [19:0] n2875;
wire     [19:0] n2876;
wire     [19:0] n2878;
wire            n2879;
wire            n288;
wire      [3:0] n2880;
wire     [19:0] n2883;
wire            n2884;
wire     [19:0] n2887;
wire            n2888;
wire      [5:0] n289;
wire     [19:0] n2891;
wire            n2892;
wire     [19:0] n2895;
wire     [19:0] n2896;
wire     [19:0] n2897;
wire     [19:0] n2898;
wire     [19:0] n2899;
wire            n29;
wire            n290;
wire     [19:0] n2900;
wire     [19:0] n2902;
wire            n2903;
wire      [3:0] n2904;
wire     [19:0] n2907;
wire            n2908;
wire      [7:0] n291;
wire     [19:0] n2911;
wire            n2912;
wire     [19:0] n2915;
wire            n2916;
wire     [19:0] n2919;
wire            n292;
wire     [19:0] n2920;
wire     [19:0] n2921;
wire     [19:0] n2922;
wire     [19:0] n2923;
wire     [19:0] n2924;
wire     [19:0] n2926;
wire            n2927;
wire      [3:0] n2928;
wire            n293;
wire     [19:0] n2931;
wire            n2932;
wire     [19:0] n2935;
wire            n2936;
wire     [19:0] n2939;
wire            n294;
wire            n2940;
wire     [19:0] n2943;
wire     [19:0] n2944;
wire     [19:0] n2945;
wire     [19:0] n2946;
wire     [19:0] n2947;
wire     [19:0] n2948;
wire      [5:0] n295;
wire     [19:0] n2950;
wire     [19:0] n2951;
wire     [31:0] n2952;
wire      [7:0] n2955;
wire     [19:0] n2956;
wire     [19:0] n2958;
wire            n2959;
wire            n296;
wire      [3:0] n2960;
wire     [19:0] n2963;
wire            n2964;
wire     [19:0] n2967;
wire            n2968;
wire      [7:0] n297;
wire     [19:0] n2971;
wire            n2972;
wire     [19:0] n2975;
wire     [19:0] n2976;
wire     [19:0] n2977;
wire     [19:0] n2978;
wire     [19:0] n2979;
wire            n298;
wire            n2980;
wire      [3:0] n2981;
wire     [19:0] n2984;
wire            n2985;
wire     [19:0] n2988;
wire            n2989;
wire            n299;
wire     [19:0] n2992;
wire            n2993;
wire     [19:0] n2996;
wire     [19:0] n2997;
wire     [19:0] n2998;
wire     [19:0] n2999;
wire            n3;
wire            n30;
wire            n300;
wire     [19:0] n3000;
wire            n3001;
wire     [19:0] n3004;
wire            n3005;
wire     [19:0] n3008;
wire            n3009;
wire      [5:0] n301;
wire     [19:0] n3012;
wire            n3013;
wire     [19:0] n3016;
wire     [19:0] n3017;
wire     [19:0] n3018;
wire     [19:0] n3019;
wire            n302;
wire     [19:0] n3020;
wire     [19:0] n3021;
wire     [19:0] n3023;
wire            n3024;
wire      [3:0] n3025;
wire     [19:0] n3028;
wire            n3029;
wire      [7:0] n303;
wire     [19:0] n3032;
wire            n3033;
wire     [19:0] n3036;
wire            n3037;
wire            n304;
wire     [19:0] n3040;
wire     [19:0] n3041;
wire     [19:0] n3042;
wire     [19:0] n3043;
wire     [19:0] n3044;
wire            n3045;
wire     [19:0] n3048;
wire            n3049;
wire            n305;
wire     [19:0] n3052;
wire            n3053;
wire     [19:0] n3056;
wire            n3057;
wire            n306;
wire     [19:0] n3060;
wire     [19:0] n3061;
wire     [19:0] n3062;
wire     [19:0] n3063;
wire     [19:0] n3064;
wire     [19:0] n3065;
wire     [19:0] n3067;
wire            n3068;
wire      [3:0] n3069;
wire      [5:0] n307;
wire     [19:0] n3072;
wire            n3073;
wire     [19:0] n3076;
wire            n3077;
wire            n308;
wire     [19:0] n3080;
wire            n3081;
wire     [19:0] n3084;
wire     [19:0] n3085;
wire     [19:0] n3086;
wire     [19:0] n3087;
wire     [19:0] n3088;
wire     [19:0] n3089;
wire      [7:0] n309;
wire     [19:0] n3091;
wire            n3092;
wire      [3:0] n3093;
wire     [19:0] n3096;
wire            n3097;
wire            n31;
wire            n310;
wire     [19:0] n3100;
wire            n3101;
wire     [19:0] n3104;
wire            n3105;
wire     [19:0] n3108;
wire     [19:0] n3109;
wire            n311;
wire     [19:0] n3110;
wire     [19:0] n3111;
wire     [19:0] n3112;
wire     [19:0] n3113;
wire     [19:0] n3115;
wire            n3116;
wire      [3:0] n3117;
wire            n312;
wire     [19:0] n3120;
wire            n3121;
wire     [19:0] n3124;
wire            n3125;
wire     [19:0] n3128;
wire            n3129;
wire      [5:0] n313;
wire     [19:0] n3132;
wire     [19:0] n3133;
wire     [19:0] n3134;
wire     [19:0] n3135;
wire     [19:0] n3136;
wire     [19:0] n3137;
wire     [19:0] n3139;
wire            n314;
wire            n3140;
wire      [3:0] n3141;
wire     [19:0] n3144;
wire            n3145;
wire     [19:0] n3148;
wire            n3149;
wire      [7:0] n315;
wire     [19:0] n3152;
wire            n3153;
wire     [19:0] n3156;
wire     [19:0] n3157;
wire     [19:0] n3158;
wire     [19:0] n3159;
wire            n316;
wire     [19:0] n3160;
wire     [19:0] n3161;
wire     [19:0] n3163;
wire     [19:0] n3164;
wire     [31:0] n3165;
wire      [7:0] n3168;
wire     [19:0] n3169;
wire            n317;
wire     [19:0] n3171;
wire            n3172;
wire      [3:0] n3173;
wire     [19:0] n3176;
wire            n3177;
wire            n318;
wire     [19:0] n3180;
wire            n3181;
wire     [19:0] n3184;
wire            n3185;
wire     [19:0] n3188;
wire     [19:0] n3189;
wire            n319;
wire     [19:0] n3190;
wire     [19:0] n3191;
wire     [19:0] n3192;
wire            n3193;
wire      [3:0] n3194;
wire     [19:0] n3197;
wire            n3198;
wire            n320;
wire     [19:0] n3201;
wire            n3202;
wire     [19:0] n3205;
wire            n3206;
wire     [19:0] n3209;
wire            n321;
wire     [19:0] n3210;
wire     [19:0] n3211;
wire     [19:0] n3212;
wire     [19:0] n3213;
wire            n3214;
wire     [19:0] n3217;
wire            n3218;
wire            n322;
wire     [19:0] n3221;
wire            n3222;
wire     [19:0] n3225;
wire            n3226;
wire     [19:0] n3229;
wire            n323;
wire     [19:0] n3230;
wire     [19:0] n3231;
wire     [19:0] n3232;
wire     [19:0] n3233;
wire     [19:0] n3234;
wire     [19:0] n3236;
wire            n3237;
wire      [3:0] n3238;
wire            n324;
wire     [19:0] n3241;
wire            n3242;
wire     [19:0] n3245;
wire            n3246;
wire     [19:0] n3249;
wire            n325;
wire            n3250;
wire     [19:0] n3253;
wire     [19:0] n3254;
wire     [19:0] n3255;
wire     [19:0] n3256;
wire     [19:0] n3257;
wire            n3258;
wire            n326;
wire     [19:0] n3261;
wire            n3262;
wire     [19:0] n3265;
wire            n3266;
wire     [19:0] n3269;
wire            n327;
wire            n3270;
wire     [19:0] n3273;
wire     [19:0] n3274;
wire     [19:0] n3275;
wire     [19:0] n3276;
wire     [19:0] n3277;
wire     [19:0] n3278;
wire            n328;
wire     [19:0] n3280;
wire            n3281;
wire      [3:0] n3282;
wire     [19:0] n3285;
wire            n3286;
wire     [19:0] n3289;
wire            n329;
wire            n3290;
wire     [19:0] n3293;
wire            n3294;
wire     [19:0] n3297;
wire     [19:0] n3298;
wire     [19:0] n3299;
wire            n33;
wire            n330;
wire     [19:0] n3300;
wire     [19:0] n3301;
wire     [19:0] n3302;
wire     [19:0] n3304;
wire            n3305;
wire      [3:0] n3306;
wire     [19:0] n3309;
wire            n331;
wire            n3310;
wire     [19:0] n3313;
wire            n3314;
wire     [19:0] n3317;
wire            n3318;
wire            n332;
wire     [19:0] n3321;
wire     [19:0] n3322;
wire     [19:0] n3323;
wire     [19:0] n3324;
wire     [19:0] n3325;
wire     [19:0] n3326;
wire     [19:0] n3328;
wire            n3329;
wire            n333;
wire      [3:0] n3330;
wire     [19:0] n3333;
wire            n3334;
wire     [19:0] n3337;
wire            n3338;
wire            n334;
wire     [19:0] n3341;
wire            n3342;
wire     [19:0] n3345;
wire     [19:0] n3346;
wire     [19:0] n3347;
wire     [19:0] n3348;
wire     [19:0] n3349;
wire            n335;
wire     [19:0] n3350;
wire     [19:0] n3352;
wire            n3353;
wire      [3:0] n3354;
wire     [19:0] n3357;
wire            n3358;
wire            n336;
wire     [19:0] n3361;
wire            n3362;
wire     [19:0] n3365;
wire            n3366;
wire     [19:0] n3369;
wire            n337;
wire     [19:0] n3370;
wire     [19:0] n3371;
wire     [19:0] n3372;
wire     [19:0] n3373;
wire     [19:0] n3374;
wire     [19:0] n3376;
wire     [19:0] n3377;
wire     [31:0] n3378;
wire            n338;
wire      [7:0] n3381;
wire     [19:0] n3382;
wire     [19:0] n3384;
wire            n3385;
wire      [3:0] n3386;
wire     [19:0] n3389;
wire            n339;
wire            n3390;
wire     [19:0] n3393;
wire            n3394;
wire     [19:0] n3397;
wire            n3398;
wire            n34;
wire            n340;
wire     [19:0] n3401;
wire     [19:0] n3402;
wire     [19:0] n3403;
wire     [19:0] n3404;
wire     [19:0] n3405;
wire            n3406;
wire      [3:0] n3407;
wire            n341;
wire     [19:0] n3410;
wire            n3411;
wire     [19:0] n3414;
wire            n3415;
wire     [19:0] n3418;
wire            n3419;
wire            n342;
wire     [19:0] n3422;
wire     [19:0] n3423;
wire     [19:0] n3424;
wire     [19:0] n3425;
wire     [19:0] n3426;
wire            n3427;
wire            n343;
wire     [19:0] n3430;
wire            n3431;
wire     [19:0] n3434;
wire            n3435;
wire     [19:0] n3438;
wire            n3439;
wire            n344;
wire     [19:0] n3442;
wire     [19:0] n3443;
wire     [19:0] n3444;
wire     [19:0] n3445;
wire     [19:0] n3446;
wire     [19:0] n3447;
wire     [19:0] n3449;
wire      [2:0] n345;
wire            n3450;
wire      [3:0] n3451;
wire     [19:0] n3454;
wire            n3455;
wire     [19:0] n3458;
wire            n3459;
wire      [5:0] n346;
wire     [19:0] n3462;
wire            n3463;
wire     [19:0] n3466;
wire     [19:0] n3467;
wire     [19:0] n3468;
wire     [19:0] n3469;
wire     [15:0] n347;
wire     [19:0] n3470;
wire            n3471;
wire     [19:0] n3474;
wire            n3475;
wire     [19:0] n3478;
wire            n3479;
wire      [4:0] n348;
wire     [19:0] n3482;
wire            n3483;
wire     [19:0] n3486;
wire     [19:0] n3487;
wire     [19:0] n3488;
wire     [19:0] n3489;
wire            n349;
wire     [19:0] n3490;
wire     [19:0] n3491;
wire     [19:0] n3493;
wire            n3494;
wire      [3:0] n3495;
wire     [19:0] n3498;
wire            n3499;
wire            n35;
wire            n350;
wire     [19:0] n3502;
wire            n3503;
wire     [19:0] n3506;
wire            n3507;
wire            n351;
wire     [19:0] n3510;
wire     [19:0] n3511;
wire     [19:0] n3512;
wire     [19:0] n3513;
wire     [19:0] n3514;
wire     [19:0] n3515;
wire     [19:0] n3517;
wire            n3518;
wire      [3:0] n3519;
wire            n352;
wire     [19:0] n3522;
wire            n3523;
wire     [19:0] n3526;
wire            n3527;
wire            n353;
wire     [19:0] n3530;
wire            n3531;
wire     [19:0] n3534;
wire     [19:0] n3535;
wire     [19:0] n3536;
wire     [19:0] n3537;
wire     [19:0] n3538;
wire     [19:0] n3539;
wire     [19:0] n3541;
wire            n3542;
wire      [3:0] n3543;
wire     [19:0] n3546;
wire            n3547;
wire     [31:0] n355;
wire     [19:0] n3550;
wire            n3551;
wire     [19:0] n3554;
wire            n3555;
wire     [19:0] n3558;
wire     [19:0] n3559;
wire     [19:0] n3560;
wire     [19:0] n3561;
wire     [19:0] n3562;
wire     [19:0] n3563;
wire     [19:0] n3565;
wire            n3566;
wire      [3:0] n3567;
wire     [31:0] n357;
wire     [19:0] n3570;
wire            n3571;
wire     [19:0] n3574;
wire            n3575;
wire     [19:0] n3578;
wire            n3579;
wire     [19:0] n3582;
wire     [19:0] n3583;
wire     [19:0] n3584;
wire     [19:0] n3585;
wire     [19:0] n3586;
wire     [19:0] n3587;
wire     [19:0] n3589;
wire     [31:0] n359;
wire     [19:0] n3590;
wire     [31:0] n3591;
wire      [7:0] n3594;
wire     [19:0] n3595;
wire     [19:0] n3597;
wire            n3598;
wire      [3:0] n3599;
wire            n36;
wire     [19:0] n3602;
wire            n3603;
wire     [19:0] n3606;
wire            n3607;
wire     [31:0] n361;
wire     [19:0] n3610;
wire            n3611;
wire     [19:0] n3614;
wire     [19:0] n3615;
wire     [19:0] n3616;
wire     [19:0] n3617;
wire     [19:0] n3618;
wire            n3619;
wire      [3:0] n3620;
wire     [19:0] n3623;
wire            n3624;
wire     [19:0] n3627;
wire            n3628;
wire     [31:0] n363;
wire     [19:0] n3631;
wire            n3632;
wire     [19:0] n3635;
wire     [19:0] n3636;
wire     [19:0] n3637;
wire     [19:0] n3638;
wire     [19:0] n3639;
wire            n3640;
wire     [19:0] n3643;
wire            n3644;
wire     [19:0] n3647;
wire            n3648;
wire     [31:0] n365;
wire     [19:0] n3651;
wire            n3652;
wire     [19:0] n3655;
wire     [19:0] n3656;
wire     [19:0] n3657;
wire     [19:0] n3658;
wire     [19:0] n3659;
wire     [19:0] n3660;
wire     [19:0] n3662;
wire            n3663;
wire      [3:0] n3664;
wire     [19:0] n3667;
wire            n3668;
wire     [31:0] n367;
wire     [19:0] n3671;
wire            n3672;
wire     [19:0] n3675;
wire            n3676;
wire     [19:0] n3679;
wire     [19:0] n3680;
wire     [19:0] n3681;
wire     [19:0] n3682;
wire     [19:0] n3683;
wire            n3684;
wire     [19:0] n3687;
wire            n3688;
wire     [31:0] n369;
wire     [19:0] n3691;
wire            n3692;
wire     [19:0] n3695;
wire            n3696;
wire     [19:0] n3699;
wire            n37;
wire     [19:0] n3700;
wire     [19:0] n3701;
wire     [19:0] n3702;
wire     [19:0] n3703;
wire     [19:0] n3704;
wire     [19:0] n3706;
wire            n3707;
wire      [3:0] n3708;
wire     [31:0] n371;
wire     [19:0] n3711;
wire            n3712;
wire     [19:0] n3715;
wire            n3716;
wire     [19:0] n3719;
wire            n3720;
wire     [19:0] n3723;
wire     [19:0] n3724;
wire     [19:0] n3725;
wire     [19:0] n3726;
wire     [19:0] n3727;
wire     [19:0] n3728;
wire     [31:0] n373;
wire     [19:0] n3730;
wire            n3731;
wire      [3:0] n3732;
wire     [19:0] n3735;
wire            n3736;
wire     [19:0] n3739;
wire            n3740;
wire     [19:0] n3743;
wire            n3744;
wire     [19:0] n3747;
wire     [19:0] n3748;
wire     [19:0] n3749;
wire     [31:0] n375;
wire     [19:0] n3750;
wire     [19:0] n3751;
wire     [19:0] n3752;
wire     [19:0] n3754;
wire            n3755;
wire      [3:0] n3756;
wire     [19:0] n3759;
wire            n3760;
wire     [19:0] n3763;
wire            n3764;
wire     [19:0] n3767;
wire            n3768;
wire     [31:0] n377;
wire     [19:0] n3771;
wire     [19:0] n3772;
wire     [19:0] n3773;
wire     [19:0] n3774;
wire     [19:0] n3775;
wire     [19:0] n3776;
wire     [19:0] n3778;
wire            n3779;
wire      [3:0] n3780;
wire     [19:0] n3783;
wire            n3784;
wire     [19:0] n3787;
wire            n3788;
wire     [31:0] n379;
wire     [19:0] n3791;
wire            n3792;
wire     [19:0] n3795;
wire     [19:0] n3796;
wire     [19:0] n3797;
wire     [19:0] n3798;
wire     [19:0] n3799;
wire            n38;
wire     [19:0] n3800;
wire     [19:0] n3802;
wire     [19:0] n3803;
wire     [31:0] n3804;
wire      [7:0] n3807;
wire     [19:0] n3808;
wire     [31:0] n381;
wire     [19:0] n3810;
wire            n3811;
wire      [3:0] n3812;
wire     [19:0] n3815;
wire            n3816;
wire     [19:0] n3819;
wire            n3820;
wire     [19:0] n3823;
wire            n3824;
wire     [19:0] n3827;
wire     [19:0] n3828;
wire     [19:0] n3829;
wire     [31:0] n383;
wire     [19:0] n3830;
wire     [19:0] n3831;
wire            n3832;
wire      [3:0] n3833;
wire     [19:0] n3836;
wire            n3837;
wire     [19:0] n3840;
wire            n3841;
wire     [19:0] n3844;
wire            n3845;
wire     [19:0] n3848;
wire     [19:0] n3849;
wire     [31:0] n385;
wire     [19:0] n3850;
wire     [19:0] n3851;
wire     [19:0] n3852;
wire            n3853;
wire     [19:0] n3856;
wire            n3857;
wire     [19:0] n3860;
wire            n3861;
wire     [19:0] n3864;
wire            n3865;
wire     [19:0] n3868;
wire     [19:0] n3869;
wire     [31:0] n387;
wire     [19:0] n3870;
wire     [19:0] n3871;
wire     [19:0] n3872;
wire     [19:0] n3873;
wire     [19:0] n3875;
wire            n3876;
wire      [3:0] n3877;
wire     [19:0] n3880;
wire            n3881;
wire     [19:0] n3884;
wire            n3885;
wire     [19:0] n3888;
wire            n3889;
wire     [31:0] n389;
wire     [19:0] n3892;
wire     [19:0] n3893;
wire     [19:0] n3894;
wire     [19:0] n3895;
wire     [19:0] n3896;
wire            n3897;
wire            n39;
wire            n390;
wire     [19:0] n3900;
wire            n3901;
wire     [19:0] n3904;
wire            n3905;
wire     [19:0] n3908;
wire            n3909;
wire     [19:0] n3912;
wire     [19:0] n3913;
wire     [19:0] n3914;
wire     [19:0] n3915;
wire     [19:0] n3916;
wire     [19:0] n3917;
wire     [19:0] n3919;
wire     [31:0] n392;
wire            n3920;
wire      [3:0] n3921;
wire     [19:0] n3924;
wire            n3925;
wire     [19:0] n3928;
wire            n3929;
wire     [19:0] n3932;
wire            n3933;
wire     [19:0] n3936;
wire     [19:0] n3937;
wire     [19:0] n3938;
wire     [19:0] n3939;
wire     [31:0] n394;
wire     [19:0] n3940;
wire     [19:0] n3941;
wire     [19:0] n3943;
wire            n3944;
wire      [3:0] n3945;
wire     [19:0] n3948;
wire            n3949;
wire     [31:0] n395;
wire     [19:0] n3952;
wire            n3953;
wire     [19:0] n3956;
wire            n3957;
wire     [31:0] n396;
wire     [19:0] n3960;
wire     [19:0] n3961;
wire     [19:0] n3962;
wire     [19:0] n3963;
wire     [19:0] n3964;
wire     [19:0] n3965;
wire     [19:0] n3967;
wire            n3968;
wire      [3:0] n3969;
wire     [31:0] n397;
wire     [19:0] n3972;
wire            n3973;
wire     [19:0] n3976;
wire            n3977;
wire      [1:0] n398;
wire     [19:0] n3980;
wire            n3981;
wire     [19:0] n3984;
wire     [19:0] n3985;
wire     [19:0] n3986;
wire     [19:0] n3987;
wire     [19:0] n3988;
wire     [19:0] n3989;
wire     [19:0] n3991;
wire            n3992;
wire      [3:0] n3993;
wire     [19:0] n3996;
wire            n3997;
wire            n4;
wire            n40;
wire            n400;
wire     [19:0] n4000;
wire            n4001;
wire     [19:0] n4004;
wire            n4005;
wire     [19:0] n4008;
wire     [19:0] n4009;
wire     [19:0] n4010;
wire     [19:0] n4011;
wire     [19:0] n4012;
wire     [19:0] n4013;
wire     [19:0] n4015;
wire     [19:0] n4016;
wire     [31:0] n4017;
wire      [7:0] n4020;
wire     [19:0] n4021;
wire     [19:0] n4023;
wire            n4024;
wire      [3:0] n4025;
wire     [19:0] n4028;
wire            n4029;
wire      [3:0] n403;
wire     [19:0] n4032;
wire            n4033;
wire     [19:0] n4036;
wire            n4037;
wire     [19:0] n4040;
wire     [19:0] n4041;
wire     [19:0] n4042;
wire     [19:0] n4043;
wire     [19:0] n4044;
wire            n4045;
wire      [3:0] n4046;
wire     [19:0] n4049;
wire            n4050;
wire     [19:0] n4053;
wire            n4054;
wire     [19:0] n4057;
wire            n4058;
wire     [19:0] n406;
wire     [19:0] n4061;
wire     [19:0] n4062;
wire     [19:0] n4063;
wire     [19:0] n4064;
wire     [19:0] n4065;
wire            n4066;
wire     [19:0] n4069;
wire            n407;
wire            n4070;
wire     [19:0] n4073;
wire            n4074;
wire     [19:0] n4077;
wire            n4078;
wire     [19:0] n4081;
wire     [19:0] n4082;
wire     [19:0] n4083;
wire     [19:0] n4084;
wire     [19:0] n4085;
wire     [19:0] n4086;
wire     [19:0] n4088;
wire            n4089;
wire      [3:0] n4090;
wire     [19:0] n4093;
wire            n4094;
wire     [19:0] n4097;
wire            n4098;
wire     [19:0] n410;
wire     [19:0] n4101;
wire            n4102;
wire     [19:0] n4105;
wire     [19:0] n4106;
wire     [19:0] n4107;
wire     [19:0] n4108;
wire     [19:0] n4109;
wire            n411;
wire            n4110;
wire     [19:0] n4113;
wire            n4114;
wire     [19:0] n4117;
wire            n4118;
wire     [19:0] n4121;
wire            n4122;
wire     [19:0] n4125;
wire     [19:0] n4126;
wire     [19:0] n4127;
wire     [19:0] n4128;
wire     [19:0] n4129;
wire     [19:0] n4130;
wire     [19:0] n4132;
wire            n4133;
wire      [3:0] n4134;
wire     [19:0] n4137;
wire            n4138;
wire     [19:0] n414;
wire     [19:0] n4141;
wire            n4142;
wire     [19:0] n4145;
wire            n4146;
wire     [19:0] n4149;
wire            n415;
wire     [19:0] n4150;
wire     [19:0] n4151;
wire     [19:0] n4152;
wire     [19:0] n4153;
wire     [19:0] n4154;
wire     [19:0] n4156;
wire            n4157;
wire      [3:0] n4158;
wire     [19:0] n4161;
wire            n4162;
wire     [19:0] n4165;
wire            n4166;
wire     [19:0] n4169;
wire            n4170;
wire     [19:0] n4173;
wire     [19:0] n4174;
wire     [19:0] n4175;
wire     [19:0] n4176;
wire     [19:0] n4177;
wire     [19:0] n4178;
wire     [19:0] n418;
wire     [19:0] n4180;
wire            n4181;
wire      [3:0] n4182;
wire     [19:0] n4185;
wire            n4186;
wire     [19:0] n4189;
wire            n4190;
wire     [19:0] n4193;
wire            n4194;
wire     [19:0] n4197;
wire     [19:0] n4198;
wire     [19:0] n4199;
wire            n42;
wire     [19:0] n420;
wire     [19:0] n4200;
wire     [19:0] n4201;
wire     [19:0] n4202;
wire     [19:0] n4204;
wire            n4205;
wire      [3:0] n4206;
wire     [19:0] n4209;
wire     [19:0] n421;
wire            n4210;
wire     [19:0] n4213;
wire            n4214;
wire     [19:0] n4217;
wire            n4218;
wire     [19:0] n422;
wire     [19:0] n4221;
wire     [19:0] n4222;
wire     [19:0] n4223;
wire     [19:0] n4224;
wire     [19:0] n4225;
wire     [19:0] n4226;
wire     [19:0] n4228;
wire     [19:0] n4229;
wire     [19:0] n423;
wire     [31:0] n4230;
wire      [7:0] n4233;
wire     [19:0] n4234;
wire     [19:0] n4236;
wire            n4237;
wire      [3:0] n4238;
wire      [7:0] n424;
wire     [19:0] n4241;
wire            n4242;
wire     [19:0] n4245;
wire            n4246;
wire     [19:0] n4249;
wire            n4250;
wire     [19:0] n4253;
wire     [19:0] n4254;
wire     [19:0] n4255;
wire     [19:0] n4256;
wire     [19:0] n4257;
wire            n4258;
wire      [3:0] n4259;
wire      [7:0] n426;
wire     [19:0] n4262;
wire            n4263;
wire     [19:0] n4266;
wire            n4267;
wire     [31:0] n427;
wire     [19:0] n4270;
wire            n4271;
wire     [19:0] n4274;
wire     [19:0] n4275;
wire     [19:0] n4276;
wire     [19:0] n4277;
wire     [19:0] n4278;
wire            n4279;
wire            n428;
wire     [19:0] n4282;
wire            n4283;
wire     [19:0] n4286;
wire            n4287;
wire     [19:0] n4290;
wire            n4291;
wire     [19:0] n4294;
wire     [19:0] n4295;
wire     [19:0] n4296;
wire     [19:0] n4297;
wire     [19:0] n4298;
wire     [19:0] n4299;
wire            n43;
wire      [3:0] n430;
wire     [19:0] n4301;
wire            n4302;
wire      [3:0] n4303;
wire     [19:0] n4306;
wire            n4307;
wire     [19:0] n4310;
wire            n4311;
wire     [19:0] n4314;
wire            n4315;
wire     [19:0] n4318;
wire     [19:0] n4319;
wire     [19:0] n4320;
wire     [19:0] n4321;
wire     [19:0] n4322;
wire            n4323;
wire     [19:0] n4326;
wire            n4327;
wire     [19:0] n433;
wire     [19:0] n4330;
wire            n4331;
wire     [19:0] n4334;
wire            n4335;
wire     [19:0] n4338;
wire     [19:0] n4339;
wire            n434;
wire     [19:0] n4340;
wire     [19:0] n4341;
wire     [19:0] n4342;
wire     [19:0] n4343;
wire     [19:0] n4345;
wire            n4346;
wire      [3:0] n4347;
wire     [19:0] n4350;
wire            n4351;
wire     [19:0] n4354;
wire            n4355;
wire     [19:0] n4358;
wire            n4359;
wire     [19:0] n4362;
wire     [19:0] n4363;
wire     [19:0] n4364;
wire     [19:0] n4365;
wire     [19:0] n4366;
wire     [19:0] n4367;
wire     [19:0] n4369;
wire     [19:0] n437;
wire            n4370;
wire      [3:0] n4371;
wire     [19:0] n4374;
wire            n4375;
wire     [19:0] n4378;
wire            n4379;
wire            n438;
wire     [19:0] n4382;
wire            n4383;
wire     [19:0] n4386;
wire     [19:0] n4387;
wire     [19:0] n4388;
wire     [19:0] n4389;
wire     [19:0] n4390;
wire     [19:0] n4391;
wire     [19:0] n4393;
wire            n4394;
wire      [3:0] n4395;
wire     [19:0] n4398;
wire            n4399;
wire            n44;
wire     [19:0] n4402;
wire            n4403;
wire     [19:0] n4406;
wire            n4407;
wire     [19:0] n441;
wire     [19:0] n4410;
wire     [19:0] n4411;
wire     [19:0] n4412;
wire     [19:0] n4413;
wire     [19:0] n4414;
wire     [19:0] n4415;
wire     [19:0] n4417;
wire            n4418;
wire      [3:0] n4419;
wire            n442;
wire     [19:0] n4422;
wire            n4423;
wire     [19:0] n4426;
wire            n4427;
wire     [19:0] n4430;
wire            n4431;
wire     [19:0] n4434;
wire     [19:0] n4435;
wire     [19:0] n4436;
wire     [19:0] n4437;
wire     [19:0] n4438;
wire     [19:0] n4439;
wire     [19:0] n4441;
wire     [19:0] n445;
wire     [19:0] n446;
wire     [19:0] n447;
wire     [19:0] n448;
wire     [19:0] n449;
wire      [7:0] n450;
wire      [7:0] n452;
wire     [31:0] n453;
wire            n454;
wire      [3:0] n455;
wire     [19:0] n458;
wire            n459;
wire            n46;
wire     [19:0] n462;
wire            n463;
wire     [19:0] n466;
wire            n467;
wire            n47;
wire     [19:0] n470;
wire     [19:0] n471;
wire     [19:0] n472;
wire     [19:0] n473;
wire     [19:0] n474;
wire      [7:0] n475;
wire      [7:0] n477;
wire     [31:0] n478;
wire            n479;
wire      [3:0] n480;
wire     [19:0] n483;
wire            n484;
wire     [19:0] n487;
wire            n488;
wire            n49;
wire     [19:0] n491;
wire            n492;
wire     [19:0] n495;
wire     [19:0] n496;
wire     [19:0] n497;
wire     [19:0] n498;
wire     [19:0] n499;
wire            n5;
wire      [7:0] n500;
wire      [7:0] n502;
wire     [31:0] n503;
wire            n504;
wire      [3:0] n505;
wire     [19:0] n508;
wire            n509;
wire            n51;
wire     [19:0] n512;
wire            n513;
wire     [19:0] n516;
wire            n517;
wire     [19:0] n520;
wire     [19:0] n521;
wire     [19:0] n522;
wire     [19:0] n523;
wire     [19:0] n524;
wire      [7:0] n525;
wire      [7:0] n527;
wire     [31:0] n528;
wire            n529;
wire            n53;
wire      [3:0] n530;
wire     [19:0] n533;
wire            n534;
wire     [19:0] n537;
wire            n538;
wire     [19:0] n541;
wire            n542;
wire     [19:0] n545;
wire     [19:0] n546;
wire     [19:0] n547;
wire     [19:0] n548;
wire     [19:0] n549;
wire            n55;
wire      [7:0] n550;
wire      [7:0] n552;
wire     [31:0] n553;
wire            n554;
wire      [3:0] n555;
wire     [19:0] n558;
wire            n559;
wire     [19:0] n562;
wire            n563;
wire     [19:0] n566;
wire            n567;
wire            n57;
wire     [19:0] n570;
wire     [19:0] n571;
wire     [19:0] n572;
wire     [19:0] n573;
wire     [19:0] n574;
wire      [7:0] n575;
wire      [7:0] n577;
wire     [31:0] n578;
wire            n579;
wire      [3:0] n580;
wire     [19:0] n583;
wire            n584;
wire     [19:0] n587;
wire            n588;
wire            n59;
wire     [19:0] n591;
wire            n592;
wire     [19:0] n595;
wire     [19:0] n596;
wire     [19:0] n597;
wire     [19:0] n598;
wire     [19:0] n599;
wire            n6;
wire      [7:0] n600;
wire      [7:0] n602;
wire     [31:0] n603;
wire            n604;
wire      [3:0] n605;
wire     [19:0] n608;
wire            n609;
wire            n61;
wire     [19:0] n612;
wire            n613;
wire     [19:0] n616;
wire            n617;
wire     [19:0] n620;
wire     [19:0] n621;
wire     [19:0] n622;
wire     [19:0] n623;
wire     [19:0] n624;
wire      [7:0] n625;
wire      [7:0] n627;
wire     [31:0] n628;
wire            n629;
wire            n63;
wire      [3:0] n631;
wire     [19:0] n634;
wire            n635;
wire     [19:0] n638;
wire            n639;
wire     [19:0] n642;
wire            n643;
wire     [19:0] n646;
wire     [19:0] n647;
wire     [19:0] n648;
wire     [19:0] n649;
wire            n65;
wire     [19:0] n650;
wire      [7:0] n651;
wire      [7:0] n653;
wire     [31:0] n654;
wire            n655;
wire      [3:0] n657;
wire     [19:0] n660;
wire            n661;
wire     [19:0] n664;
wire            n665;
wire     [19:0] n668;
wire            n669;
wire            n67;
wire     [19:0] n672;
wire     [19:0] n673;
wire     [19:0] n674;
wire     [19:0] n675;
wire     [19:0] n676;
wire      [7:0] n677;
wire      [7:0] n679;
wire     [31:0] n680;
wire            n681;
wire      [3:0] n682;
wire     [19:0] n685;
wire            n686;
wire     [19:0] n689;
wire            n69;
wire            n690;
wire     [19:0] n693;
wire            n694;
wire     [19:0] n697;
wire     [19:0] n698;
wire     [19:0] n699;
wire            n7;
wire     [19:0] n700;
wire     [19:0] n701;
wire      [7:0] n702;
wire      [7:0] n704;
wire     [31:0] n705;
wire            n706;
wire      [3:0] n707;
wire            n71;
wire     [19:0] n710;
wire            n711;
wire     [19:0] n714;
wire            n715;
wire     [19:0] n718;
wire            n719;
wire     [19:0] n722;
wire     [19:0] n723;
wire     [19:0] n724;
wire     [19:0] n725;
wire     [19:0] n726;
wire      [7:0] n727;
wire      [7:0] n729;
wire            n73;
wire     [31:0] n730;
wire            n731;
wire      [3:0] n732;
wire     [19:0] n735;
wire            n736;
wire     [19:0] n739;
wire            n740;
wire     [19:0] n743;
wire            n744;
wire     [19:0] n747;
wire     [19:0] n748;
wire     [19:0] n749;
wire            n75;
wire     [19:0] n750;
wire     [19:0] n751;
wire      [7:0] n752;
wire      [7:0] n754;
wire     [31:0] n755;
wire            n756;
wire      [3:0] n757;
wire     [19:0] n760;
wire            n761;
wire     [19:0] n764;
wire            n765;
wire     [19:0] n768;
wire            n769;
wire            n77;
wire     [19:0] n772;
wire     [19:0] n773;
wire     [19:0] n774;
wire     [19:0] n775;
wire     [19:0] n776;
wire      [7:0] n777;
wire      [7:0] n779;
wire     [31:0] n780;
wire            n781;
wire      [3:0] n782;
wire     [19:0] n785;
wire            n786;
wire     [19:0] n789;
wire            n79;
wire            n790;
wire     [19:0] n793;
wire            n794;
wire     [19:0] n797;
wire     [19:0] n798;
wire     [19:0] n799;
wire            n8;
wire     [19:0] n800;
wire     [19:0] n801;
wire      [7:0] n802;
wire      [7:0] n804;
wire      [5:0] n805;
wire      [5:0] n806;
wire      [5:0] n807;
wire      [5:0] n808;
wire      [5:0] n809;
wire            n81;
wire      [5:0] n810;
wire      [5:0] n811;
wire      [5:0] n812;
wire      [5:0] n813;
wire      [5:0] n814;
wire      [5:0] n815;
wire      [5:0] n816;
wire      [5:0] n817;
wire      [5:0] n818;
wire      [5:0] n819;
wire      [5:0] n820;
wire      [5:0] n821;
wire      [5:0] n822;
wire      [5:0] n823;
wire      [5:0] n824;
wire      [5:0] n825;
wire      [5:0] n826;
wire      [5:0] n827;
wire      [5:0] n828;
wire            n829;
wire            n83;
wire            n830;
wire      [7:0] n831;
wire      [7:0] n832;
wire      [7:0] n833;
wire            n834;
wire            n835;
wire      [7:0] n836;
wire      [7:0] n837;
wire      [7:0] n838;
wire            n839;
wire            n840;
wire      [7:0] n841;
wire      [7:0] n842;
wire      [7:0] n843;
wire            n844;
wire            n845;
wire      [7:0] n846;
wire      [7:0] n847;
wire      [7:0] n848;
wire            n849;
wire            n85;
wire            n850;
wire      [7:0] n851;
wire      [7:0] n852;
wire      [7:0] n853;
wire            n854;
wire            n855;
wire      [7:0] n856;
wire      [7:0] n857;
wire      [7:0] n858;
wire            n859;
wire            n860;
wire      [7:0] n861;
wire      [7:0] n862;
wire      [7:0] n863;
wire            n864;
wire            n865;
wire      [7:0] n866;
wire      [7:0] n867;
wire      [7:0] n868;
wire            n869;
wire            n87;
wire            n870;
wire      [7:0] n871;
wire      [7:0] n872;
wire      [7:0] n873;
wire            n874;
wire            n875;
wire      [7:0] n876;
wire      [7:0] n877;
wire      [7:0] n878;
wire            n879;
wire            n880;
wire      [7:0] n881;
wire      [7:0] n882;
wire      [7:0] n883;
wire            n884;
wire            n885;
wire      [7:0] n886;
wire      [7:0] n887;
wire      [7:0] n888;
wire            n889;
wire            n89;
wire            n890;
wire            n891;
wire      [3:0] n892;
wire     [19:0] n893;
wire      [3:0] n894;
wire     [19:0] n895;
wire      [3:0] n896;
wire     [19:0] n897;
wire      [3:0] n898;
wire     [19:0] n899;
wire      [3:0] n900;
wire     [19:0] n901;
wire      [3:0] n902;
wire     [19:0] n903;
wire      [3:0] n904;
wire     [19:0] n905;
wire      [3:0] n906;
wire     [19:0] n907;
wire      [3:0] n908;
wire     [19:0] n909;
wire            n91;
wire      [3:0] n910;
wire     [19:0] n911;
wire      [3:0] n912;
wire     [19:0] n913;
wire      [3:0] n914;
wire     [19:0] n915;
wire      [3:0] n916;
wire     [19:0] n917;
wire      [3:0] n918;
wire     [19:0] n919;
wire      [3:0] n920;
wire     [19:0] n921;
wire      [3:0] n922;
wire     [19:0] n923;
wire            n924;
wire            n925;
wire            n926;
wire      [3:0] n927;
wire     [19:0] n928;
wire      [3:0] n929;
wire            n93;
wire     [19:0] n930;
wire      [3:0] n931;
wire     [19:0] n932;
wire      [3:0] n933;
wire     [19:0] n934;
wire      [3:0] n935;
wire     [19:0] n936;
wire      [3:0] n937;
wire     [19:0] n938;
wire      [3:0] n939;
wire     [19:0] n940;
wire      [3:0] n941;
wire     [19:0] n942;
wire      [3:0] n943;
wire     [19:0] n944;
wire      [3:0] n945;
wire     [19:0] n946;
wire      [3:0] n947;
wire     [19:0] n948;
wire      [3:0] n949;
wire            n95;
wire     [19:0] n950;
wire      [3:0] n951;
wire     [19:0] n952;
wire      [3:0] n953;
wire     [19:0] n954;
wire      [3:0] n955;
wire     [19:0] n956;
wire      [3:0] n957;
wire     [19:0] n958;
wire            n959;
wire            n960;
wire            n961;
wire      [3:0] n962;
wire     [19:0] n963;
wire      [3:0] n964;
wire     [19:0] n965;
wire      [3:0] n966;
wire     [19:0] n967;
wire      [3:0] n968;
wire     [19:0] n969;
wire            n97;
wire      [3:0] n970;
wire     [19:0] n971;
wire      [3:0] n972;
wire     [19:0] n973;
wire      [3:0] n974;
wire     [19:0] n975;
wire      [3:0] n976;
wire     [19:0] n977;
wire      [3:0] n978;
wire     [19:0] n979;
wire      [3:0] n980;
wire     [19:0] n981;
wire      [3:0] n982;
wire     [19:0] n983;
wire      [3:0] n984;
wire     [19:0] n985;
wire      [3:0] n986;
wire     [19:0] n987;
wire      [3:0] n988;
wire     [19:0] n989;
wire            n99;
wire      [3:0] n990;
wire     [19:0] n991;
wire      [3:0] n992;
wire     [19:0] n993;
wire            n994;
wire            n995;
wire            n996;
wire      [3:0] n997;
wire     [19:0] n998;
wire      [3:0] n999;
wire            output_port_ready;
wire     [31:0] pe0_act_buffer_addr0;
wire     [31:0] pe0_act_buffer_addr1;
wire     [31:0] pe0_act_buffer_addr10;
wire     [31:0] pe0_act_buffer_addr11;
wire     [31:0] pe0_act_buffer_addr12;
wire     [31:0] pe0_act_buffer_addr13;
wire     [31:0] pe0_act_buffer_addr14;
wire     [31:0] pe0_act_buffer_addr15;
wire     [31:0] pe0_act_buffer_addr2;
wire     [31:0] pe0_act_buffer_addr3;
wire     [31:0] pe0_act_buffer_addr4;
wire     [31:0] pe0_act_buffer_addr5;
wire     [31:0] pe0_act_buffer_addr6;
wire     [31:0] pe0_act_buffer_addr7;
wire     [31:0] pe0_act_buffer_addr8;
wire     [31:0] pe0_act_buffer_addr9;
wire     [31:0] pe0_act_buffer_addr_n1035;
wire     [31:0] pe0_act_buffer_addr_n1249;
wire     [31:0] pe0_act_buffer_addr_n1462;
wire     [31:0] pe0_act_buffer_addr_n1675;
wire     [31:0] pe0_act_buffer_addr_n1888;
wire     [31:0] pe0_act_buffer_addr_n2101;
wire     [31:0] pe0_act_buffer_addr_n2314;
wire     [31:0] pe0_act_buffer_addr_n2527;
wire     [31:0] pe0_act_buffer_addr_n2740;
wire     [31:0] pe0_act_buffer_addr_n2953;
wire     [31:0] pe0_act_buffer_addr_n3166;
wire     [31:0] pe0_act_buffer_addr_n3379;
wire     [31:0] pe0_act_buffer_addr_n3592;
wire     [31:0] pe0_act_buffer_addr_n3805;
wire     [31:0] pe0_act_buffer_addr_n4018;
wire     [31:0] pe0_act_buffer_addr_n4231;
wire      [7:0] pe0_act_buffer_data0;
wire      [7:0] pe0_act_buffer_data1;
wire      [7:0] pe0_act_buffer_data10;
wire      [7:0] pe0_act_buffer_data11;
wire      [7:0] pe0_act_buffer_data12;
wire      [7:0] pe0_act_buffer_data13;
wire      [7:0] pe0_act_buffer_data14;
wire      [7:0] pe0_act_buffer_data15;
wire      [7:0] pe0_act_buffer_data2;
wire      [7:0] pe0_act_buffer_data3;
wire      [7:0] pe0_act_buffer_data4;
wire      [7:0] pe0_act_buffer_data5;
wire      [7:0] pe0_act_buffer_data6;
wire      [7:0] pe0_act_buffer_data7;
wire      [7:0] pe0_act_buffer_data8;
wire      [7:0] pe0_act_buffer_data9;
wire      [7:0] pe0_act_buffer_data_n1036;
wire      [7:0] pe0_act_buffer_data_n1250;
wire      [7:0] pe0_act_buffer_data_n1463;
wire      [7:0] pe0_act_buffer_data_n1676;
wire      [7:0] pe0_act_buffer_data_n1889;
wire      [7:0] pe0_act_buffer_data_n2102;
wire      [7:0] pe0_act_buffer_data_n2315;
wire      [7:0] pe0_act_buffer_data_n2528;
wire      [7:0] pe0_act_buffer_data_n2741;
wire      [7:0] pe0_act_buffer_data_n2954;
wire      [7:0] pe0_act_buffer_data_n3167;
wire      [7:0] pe0_act_buffer_data_n3380;
wire      [7:0] pe0_act_buffer_data_n3593;
wire      [7:0] pe0_act_buffer_data_n3806;
wire      [7:0] pe0_act_buffer_data_n4019;
wire      [7:0] pe0_act_buffer_data_n4232;
wire            pe0_act_buffer_wen0;
wire            pe0_act_buffer_wen1;
wire            pe0_act_buffer_wen10;
wire            pe0_act_buffer_wen11;
wire            pe0_act_buffer_wen12;
wire            pe0_act_buffer_wen13;
wire            pe0_act_buffer_wen14;
wire            pe0_act_buffer_wen15;
wire            pe0_act_buffer_wen2;
wire            pe0_act_buffer_wen3;
wire            pe0_act_buffer_wen4;
wire            pe0_act_buffer_wen5;
wire            pe0_act_buffer_wen6;
wire            pe0_act_buffer_wen7;
wire            pe0_act_buffer_wen8;
wire            pe0_act_buffer_wen9;
wire            pe0_act_reg_port_valid;
wire            rst;
wire            rva_in_valid;
wire     [15:0] wstrb;
assign __ILA_pe_act_valid__ = 1'b1 ;
assign bv_1_1_n0 = 1'h1 ;
assign n1 =  ( axi_rw ) == ( bv_1_1_n0 )  ;
assign bv_24_8388624_n2 = 24'h800010 ;
assign n3 =  ( addr ) == ( bv_24_8388624_n2 )  ;
assign n4 =  ( rva_in_valid ) & ( rva_in_ready )  ;
assign n5 =  ( n4 ) == ( bv_1_1_n0 )  ;
assign n6 =  ( n3 ) & (n5 )  ;
assign n7 =  ( n1 ) & (n6 )  ;
assign __ILA_pe_act_decode_of_PE0_CONFIG_ACT_MNGR__ = n7 ;
assign __ILA_pe_act_acc_decode__[0] = __ILA_pe_act_decode_of_PE0_CONFIG_ACT_MNGR__ ;
assign n8 =  ( axi_rw ) == ( bv_1_1_n0 )  ;
assign bv_24_8388640_n9 = 24'h800020 ;
assign n10 =  ( addr ) == ( bv_24_8388640_n9 )  ;
assign n11 =  ( n4 ) == ( bv_1_1_n0 )  ;
assign n12 =  ( n10 ) & (n11 )  ;
assign n13 =  ( n8 ) & (n12 )  ;
assign __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_0_15__ = n13 ;
assign __ILA_pe_act_acc_decode__[1] = __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_0_15__ ;
assign n14 =  ( axi_rw ) == ( bv_1_1_n0 )  ;
assign bv_24_8388656_n15 = 24'h800030 ;
assign n16 =  ( addr ) == ( bv_24_8388656_n15 )  ;
assign n17 =  ( n4 ) == ( bv_1_1_n0 )  ;
assign n18 =  ( n16 ) & (n17 )  ;
assign n19 =  ( n14 ) & (n18 )  ;
assign __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_16_31__ = n19 ;
assign __ILA_pe_act_acc_decode__[2] = __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_16_31__ ;
assign n20 =  ( axi_rw ) == ( bv_1_1_n0 )  ;
assign bv_24_9437184_n21 = 24'h900000 ;
assign n22 =  ( addr ) == ( bv_24_9437184_n21 )  ;
assign n23 =  ( addr ) > ( bv_24_9437184_n21 )  ;
assign n24 =  ( n22 ) | ( n23 )  ;
assign bv_24_9437680_n25 = 24'h9001f0 ;
assign n26 =  ( addr ) == ( bv_24_9437680_n25 )  ;
assign n27 =  ( addr ) < ( bv_24_9437680_n25 )  ;
assign n28 =  ( n26 ) | ( n27 )  ;
assign n29 =  ( n24 ) & (n28 )  ;
assign n30 =  ( n20 ) & (n29 )  ;
assign __ILA_pe_act_decode_of_PE0_ACT_STORE_BUFFER__ = n30 ;
assign __ILA_pe_act_acc_decode__[3] = __ILA_pe_act_decode_of_PE0_ACT_STORE_BUFFER__ ;
assign n31 =  ( pe0_act_mngr_is_valid ) == ( bv_1_1_n0 )  ;
assign bv_1_0_n32 = 1'h0 ;
assign n33 =  ( pe0_act_is_start_reg ) == ( bv_1_0_n32 )  ;
assign n34 =  ( n31 ) & (n33 )  ;
assign n35 =  ( act_start ) == ( bv_1_1_n0 )  ;
assign n36 =  ( act_start_valid ) == ( bv_1_1_n0 )  ;
assign n37 =  ( n35 ) & (n36 )  ;
assign n38 =  ( act_start_ready ) == ( bv_1_1_n0 )  ;
assign n39 =  ( n37 ) & (n38 )  ;
assign n40 =  ( n34 ) & (n39 )  ;
assign bv_2_0_n41 = 2'h0 ;
assign n42 =  ( pe0_act_state ) == ( bv_2_0_n41 )  ;
assign n43 =  ( n40 ) & (n42 )  ;
assign __ILA_pe_act_decode_of_PE0_act_child_initiate__ = n43 ;
assign __ILA_pe_act_acc_decode__[4] = __ILA_pe_act_decode_of_PE0_act_child_initiate__ ;
assign n44 =  ( pe0_act_is_start_reg ) == ( bv_1_1_n0 )  ;
assign bv_2_1_n45 = 2'h1 ;
assign n46 =  ( pe0_act_state ) == ( bv_2_1_n45 )  ;
assign n47 =  ( n44 ) & (n46 )  ;
assign bv_6_31_n48 = 6'h1f ;
assign n49 =  ( pe0_act_instruction_counter ) == ( bv_6_31_n48 )  ;
assign bv_6_30_n50 = 6'h1e ;
assign n51 =  ( pe0_act_instruction_counter ) == ( bv_6_30_n50 )  ;
assign bv_6_29_n52 = 6'h1d ;
assign n53 =  ( pe0_act_instruction_counter ) == ( bv_6_29_n52 )  ;
assign bv_6_28_n54 = 6'h1c ;
assign n55 =  ( pe0_act_instruction_counter ) == ( bv_6_28_n54 )  ;
assign bv_6_27_n56 = 6'h1b ;
assign n57 =  ( pe0_act_instruction_counter ) == ( bv_6_27_n56 )  ;
assign bv_6_26_n58 = 6'h1a ;
assign n59 =  ( pe0_act_instruction_counter ) == ( bv_6_26_n58 )  ;
assign bv_6_25_n60 = 6'h19 ;
assign n61 =  ( pe0_act_instruction_counter ) == ( bv_6_25_n60 )  ;
assign bv_6_24_n62 = 6'h18 ;
assign n63 =  ( pe0_act_instruction_counter ) == ( bv_6_24_n62 )  ;
assign bv_6_23_n64 = 6'h17 ;
assign n65 =  ( pe0_act_instruction_counter ) == ( bv_6_23_n64 )  ;
assign bv_6_22_n66 = 6'h16 ;
assign n67 =  ( pe0_act_instruction_counter ) == ( bv_6_22_n66 )  ;
assign bv_6_21_n68 = 6'h15 ;
assign n69 =  ( pe0_act_instruction_counter ) == ( bv_6_21_n68 )  ;
assign bv_6_20_n70 = 6'h14 ;
assign n71 =  ( pe0_act_instruction_counter ) == ( bv_6_20_n70 )  ;
assign bv_6_19_n72 = 6'h13 ;
assign n73 =  ( pe0_act_instruction_counter ) == ( bv_6_19_n72 )  ;
assign bv_6_18_n74 = 6'h12 ;
assign n75 =  ( pe0_act_instruction_counter ) == ( bv_6_18_n74 )  ;
assign bv_6_17_n76 = 6'h11 ;
assign n77 =  ( pe0_act_instruction_counter ) == ( bv_6_17_n76 )  ;
assign bv_6_16_n78 = 6'h10 ;
assign n79 =  ( pe0_act_instruction_counter ) == ( bv_6_16_n78 )  ;
assign bv_6_15_n80 = 6'hf ;
assign n81 =  ( pe0_act_instruction_counter ) == ( bv_6_15_n80 )  ;
assign bv_6_14_n82 = 6'he ;
assign n83 =  ( pe0_act_instruction_counter ) == ( bv_6_14_n82 )  ;
assign bv_6_13_n84 = 6'hd ;
assign n85 =  ( pe0_act_instruction_counter ) == ( bv_6_13_n84 )  ;
assign bv_6_12_n86 = 6'hc ;
assign n87 =  ( pe0_act_instruction_counter ) == ( bv_6_12_n86 )  ;
assign bv_6_11_n88 = 6'hb ;
assign n89 =  ( pe0_act_instruction_counter ) == ( bv_6_11_n88 )  ;
assign bv_6_10_n90 = 6'ha ;
assign n91 =  ( pe0_act_instruction_counter ) == ( bv_6_10_n90 )  ;
assign bv_6_9_n92 = 6'h9 ;
assign n93 =  ( pe0_act_instruction_counter ) == ( bv_6_9_n92 )  ;
assign bv_6_8_n94 = 6'h8 ;
assign n95 =  ( pe0_act_instruction_counter ) == ( bv_6_8_n94 )  ;
assign bv_6_7_n96 = 6'h7 ;
assign n97 =  ( pe0_act_instruction_counter ) == ( bv_6_7_n96 )  ;
assign bv_6_6_n98 = 6'h6 ;
assign n99 =  ( pe0_act_instruction_counter ) == ( bv_6_6_n98 )  ;
assign bv_6_5_n100 = 6'h5 ;
assign n101 =  ( pe0_act_instruction_counter ) == ( bv_6_5_n100 )  ;
assign bv_6_4_n102 = 6'h4 ;
assign n103 =  ( pe0_act_instruction_counter ) == ( bv_6_4_n102 )  ;
assign bv_6_3_n104 = 6'h3 ;
assign n105 =  ( pe0_act_instruction_counter ) == ( bv_6_3_n104 )  ;
assign bv_6_2_n106 = 6'h2 ;
assign n107 =  ( pe0_act_instruction_counter ) == ( bv_6_2_n106 )  ;
assign bv_6_1_n108 = 6'h1 ;
assign n109 =  ( pe0_act_instruction_counter ) == ( bv_6_1_n108 )  ;
assign bv_6_0_n110 = 6'h0 ;
assign n111 =  ( pe0_act_instruction_counter ) == ( bv_6_0_n110 )  ;
assign n112 =  ( n111 ) ? ( act_vector_0_15_Inst_0 ) : ( act_vector_0_15_Inst_0 ) ;
assign n113 =  ( n109 ) ? ( act_vector_0_15_Inst_1 ) : ( n112 ) ;
assign n114 =  ( n107 ) ? ( act_vector_0_15_Inst_2 ) : ( n113 ) ;
assign n115 =  ( n105 ) ? ( act_vector_0_15_Inst_3 ) : ( n114 ) ;
assign n116 =  ( n103 ) ? ( act_vector_0_15_Inst_4 ) : ( n115 ) ;
assign n117 =  ( n101 ) ? ( act_vector_0_15_Inst_5 ) : ( n116 ) ;
assign n118 =  ( n99 ) ? ( act_vector_0_15_Inst_6 ) : ( n117 ) ;
assign n119 =  ( n97 ) ? ( act_vector_0_15_Inst_7 ) : ( n118 ) ;
assign n120 =  ( n95 ) ? ( act_vector_0_15_Inst_8 ) : ( n119 ) ;
assign n121 =  ( n93 ) ? ( act_vector_0_15_Inst_9 ) : ( n120 ) ;
assign n122 =  ( n91 ) ? ( act_vector_0_15_Inst_10 ) : ( n121 ) ;
assign n123 =  ( n89 ) ? ( act_vector_0_15_Inst_11 ) : ( n122 ) ;
assign n124 =  ( n87 ) ? ( act_vector_0_15_Inst_12 ) : ( n123 ) ;
assign n125 =  ( n85 ) ? ( act_vector_0_15_Inst_13 ) : ( n124 ) ;
assign n126 =  ( n83 ) ? ( act_vector_0_15_Inst_14 ) : ( n125 ) ;
assign n127 =  ( n81 ) ? ( act_vector_0_15_Inst_15 ) : ( n126 ) ;
assign n128 =  ( n79 ) ? ( act_vector_16_31_Inst_0 ) : ( n127 ) ;
assign n129 =  ( n77 ) ? ( act_vector_16_31_Inst_1 ) : ( n128 ) ;
assign n130 =  ( n75 ) ? ( act_vector_16_31_Inst_2 ) : ( n129 ) ;
assign n131 =  ( n73 ) ? ( act_vector_16_31_Inst_3 ) : ( n130 ) ;
assign n132 =  ( n71 ) ? ( act_vector_16_31_Inst_4 ) : ( n131 ) ;
assign n133 =  ( n69 ) ? ( act_vector_16_31_Inst_5 ) : ( n132 ) ;
assign n134 =  ( n67 ) ? ( act_vector_16_31_Inst_6 ) : ( n133 ) ;
assign n135 =  ( n65 ) ? ( act_vector_16_31_Inst_7 ) : ( n134 ) ;
assign n136 =  ( n63 ) ? ( act_vector_16_31_Inst_8 ) : ( n135 ) ;
assign n137 =  ( n61 ) ? ( act_vector_16_31_Inst_9 ) : ( n136 ) ;
assign n138 =  ( n59 ) ? ( act_vector_16_31_Inst_10 ) : ( n137 ) ;
assign n139 =  ( n57 ) ? ( act_vector_16_31_Inst_11 ) : ( n138 ) ;
assign n140 =  ( n55 ) ? ( act_vector_16_31_Inst_12 ) : ( n139 ) ;
assign n141 =  ( n53 ) ? ( act_vector_16_31_Inst_13 ) : ( n140 ) ;
assign n142 =  ( n51 ) ? ( act_vector_16_31_Inst_14 ) : ( n141 ) ;
assign n143 =  ( n49 ) ? ( act_vector_16_31_Inst_15 ) : ( n142 ) ;
assign n144 = n143[7:4] ;
assign bv_4_1_n145 = 4'h1 ;
assign n146 =  ( n144 ) == ( bv_4_1_n145 )  ;
assign n147 =  ( n47 ) & (n146 )  ;
assign n148 =  ( pe0_act_mngr_is_zero_first ) == ( bv_1_1_n0 )  ;
assign n149 =  ( n147 ) & (n148 )  ;
assign __ILA_pe_act_decode_of_PE0_act_child_op_load_zero__ = n149 ;
assign __ILA_pe_act_acc_decode__[5] = __ILA_pe_act_decode_of_PE0_act_child_op_load_zero__ ;
assign n150 =  ( pe0_act_is_start_reg ) == ( bv_1_1_n0 )  ;
assign n151 =  ( pe0_act_state ) == ( bv_2_1_n45 )  ;
assign n152 =  ( n150 ) & (n151 )  ;
assign n153 =  ( n144 ) == ( bv_4_1_n145 )  ;
assign n154 =  ( n152 ) & (n153 )  ;
assign n155 =  ( pe0_act_mngr_is_zero_first ) == ( bv_1_0_n32 )  ;
assign n156 =  ( n154 ) & (n155 )  ;
assign __ILA_pe_act_decode_of_PE0_act_child_op_load__ = n156 ;
assign __ILA_pe_act_acc_decode__[6] = __ILA_pe_act_decode_of_PE0_act_child_op_load__ ;
assign n157 =  ( pe0_act_is_start_reg ) == ( bv_1_1_n0 )  ;
assign n158 =  ( pe0_act_state ) == ( bv_2_1_n45 )  ;
assign n159 =  ( n157 ) & (n158 )  ;
assign bv_4_2_n160 = 4'h2 ;
assign n161 =  ( n144 ) == ( bv_4_2_n160 )  ;
assign n162 =  ( n159 ) & (n161 )  ;
assign __ILA_pe_act_decode_of_PE0_act_child_op_store__ = n162 ;
assign __ILA_pe_act_acc_decode__[7] = __ILA_pe_act_decode_of_PE0_act_child_op_store__ ;
assign n163 =  ( pe0_act_is_start_reg ) == ( bv_1_1_n0 )  ;
assign n164 =  ( pe0_act_state ) == ( bv_2_1_n45 )  ;
assign n165 =  ( n163 ) & (n164 )  ;
assign bv_4_3_n166 = 4'h3 ;
assign n167 =  ( n144 ) == ( bv_4_3_n166 )  ;
assign n168 =  ( n165 ) & (n167 )  ;
assign n169 =  ( pe0_act_reg_port_valid ) == ( bv_1_1_n0 )  ;
assign n170 =  ( act_port_ready ) == ( bv_1_1_n0 )  ;
assign n171 =  ( n169 ) & (n170 )  ;
assign n172 =  ( n168 ) & (n171 )  ;
assign __ILA_pe_act_decode_of_PE0_act_child_op_inpe__ = n172 ;
assign __ILA_pe_act_acc_decode__[8] = __ILA_pe_act_decode_of_PE0_act_child_op_inpe__ ;
assign n173 =  ( pe0_act_is_start_reg ) == ( bv_1_1_n0 )  ;
assign n174 =  ( pe0_act_state ) == ( bv_2_1_n45 )  ;
assign n175 =  ( n173 ) & (n174 )  ;
assign bv_4_4_n176 = 4'h4 ;
assign n177 =  ( n144 ) == ( bv_4_4_n176 )  ;
assign n178 =  ( n175 ) & (n177 )  ;
assign n179 =  ( output_port_valid ) == ( bv_1_0_n32 )  ;
assign n180 =  ( n178 ) & (n179 )  ;
assign __ILA_pe_act_decode_of_PE0_act_child_op_outgb__ = n180 ;
assign __ILA_pe_act_acc_decode__[9] = __ILA_pe_act_decode_of_PE0_act_child_op_outgb__ ;
assign n181 =  ( pe0_act_is_start_reg ) == ( bv_1_1_n0 )  ;
assign n182 =  ( pe0_act_state ) == ( bv_2_1_n45 )  ;
assign n183 =  ( n181 ) & (n182 )  ;
assign bv_4_7_n184 = 4'h7 ;
assign n185 =  ( n144 ) == ( bv_4_7_n184 )  ;
assign n186 =  ( n183 ) & (n185 )  ;
assign __ILA_pe_act_decode_of_PE0_act_child_op_copy__ = n186 ;
assign __ILA_pe_act_acc_decode__[10] = __ILA_pe_act_decode_of_PE0_act_child_op_copy__ ;
assign n187 =  ( pe0_act_is_start_reg ) == ( bv_1_1_n0 )  ;
assign n188 =  ( pe0_act_state ) == ( bv_2_1_n45 )  ;
assign n189 =  ( n187 ) & (n188 )  ;
assign bv_4_8_n190 = 4'h8 ;
assign n191 =  ( n144 ) == ( bv_4_8_n190 )  ;
assign n192 =  ( n189 ) & (n191 )  ;
assign __ILA_pe_act_decode_of_PE0_act_child_op_eadd__ = n192 ;
assign __ILA_pe_act_acc_decode__[11] = __ILA_pe_act_decode_of_PE0_act_child_op_eadd__ ;
assign n193 =  ( pe0_act_is_start_reg ) == ( bv_1_1_n0 )  ;
assign n194 =  ( pe0_act_state ) == ( bv_2_1_n45 )  ;
assign n195 =  ( n193 ) & (n194 )  ;
assign bv_4_9_n196 = 4'h9 ;
assign n197 =  ( n144 ) == ( bv_4_9_n196 )  ;
assign n198 =  ( n195 ) & (n197 )  ;
assign __ILA_pe_act_decode_of_PE0_act_child_op_emul__ = n198 ;
assign __ILA_pe_act_acc_decode__[12] = __ILA_pe_act_decode_of_PE0_act_child_op_emul__ ;
assign n199 =  ( pe0_act_is_start_reg ) == ( bv_1_1_n0 )  ;
assign n200 =  ( pe0_act_state ) == ( bv_2_1_n45 )  ;
assign n201 =  ( n199 ) & (n200 )  ;
assign bv_4_10_n202 = 4'ha ;
assign n203 =  ( n144 ) == ( bv_4_10_n202 )  ;
assign n204 =  ( n201 ) & (n203 )  ;
assign __ILA_pe_act_decode_of_PE0_act_child_op_sigm__ = n204 ;
assign __ILA_pe_act_acc_decode__[13] = __ILA_pe_act_decode_of_PE0_act_child_op_sigm__ ;
assign n205 =  ( pe0_act_is_start_reg ) == ( bv_1_1_n0 )  ;
assign n206 =  ( pe0_act_state ) == ( bv_2_1_n45 )  ;
assign n207 =  ( n205 ) & (n206 )  ;
assign bv_4_11_n208 = 4'hb ;
assign n209 =  ( n144 ) == ( bv_4_11_n208 )  ;
assign n210 =  ( n207 ) & (n209 )  ;
assign __ILA_pe_act_decode_of_PE0_act_child_op_tanh__ = n210 ;
assign __ILA_pe_act_acc_decode__[14] = __ILA_pe_act_decode_of_PE0_act_child_op_tanh__ ;
assign n211 =  ( pe0_act_is_start_reg ) == ( bv_1_1_n0 )  ;
assign n212 =  ( pe0_act_state ) == ( bv_2_1_n45 )  ;
assign n213 =  ( n211 ) & (n212 )  ;
assign bv_4_12_n214 = 4'hc ;
assign n215 =  ( n144 ) == ( bv_4_12_n214 )  ;
assign n216 =  ( n213 ) & (n215 )  ;
assign __ILA_pe_act_decode_of_PE0_act_child_op_relu__ = n216 ;
assign __ILA_pe_act_acc_decode__[15] = __ILA_pe_act_decode_of_PE0_act_child_op_relu__ ;
assign n217 =  ( pe0_act_is_start_reg ) == ( bv_1_1_n0 )  ;
assign n218 =  ( pe0_act_state ) == ( bv_2_1_n45 )  ;
assign n219 =  ( n217 ) & (n218 )  ;
assign bv_4_13_n220 = 4'hd ;
assign n221 =  ( n144 ) == ( bv_4_13_n220 )  ;
assign n222 =  ( n219 ) & (n221 )  ;
assign __ILA_pe_act_decode_of_PE0_act_child_op_onex__ = n222 ;
assign __ILA_pe_act_acc_decode__[16] = __ILA_pe_act_decode_of_PE0_act_child_op_onex__ ;
assign n223 =  ( pe0_act_is_start_reg ) == ( bv_1_1_n0 )  ;
assign bv_2_2_n224 = 2'h2 ;
assign n225 =  ( pe0_act_state ) == ( bv_2_2_n224 )  ;
assign n226 =  ( output_port_valid ) == ( bv_1_0_n32 )  ;
assign n227 =  ( n225 ) & (n226 )  ;
assign n228 =  ( done_valid ) == ( bv_1_0_n32 )  ;
assign n229 =  ( n227 ) & (n228 )  ;
assign n230 =  ( n223 ) & (n229 )  ;
assign __ILA_pe_act_decode_of_PE0_act_child_reg_store__ = n230 ;
assign __ILA_pe_act_acc_decode__[17] = __ILA_pe_act_decode_of_PE0_act_child_reg_store__ ;
assign n231 =  ( pe0_act_is_start_reg ) == ( bv_1_1_n0 )  ;
assign n232 =  ( pe0_act_state ) == ( bv_2_2_n224 )  ;
assign n233 =  ( output_port_valid ) == ( bv_1_1_n0 )  ;
assign n234 =  ( output_port_ready ) == ( bv_1_1_n0 )  ;
assign n235 =  ( n233 ) & (n234 )  ;
assign n236 =  ( n232 ) & (n235 )  ;
assign n237 =  ( n231 ) & (n236 )  ;
assign __ILA_pe_act_decode_of_PE0_act_child_out_sent__ = n237 ;
assign __ILA_pe_act_acc_decode__[18] = __ILA_pe_act_decode_of_PE0_act_child_out_sent__ ;
assign n238 =  ( pe0_act_is_start_reg ) == ( bv_1_1_n0 )  ;
assign n239 =  ( pe0_act_state ) == ( bv_2_2_n224 )  ;
assign n240 =  ( done_valid ) == ( bv_1_1_n0 )  ;
assign n241 =  ( done_ready ) == ( bv_1_1_n0 )  ;
assign n242 =  ( n240 ) & (n241 )  ;
assign n243 =  ( n239 ) & (n242 )  ;
assign n244 =  ( n238 ) & (n243 )  ;
assign __ILA_pe_act_decode_of_PE0_act_child_done_sent__ = n244 ;
assign __ILA_pe_act_acc_decode__[19] = __ILA_pe_act_decode_of_PE0_act_child_done_sent__ ;
assign n245 =  ( pe0_act_output_counter ) + ( pe0_act_mngr_output_addr_base )  ;
assign n246 =  ( pe0_act_mngr_num_inst ) - ( bv_6_1_n108 )  ;
assign n247 =  ( pe0_act_instruction_counter ) == ( n246 )  ;
assign bv_8_1_n248 = 8'h1 ;
assign n249 =  ( pe0_act_mngr_num_output ) - ( bv_8_1_n248 )  ;
assign n250 =  ( pe0_act_output_counter ) == ( n249 )  ;
assign n251 =  ( n247 ) & (n250 )  ;
assign n252 =  ( n251 ) ? ( bv_1_1_n0 ) : ( done ) ;
assign n253 =  ( pe0_act_mngr_num_inst ) - ( bv_6_1_n108 )  ;
assign n254 =  ( pe0_act_instruction_counter ) == ( n253 )  ;
assign n255 =  ( pe0_act_mngr_num_output ) - ( bv_8_1_n248 )  ;
assign n256 =  ( pe0_act_output_counter ) == ( n255 )  ;
assign n257 =  ( n254 ) & (n256 )  ;
assign n258 =  ( n257 ) ? ( bv_1_1_n0 ) : ( done ) ;
assign n259 =  ( pe0_act_mngr_num_inst ) - ( bv_6_1_n108 )  ;
assign n260 =  ( pe0_act_instruction_counter ) == ( n259 )  ;
assign n261 =  ( pe0_act_mngr_num_output ) - ( bv_8_1_n248 )  ;
assign n262 =  ( pe0_act_output_counter ) == ( n261 )  ;
assign n263 =  ( n260 ) & (n262 )  ;
assign n264 =  ( n263 ) ? ( bv_1_1_n0 ) : ( done ) ;
assign n265 =  ( pe0_act_mngr_num_inst ) - ( bv_6_1_n108 )  ;
assign n266 =  ( pe0_act_instruction_counter ) == ( n265 )  ;
assign n267 =  ( pe0_act_mngr_num_output ) - ( bv_8_1_n248 )  ;
assign n268 =  ( pe0_act_output_counter ) == ( n267 )  ;
assign n269 =  ( n266 ) & (n268 )  ;
assign n270 =  ( n269 ) ? ( bv_1_1_n0 ) : ( done ) ;
assign n271 =  ( pe0_act_mngr_num_inst ) - ( bv_6_1_n108 )  ;
assign n272 =  ( pe0_act_instruction_counter ) == ( n271 )  ;
assign n273 =  ( pe0_act_mngr_num_output ) - ( bv_8_1_n248 )  ;
assign n274 =  ( pe0_act_output_counter ) == ( n273 )  ;
assign n275 =  ( n272 ) & (n274 )  ;
assign n276 =  ( n275 ) ? ( bv_1_1_n0 ) : ( done ) ;
assign n277 =  ( pe0_act_mngr_num_inst ) - ( bv_6_1_n108 )  ;
assign n278 =  ( pe0_act_instruction_counter ) == ( n277 )  ;
assign n279 =  ( pe0_act_mngr_num_output ) - ( bv_8_1_n248 )  ;
assign n280 =  ( pe0_act_output_counter ) == ( n279 )  ;
assign n281 =  ( n278 ) & (n280 )  ;
assign n282 =  ( n281 ) ? ( bv_1_1_n0 ) : ( done ) ;
assign n283 =  ( pe0_act_mngr_num_inst ) - ( bv_6_1_n108 )  ;
assign n284 =  ( pe0_act_instruction_counter ) == ( n283 )  ;
assign n285 =  ( pe0_act_mngr_num_output ) - ( bv_8_1_n248 )  ;
assign n286 =  ( pe0_act_output_counter ) == ( n285 )  ;
assign n287 =  ( n284 ) & (n286 )  ;
assign n288 =  ( n287 ) ? ( bv_1_1_n0 ) : ( done ) ;
assign n289 =  ( pe0_act_mngr_num_inst ) - ( bv_6_1_n108 )  ;
assign n290 =  ( pe0_act_instruction_counter ) == ( n289 )  ;
assign n291 =  ( pe0_act_mngr_num_output ) - ( bv_8_1_n248 )  ;
assign n292 =  ( pe0_act_output_counter ) == ( n291 )  ;
assign n293 =  ( n290 ) & (n292 )  ;
assign n294 =  ( n293 ) ? ( bv_1_1_n0 ) : ( done ) ;
assign n295 =  ( pe0_act_mngr_num_inst ) - ( bv_6_1_n108 )  ;
assign n296 =  ( pe0_act_instruction_counter ) == ( n295 )  ;
assign n297 =  ( pe0_act_mngr_num_output ) - ( bv_8_1_n248 )  ;
assign n298 =  ( pe0_act_output_counter ) == ( n297 )  ;
assign n299 =  ( n296 ) & (n298 )  ;
assign n300 =  ( n299 ) ? ( bv_1_1_n0 ) : ( done ) ;
assign n301 =  ( pe0_act_mngr_num_inst ) - ( bv_6_1_n108 )  ;
assign n302 =  ( pe0_act_instruction_counter ) == ( n301 )  ;
assign n303 =  ( pe0_act_mngr_num_output ) - ( bv_8_1_n248 )  ;
assign n304 =  ( pe0_act_output_counter ) == ( n303 )  ;
assign n305 =  ( n302 ) & (n304 )  ;
assign n306 =  ( n305 ) ? ( bv_1_1_n0 ) : ( done ) ;
assign n307 =  ( pe0_act_mngr_num_inst ) - ( bv_6_1_n108 )  ;
assign n308 =  ( pe0_act_instruction_counter ) == ( n307 )  ;
assign n309 =  ( pe0_act_mngr_num_output ) - ( bv_8_1_n248 )  ;
assign n310 =  ( pe0_act_output_counter ) == ( n309 )  ;
assign n311 =  ( n308 ) & (n310 )  ;
assign n312 =  ( n311 ) ? ( bv_1_1_n0 ) : ( done ) ;
assign n313 =  ( pe0_act_mngr_num_inst ) - ( bv_6_1_n108 )  ;
assign n314 =  ( pe0_act_instruction_counter ) == ( n313 )  ;
assign n315 =  ( pe0_act_mngr_num_output ) - ( bv_8_1_n248 )  ;
assign n316 =  ( pe0_act_output_counter ) == ( n315 )  ;
assign n317 =  ( n314 ) & (n316 )  ;
assign n318 =  ( n317 ) ? ( bv_1_1_n0 ) : ( done ) ;
assign n319 =  ( n251 ) ? ( bv_1_1_n0 ) : ( bv_1_0_n32 ) ;
assign n320 =  ( n257 ) ? ( bv_1_1_n0 ) : ( bv_1_0_n32 ) ;
assign n321 =  ( n263 ) ? ( bv_1_1_n0 ) : ( bv_1_0_n32 ) ;
assign n322 =  ( n269 ) ? ( bv_1_1_n0 ) : ( bv_1_0_n32 ) ;
assign n323 =  ( n275 ) ? ( bv_1_1_n0 ) : ( bv_1_0_n32 ) ;
assign n324 =  ( n281 ) ? ( bv_1_1_n0 ) : ( bv_1_0_n32 ) ;
assign n325 =  ( n287 ) ? ( bv_1_1_n0 ) : ( bv_1_0_n32 ) ;
assign n326 =  ( n293 ) ? ( bv_1_1_n0 ) : ( bv_1_0_n32 ) ;
assign n327 =  ( n299 ) ? ( bv_1_1_n0 ) : ( bv_1_0_n32 ) ;
assign n328 =  ( n305 ) ? ( bv_1_1_n0 ) : ( bv_1_0_n32 ) ;
assign n329 =  ( n311 ) ? ( bv_1_1_n0 ) : ( bv_1_0_n32 ) ;
assign n330 =  ( n317 ) ? ( bv_1_1_n0 ) : ( bv_1_0_n32 ) ;
assign n331 = data_in_0[0:0] ;
assign n332 = data_in_1[0:0] ;
assign n333 =  ( n251 ) ? ( bv_1_0_n32 ) : ( pe0_act_mngr_is_zero_first ) ;
assign n334 =  ( n257 ) ? ( bv_1_0_n32 ) : ( pe0_act_mngr_is_zero_first ) ;
assign n335 =  ( n263 ) ? ( bv_1_0_n32 ) : ( pe0_act_mngr_is_zero_first ) ;
assign n336 =  ( n269 ) ? ( bv_1_0_n32 ) : ( pe0_act_mngr_is_zero_first ) ;
assign n337 =  ( n275 ) ? ( bv_1_0_n32 ) : ( pe0_act_mngr_is_zero_first ) ;
assign n338 =  ( n281 ) ? ( bv_1_0_n32 ) : ( pe0_act_mngr_is_zero_first ) ;
assign n339 =  ( n287 ) ? ( bv_1_0_n32 ) : ( pe0_act_mngr_is_zero_first ) ;
assign n340 =  ( n293 ) ? ( bv_1_0_n32 ) : ( pe0_act_mngr_is_zero_first ) ;
assign n341 =  ( n299 ) ? ( bv_1_0_n32 ) : ( pe0_act_mngr_is_zero_first ) ;
assign n342 =  ( n305 ) ? ( bv_1_0_n32 ) : ( pe0_act_mngr_is_zero_first ) ;
assign n343 =  ( n311 ) ? ( bv_1_0_n32 ) : ( pe0_act_mngr_is_zero_first ) ;
assign n344 =  ( n317 ) ? ( bv_1_0_n32 ) : ( pe0_act_mngr_is_zero_first ) ;
assign n345 = data_in_2[2:0] ;
assign n346 = data_in_3[5:0] ;
assign n347 =  { ( data_in_7 ) , ( data_in_6 ) }  ;
assign n348 = n347[4:0] ;
assign n349 = ~ ( n162 )  ;
assign n350 =  ( 1'b1 ) & (n349 )  ;
assign n351 = ~ ( n30 )  ;
assign n352 =  ( n350 ) & (n351 )  ;
assign n353 =  ( n350 ) & (n30 )  ;
assign bv_8_0_n354 = 8'h0 ;
assign n355 =  { ( bv_8_0_n354 ) , ( addr ) }  ;
assign bv_32_9437184_n356 = 32'h900000 ;
assign n357 =  ( n355 ) - ( bv_32_9437184_n356 )  ;
assign bv_32_15_n358 = 32'hf ;
assign n359 =  ( n357 ) + ( bv_32_15_n358 )  ;
assign bv_32_14_n360 = 32'he ;
assign n361 =  ( n357 ) + ( bv_32_14_n360 )  ;
assign bv_32_13_n362 = 32'hd ;
assign n363 =  ( n357 ) + ( bv_32_13_n362 )  ;
assign bv_32_12_n364 = 32'hc ;
assign n365 =  ( n357 ) + ( bv_32_12_n364 )  ;
assign bv_32_11_n366 = 32'hb ;
assign n367 =  ( n357 ) + ( bv_32_11_n366 )  ;
assign bv_32_10_n368 = 32'ha ;
assign n369 =  ( n357 ) + ( bv_32_10_n368 )  ;
assign bv_32_9_n370 = 32'h9 ;
assign n371 =  ( n357 ) + ( bv_32_9_n370 )  ;
assign bv_32_8_n372 = 32'h8 ;
assign n373 =  ( n357 ) + ( bv_32_8_n372 )  ;
assign bv_32_7_n374 = 32'h7 ;
assign n375 =  ( n357 ) + ( bv_32_7_n374 )  ;
assign bv_32_6_n376 = 32'h6 ;
assign n377 =  ( n357 ) + ( bv_32_6_n376 )  ;
assign bv_32_5_n378 = 32'h5 ;
assign n379 =  ( n357 ) + ( bv_32_5_n378 )  ;
assign bv_32_4_n380 = 32'h4 ;
assign n381 =  ( n357 ) + ( bv_32_4_n380 )  ;
assign bv_32_3_n382 = 32'h3 ;
assign n383 =  ( n357 ) + ( bv_32_3_n382 )  ;
assign bv_32_2_n384 = 32'h2 ;
assign n385 =  ( n357 ) + ( bv_32_2_n384 )  ;
assign bv_32_1_n386 = 32'h1 ;
assign n387 =  ( n357 ) + ( bv_32_1_n386 )  ;
assign bv_32_0_n388 = 32'h0 ;
assign n389 =  ( n357 ) + ( bv_32_0_n388 )  ;
assign n390 =  ( 1'b1 ) & (n162 )  ;
assign bv_24_0_n391 = 24'h0 ;
assign n392 =  { ( bv_24_0_n391 ) , ( pe0_act_output_counter ) }  ;
assign bv_27_0_n393 = 27'h0 ;
assign n394 =  { ( bv_27_0_n393 ) , ( pe0_act_mngr_buffer_addr_base ) }  ;
assign n395 =  ( n392 ) + ( n394 )  ;
assign n396 =  ( n395 ) << ( bv_32_4_n380 )  ;
assign n397 =  ( n396 ) + ( bv_32_15_n358 )  ;
assign n398 = n143[3:2] ;
assign bv_2_3_n399 = 2'h3 ;
assign n400 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign bv_4_15_n401 = 4'hf ;
assign bv_4_0_n402 = 4'h0 ;
assign n403 =  ( bv_4_15_n401 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n404 = n403 ;
assign n406 = PE0_act_regs_3_data_n405 ;
assign n407 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n408 = n403 ;
assign n410 = PE0_act_regs_2_data_n409 ;
assign n411 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n412 = n403 ;
assign n414 = PE0_act_regs_1_data_n413 ;
assign n415 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n416 = n403 ;
assign n418 = PE0_act_regs_0_data_n417 ;
assign bv_20_0_n419 = 20'h0 ;
assign n420 =  ( n415 ) ? ( n418 ) : ( bv_20_0_n419 ) ;
assign n421 =  ( n411 ) ? ( n414 ) : ( n420 ) ;
assign n422 =  ( n407 ) ? ( n410 ) : ( n421 ) ;
assign n423 =  ( n400 ) ? ( n406 ) : ( n422 ) ;
fun_Fixed2Adaptfloat  applyFunc_n425(
    .arg0( n423 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n424 )
);
assign n426 = n424 ;
assign n427 =  ( n396 ) + ( bv_32_14_n360 )  ;
assign n428 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign bv_4_14_n429 = 4'he ;
assign n430 =  ( bv_4_14_n429 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n431 = n430 ;
assign n433 = PE0_act_regs_3_data_n432 ;
assign n434 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n435 = n430 ;
assign n437 = PE0_act_regs_2_data_n436 ;
assign n438 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n439 = n430 ;
assign n441 = PE0_act_regs_1_data_n440 ;
assign n442 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n443 = n430 ;
assign n445 = PE0_act_regs_0_data_n444 ;
assign n446 =  ( n442 ) ? ( n445 ) : ( bv_20_0_n419 ) ;
assign n447 =  ( n438 ) ? ( n441 ) : ( n446 ) ;
assign n448 =  ( n434 ) ? ( n437 ) : ( n447 ) ;
assign n449 =  ( n428 ) ? ( n433 ) : ( n448 ) ;
fun_Fixed2Adaptfloat  applyFunc_n451(
    .arg0( n449 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n450 )
);
assign n452 = n450 ;
assign n453 =  ( n396 ) + ( bv_32_13_n362 )  ;
assign n454 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n455 =  ( bv_4_13_n220 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n456 = n455 ;
assign n458 = PE0_act_regs_3_data_n457 ;
assign n459 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n460 = n455 ;
assign n462 = PE0_act_regs_2_data_n461 ;
assign n463 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n464 = n455 ;
assign n466 = PE0_act_regs_1_data_n465 ;
assign n467 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n468 = n455 ;
assign n470 = PE0_act_regs_0_data_n469 ;
assign n471 =  ( n467 ) ? ( n470 ) : ( bv_20_0_n419 ) ;
assign n472 =  ( n463 ) ? ( n466 ) : ( n471 ) ;
assign n473 =  ( n459 ) ? ( n462 ) : ( n472 ) ;
assign n474 =  ( n454 ) ? ( n458 ) : ( n473 ) ;
fun_Fixed2Adaptfloat  applyFunc_n476(
    .arg0( n474 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n475 )
);
assign n477 = n475 ;
assign n478 =  ( n396 ) + ( bv_32_12_n364 )  ;
assign n479 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n480 =  ( bv_4_12_n214 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n481 = n480 ;
assign n483 = PE0_act_regs_3_data_n482 ;
assign n484 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n485 = n480 ;
assign n487 = PE0_act_regs_2_data_n486 ;
assign n488 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n489 = n480 ;
assign n491 = PE0_act_regs_1_data_n490 ;
assign n492 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n493 = n480 ;
assign n495 = PE0_act_regs_0_data_n494 ;
assign n496 =  ( n492 ) ? ( n495 ) : ( bv_20_0_n419 ) ;
assign n497 =  ( n488 ) ? ( n491 ) : ( n496 ) ;
assign n498 =  ( n484 ) ? ( n487 ) : ( n497 ) ;
assign n499 =  ( n479 ) ? ( n483 ) : ( n498 ) ;
fun_Fixed2Adaptfloat  applyFunc_n501(
    .arg0( n499 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n500 )
);
assign n502 = n500 ;
assign n503 =  ( n396 ) + ( bv_32_11_n366 )  ;
assign n504 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n505 =  ( bv_4_11_n208 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n506 = n505 ;
assign n508 = PE0_act_regs_3_data_n507 ;
assign n509 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n510 = n505 ;
assign n512 = PE0_act_regs_2_data_n511 ;
assign n513 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n514 = n505 ;
assign n516 = PE0_act_regs_1_data_n515 ;
assign n517 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n518 = n505 ;
assign n520 = PE0_act_regs_0_data_n519 ;
assign n521 =  ( n517 ) ? ( n520 ) : ( bv_20_0_n419 ) ;
assign n522 =  ( n513 ) ? ( n516 ) : ( n521 ) ;
assign n523 =  ( n509 ) ? ( n512 ) : ( n522 ) ;
assign n524 =  ( n504 ) ? ( n508 ) : ( n523 ) ;
fun_Fixed2Adaptfloat  applyFunc_n526(
    .arg0( n524 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n525 )
);
assign n527 = n525 ;
assign n528 =  ( n396 ) + ( bv_32_10_n368 )  ;
assign n529 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n530 =  ( bv_4_10_n202 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n531 = n530 ;
assign n533 = PE0_act_regs_3_data_n532 ;
assign n534 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n535 = n530 ;
assign n537 = PE0_act_regs_2_data_n536 ;
assign n538 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n539 = n530 ;
assign n541 = PE0_act_regs_1_data_n540 ;
assign n542 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n543 = n530 ;
assign n545 = PE0_act_regs_0_data_n544 ;
assign n546 =  ( n542 ) ? ( n545 ) : ( bv_20_0_n419 ) ;
assign n547 =  ( n538 ) ? ( n541 ) : ( n546 ) ;
assign n548 =  ( n534 ) ? ( n537 ) : ( n547 ) ;
assign n549 =  ( n529 ) ? ( n533 ) : ( n548 ) ;
fun_Fixed2Adaptfloat  applyFunc_n551(
    .arg0( n549 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n550 )
);
assign n552 = n550 ;
assign n553 =  ( n396 ) + ( bv_32_9_n370 )  ;
assign n554 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n555 =  ( bv_4_9_n196 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n556 = n555 ;
assign n558 = PE0_act_regs_3_data_n557 ;
assign n559 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n560 = n555 ;
assign n562 = PE0_act_regs_2_data_n561 ;
assign n563 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n564 = n555 ;
assign n566 = PE0_act_regs_1_data_n565 ;
assign n567 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n568 = n555 ;
assign n570 = PE0_act_regs_0_data_n569 ;
assign n571 =  ( n567 ) ? ( n570 ) : ( bv_20_0_n419 ) ;
assign n572 =  ( n563 ) ? ( n566 ) : ( n571 ) ;
assign n573 =  ( n559 ) ? ( n562 ) : ( n572 ) ;
assign n574 =  ( n554 ) ? ( n558 ) : ( n573 ) ;
fun_Fixed2Adaptfloat  applyFunc_n576(
    .arg0( n574 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n575 )
);
assign n577 = n575 ;
assign n578 =  ( n396 ) + ( bv_32_8_n372 )  ;
assign n579 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n580 =  ( bv_4_8_n190 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n581 = n580 ;
assign n583 = PE0_act_regs_3_data_n582 ;
assign n584 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n585 = n580 ;
assign n587 = PE0_act_regs_2_data_n586 ;
assign n588 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n589 = n580 ;
assign n591 = PE0_act_regs_1_data_n590 ;
assign n592 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n593 = n580 ;
assign n595 = PE0_act_regs_0_data_n594 ;
assign n596 =  ( n592 ) ? ( n595 ) : ( bv_20_0_n419 ) ;
assign n597 =  ( n588 ) ? ( n591 ) : ( n596 ) ;
assign n598 =  ( n584 ) ? ( n587 ) : ( n597 ) ;
assign n599 =  ( n579 ) ? ( n583 ) : ( n598 ) ;
fun_Fixed2Adaptfloat  applyFunc_n601(
    .arg0( n599 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n600 )
);
assign n602 = n600 ;
assign n603 =  ( n396 ) + ( bv_32_7_n374 )  ;
assign n604 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n605 =  ( bv_4_7_n184 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n606 = n605 ;
assign n608 = PE0_act_regs_3_data_n607 ;
assign n609 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n610 = n605 ;
assign n612 = PE0_act_regs_2_data_n611 ;
assign n613 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n614 = n605 ;
assign n616 = PE0_act_regs_1_data_n615 ;
assign n617 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n618 = n605 ;
assign n620 = PE0_act_regs_0_data_n619 ;
assign n621 =  ( n617 ) ? ( n620 ) : ( bv_20_0_n419 ) ;
assign n622 =  ( n613 ) ? ( n616 ) : ( n621 ) ;
assign n623 =  ( n609 ) ? ( n612 ) : ( n622 ) ;
assign n624 =  ( n604 ) ? ( n608 ) : ( n623 ) ;
fun_Fixed2Adaptfloat  applyFunc_n626(
    .arg0( n624 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n625 )
);
assign n627 = n625 ;
assign n628 =  ( n396 ) + ( bv_32_6_n376 )  ;
assign n629 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign bv_4_6_n630 = 4'h6 ;
assign n631 =  ( bv_4_6_n630 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n632 = n631 ;
assign n634 = PE0_act_regs_3_data_n633 ;
assign n635 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n636 = n631 ;
assign n638 = PE0_act_regs_2_data_n637 ;
assign n639 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n640 = n631 ;
assign n642 = PE0_act_regs_1_data_n641 ;
assign n643 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n644 = n631 ;
assign n646 = PE0_act_regs_0_data_n645 ;
assign n647 =  ( n643 ) ? ( n646 ) : ( bv_20_0_n419 ) ;
assign n648 =  ( n639 ) ? ( n642 ) : ( n647 ) ;
assign n649 =  ( n635 ) ? ( n638 ) : ( n648 ) ;
assign n650 =  ( n629 ) ? ( n634 ) : ( n649 ) ;
fun_Fixed2Adaptfloat  applyFunc_n652(
    .arg0( n650 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n651 )
);
assign n653 = n651 ;
assign n654 =  ( n396 ) + ( bv_32_5_n378 )  ;
assign n655 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign bv_4_5_n656 = 4'h5 ;
assign n657 =  ( bv_4_5_n656 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n658 = n657 ;
assign n660 = PE0_act_regs_3_data_n659 ;
assign n661 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n662 = n657 ;
assign n664 = PE0_act_regs_2_data_n663 ;
assign n665 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n666 = n657 ;
assign n668 = PE0_act_regs_1_data_n667 ;
assign n669 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n670 = n657 ;
assign n672 = PE0_act_regs_0_data_n671 ;
assign n673 =  ( n669 ) ? ( n672 ) : ( bv_20_0_n419 ) ;
assign n674 =  ( n665 ) ? ( n668 ) : ( n673 ) ;
assign n675 =  ( n661 ) ? ( n664 ) : ( n674 ) ;
assign n676 =  ( n655 ) ? ( n660 ) : ( n675 ) ;
fun_Fixed2Adaptfloat  applyFunc_n678(
    .arg0( n676 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n677 )
);
assign n679 = n677 ;
assign n680 =  ( n396 ) + ( bv_32_4_n380 )  ;
assign n681 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n682 =  ( bv_4_4_n176 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n683 = n682 ;
assign n685 = PE0_act_regs_3_data_n684 ;
assign n686 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n687 = n682 ;
assign n689 = PE0_act_regs_2_data_n688 ;
assign n690 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n691 = n682 ;
assign n693 = PE0_act_regs_1_data_n692 ;
assign n694 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n695 = n682 ;
assign n697 = PE0_act_regs_0_data_n696 ;
assign n698 =  ( n694 ) ? ( n697 ) : ( bv_20_0_n419 ) ;
assign n699 =  ( n690 ) ? ( n693 ) : ( n698 ) ;
assign n700 =  ( n686 ) ? ( n689 ) : ( n699 ) ;
assign n701 =  ( n681 ) ? ( n685 ) : ( n700 ) ;
fun_Fixed2Adaptfloat  applyFunc_n703(
    .arg0( n701 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n702 )
);
assign n704 = n702 ;
assign n705 =  ( n396 ) + ( bv_32_3_n382 )  ;
assign n706 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n707 =  ( bv_4_3_n166 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n708 = n707 ;
assign n710 = PE0_act_regs_3_data_n709 ;
assign n711 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n712 = n707 ;
assign n714 = PE0_act_regs_2_data_n713 ;
assign n715 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n716 = n707 ;
assign n718 = PE0_act_regs_1_data_n717 ;
assign n719 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n720 = n707 ;
assign n722 = PE0_act_regs_0_data_n721 ;
assign n723 =  ( n719 ) ? ( n722 ) : ( bv_20_0_n419 ) ;
assign n724 =  ( n715 ) ? ( n718 ) : ( n723 ) ;
assign n725 =  ( n711 ) ? ( n714 ) : ( n724 ) ;
assign n726 =  ( n706 ) ? ( n710 ) : ( n725 ) ;
fun_Fixed2Adaptfloat  applyFunc_n728(
    .arg0( n726 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n727 )
);
assign n729 = n727 ;
assign n730 =  ( n396 ) + ( bv_32_2_n384 )  ;
assign n731 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n732 =  ( bv_4_2_n160 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n733 = n732 ;
assign n735 = PE0_act_regs_3_data_n734 ;
assign n736 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n737 = n732 ;
assign n739 = PE0_act_regs_2_data_n738 ;
assign n740 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n741 = n732 ;
assign n743 = PE0_act_regs_1_data_n742 ;
assign n744 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n745 = n732 ;
assign n747 = PE0_act_regs_0_data_n746 ;
assign n748 =  ( n744 ) ? ( n747 ) : ( bv_20_0_n419 ) ;
assign n749 =  ( n740 ) ? ( n743 ) : ( n748 ) ;
assign n750 =  ( n736 ) ? ( n739 ) : ( n749 ) ;
assign n751 =  ( n731 ) ? ( n735 ) : ( n750 ) ;
fun_Fixed2Adaptfloat  applyFunc_n753(
    .arg0( n751 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n752 )
);
assign n754 = n752 ;
assign n755 =  ( n396 ) + ( bv_32_1_n386 )  ;
assign n756 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n757 =  ( bv_4_1_n145 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n758 = n757 ;
assign n760 = PE0_act_regs_3_data_n759 ;
assign n761 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n762 = n757 ;
assign n764 = PE0_act_regs_2_data_n763 ;
assign n765 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n766 = n757 ;
assign n768 = PE0_act_regs_1_data_n767 ;
assign n769 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n770 = n757 ;
assign n772 = PE0_act_regs_0_data_n771 ;
assign n773 =  ( n769 ) ? ( n772 ) : ( bv_20_0_n419 ) ;
assign n774 =  ( n765 ) ? ( n768 ) : ( n773 ) ;
assign n775 =  ( n761 ) ? ( n764 ) : ( n774 ) ;
assign n776 =  ( n756 ) ? ( n760 ) : ( n775 ) ;
fun_Fixed2Adaptfloat  applyFunc_n778(
    .arg0( n776 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n777 )
);
assign n779 = n777 ;
assign n780 =  ( n396 ) + ( bv_32_0_n388 )  ;
assign n781 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n782 =  ( bv_4_0_n402 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n783 = n782 ;
assign n785 = PE0_act_regs_3_data_n784 ;
assign n786 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n787 = n782 ;
assign n789 = PE0_act_regs_2_data_n788 ;
assign n790 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n791 = n782 ;
assign n793 = PE0_act_regs_1_data_n792 ;
assign n794 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n795 = n782 ;
assign n797 = PE0_act_regs_0_data_n796 ;
assign n798 =  ( n794 ) ? ( n797 ) : ( bv_20_0_n419 ) ;
assign n799 =  ( n790 ) ? ( n793 ) : ( n798 ) ;
assign n800 =  ( n786 ) ? ( n789 ) : ( n799 ) ;
assign n801 =  ( n781 ) ? ( n785 ) : ( n800 ) ;
fun_Fixed2Adaptfloat  applyFunc_n803(
    .arg0( n801 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n802 )
);
assign n804 = n802 ;
assign pe0_act_buffer_addr0 = n390 ? (n397) : (n353 ? (n359) : (0)) ;
assign pe0_act_buffer_data0 = n390 ? (n426) : (n353 ? (data_in_15) : ('d0)) ;
assign pe0_act_buffer_wen0 = (n390) ? ( 1'b1 ) : ((n353) ? ( 1'b1 ) : (1'b0)) ;
assign pe0_act_buffer_addr1 = n390 ? (n427) : (n353 ? (n361) : (0)) ;
assign pe0_act_buffer_data1 = n390 ? (n452) : (n353 ? (data_in_14) : ('d0)) ;
assign pe0_act_buffer_wen1 = (n390) ? ( 1'b1 ) : ((n353) ? ( 1'b1 ) : (1'b0)) ;
assign pe0_act_buffer_addr2 = n390 ? (n453) : (n353 ? (n363) : (0)) ;
assign pe0_act_buffer_data2 = n390 ? (n477) : (n353 ? (data_in_13) : ('d0)) ;
assign pe0_act_buffer_wen2 = (n390) ? ( 1'b1 ) : ((n353) ? ( 1'b1 ) : (1'b0)) ;
assign pe0_act_buffer_addr3 = n390 ? (n478) : (n353 ? (n365) : (0)) ;
assign pe0_act_buffer_data3 = n390 ? (n502) : (n353 ? (data_in_12) : ('d0)) ;
assign pe0_act_buffer_wen3 = (n390) ? ( 1'b1 ) : ((n353) ? ( 1'b1 ) : (1'b0)) ;
assign pe0_act_buffer_addr4 = n390 ? (n503) : (n353 ? (n367) : (0)) ;
assign pe0_act_buffer_data4 = n390 ? (n527) : (n353 ? (data_in_11) : ('d0)) ;
assign pe0_act_buffer_wen4 = (n390) ? ( 1'b1 ) : ((n353) ? ( 1'b1 ) : (1'b0)) ;
assign pe0_act_buffer_addr5 = n390 ? (n528) : (n353 ? (n369) : (0)) ;
assign pe0_act_buffer_data5 = n390 ? (n552) : (n353 ? (data_in_10) : ('d0)) ;
assign pe0_act_buffer_wen5 = (n390) ? ( 1'b1 ) : ((n353) ? ( 1'b1 ) : (1'b0)) ;
assign pe0_act_buffer_addr6 = n390 ? (n553) : (n353 ? (n371) : (0)) ;
assign pe0_act_buffer_data6 = n390 ? (n577) : (n353 ? (data_in_9) : ('d0)) ;
assign pe0_act_buffer_wen6 = (n390) ? ( 1'b1 ) : ((n353) ? ( 1'b1 ) : (1'b0)) ;
assign pe0_act_buffer_addr7 = n390 ? (n578) : (n353 ? (n373) : (0)) ;
assign pe0_act_buffer_data7 = n390 ? (n602) : (n353 ? (data_in_8) : ('d0)) ;
assign pe0_act_buffer_wen7 = (n390) ? ( 1'b1 ) : ((n353) ? ( 1'b1 ) : (1'b0)) ;
assign pe0_act_buffer_addr8 = n390 ? (n603) : (n353 ? (n375) : (0)) ;
assign pe0_act_buffer_data8 = n390 ? (n627) : (n353 ? (data_in_7) : ('d0)) ;
assign pe0_act_buffer_wen8 = (n390) ? ( 1'b1 ) : ((n353) ? ( 1'b1 ) : (1'b0)) ;
assign pe0_act_buffer_addr9 = n390 ? (n628) : (n353 ? (n377) : (0)) ;
assign pe0_act_buffer_data9 = n390 ? (n653) : (n353 ? (data_in_6) : ('d0)) ;
assign pe0_act_buffer_wen9 = (n390) ? ( 1'b1 ) : ((n353) ? ( 1'b1 ) : (1'b0)) ;
assign pe0_act_buffer_addr10 = n390 ? (n654) : (n353 ? (n379) : (0)) ;
assign pe0_act_buffer_data10 = n390 ? (n679) : (n353 ? (data_in_5) : ('d0)) ;
assign pe0_act_buffer_wen10 = (n390) ? ( 1'b1 ) : ((n353) ? ( 1'b1 ) : (1'b0)) ;
assign pe0_act_buffer_addr11 = n390 ? (n680) : (n353 ? (n381) : (0)) ;
assign pe0_act_buffer_data11 = n390 ? (n704) : (n353 ? (data_in_4) : ('d0)) ;
assign pe0_act_buffer_wen11 = (n390) ? ( 1'b1 ) : ((n353) ? ( 1'b1 ) : (1'b0)) ;
assign pe0_act_buffer_addr12 = n390 ? (n705) : (n353 ? (n383) : (0)) ;
assign pe0_act_buffer_data12 = n390 ? (n729) : (n353 ? (data_in_3) : ('d0)) ;
assign pe0_act_buffer_wen12 = (n390) ? ( 1'b1 ) : ((n353) ? ( 1'b1 ) : (1'b0)) ;
assign pe0_act_buffer_addr13 = n390 ? (n730) : (n353 ? (n385) : (0)) ;
assign pe0_act_buffer_data13 = n390 ? (n754) : (n353 ? (data_in_2) : ('d0)) ;
assign pe0_act_buffer_wen13 = (n390) ? ( 1'b1 ) : ((n353) ? ( 1'b1 ) : (1'b0)) ;
assign pe0_act_buffer_addr14 = n390 ? (n755) : (n353 ? (n387) : (0)) ;
assign pe0_act_buffer_data14 = n390 ? (n779) : (n353 ? (data_in_1) : ('d0)) ;
assign pe0_act_buffer_wen14 = (n390) ? ( 1'b1 ) : ((n353) ? ( 1'b1 ) : (1'b0)) ;
assign pe0_act_buffer_addr15 = n390 ? (n780) : (n353 ? (n389) : (0)) ;
assign pe0_act_buffer_data15 = n390 ? (n804) : (n353 ? (data_in_0) : ('d0)) ;
assign pe0_act_buffer_wen15 = (n390) ? ( 1'b1 ) : ((n353) ? ( 1'b1 ) : (1'b0)) ;
assign n805 =  ( pe0_act_instruction_counter ) + ( bv_6_1_n108 )  ;
assign n806 =  ( n247 ) ? ( bv_6_0_n110 ) : ( n805 ) ;
assign n807 =  ( pe0_act_instruction_counter ) + ( bv_6_1_n108 )  ;
assign n808 =  ( n254 ) ? ( bv_6_0_n110 ) : ( n807 ) ;
assign n809 =  ( pe0_act_instruction_counter ) + ( bv_6_1_n108 )  ;
assign n810 =  ( n260 ) ? ( bv_6_0_n110 ) : ( n809 ) ;
assign n811 =  ( pe0_act_instruction_counter ) + ( bv_6_1_n108 )  ;
assign n812 =  ( n266 ) ? ( bv_6_0_n110 ) : ( n811 ) ;
assign n813 =  ( pe0_act_instruction_counter ) + ( bv_6_1_n108 )  ;
assign n814 =  ( n272 ) ? ( bv_6_0_n110 ) : ( n813 ) ;
assign n815 =  ( pe0_act_instruction_counter ) + ( bv_6_1_n108 )  ;
assign n816 =  ( n278 ) ? ( bv_6_0_n110 ) : ( n815 ) ;
assign n817 =  ( pe0_act_instruction_counter ) + ( bv_6_1_n108 )  ;
assign n818 =  ( n284 ) ? ( bv_6_0_n110 ) : ( n817 ) ;
assign n819 =  ( pe0_act_instruction_counter ) + ( bv_6_1_n108 )  ;
assign n820 =  ( n290 ) ? ( bv_6_0_n110 ) : ( n819 ) ;
assign n821 =  ( pe0_act_instruction_counter ) + ( bv_6_1_n108 )  ;
assign n822 =  ( n296 ) ? ( bv_6_0_n110 ) : ( n821 ) ;
assign n823 =  ( pe0_act_instruction_counter ) + ( bv_6_1_n108 )  ;
assign n824 =  ( n302 ) ? ( bv_6_0_n110 ) : ( n823 ) ;
assign n825 =  ( pe0_act_instruction_counter ) + ( bv_6_1_n108 )  ;
assign n826 =  ( n308 ) ? ( bv_6_0_n110 ) : ( n825 ) ;
assign n827 =  ( pe0_act_instruction_counter ) + ( bv_6_1_n108 )  ;
assign n828 =  ( n314 ) ? ( bv_6_0_n110 ) : ( n827 ) ;
assign n829 = ~ ( n250 )  ;
assign n830 =  ( n247 ) & (n829 )  ;
assign n831 =  ( pe0_act_output_counter ) + ( bv_8_1_n248 )  ;
assign n832 =  ( n830 ) ? ( n831 ) : ( pe0_act_output_counter ) ;
assign n833 =  ( n251 ) ? ( bv_8_0_n354 ) : ( n832 ) ;
assign n834 = ~ ( n256 )  ;
assign n835 =  ( n254 ) & (n834 )  ;
assign n836 =  ( pe0_act_output_counter ) + ( bv_8_1_n248 )  ;
assign n837 =  ( n835 ) ? ( n836 ) : ( pe0_act_output_counter ) ;
assign n838 =  ( n257 ) ? ( bv_8_0_n354 ) : ( n837 ) ;
assign n839 = ~ ( n262 )  ;
assign n840 =  ( n260 ) & (n839 )  ;
assign n841 =  ( pe0_act_output_counter ) + ( bv_8_1_n248 )  ;
assign n842 =  ( n840 ) ? ( n841 ) : ( pe0_act_output_counter ) ;
assign n843 =  ( n263 ) ? ( bv_8_0_n354 ) : ( n842 ) ;
assign n844 = ~ ( n268 )  ;
assign n845 =  ( n266 ) & (n844 )  ;
assign n846 =  ( pe0_act_output_counter ) + ( bv_8_1_n248 )  ;
assign n847 =  ( n845 ) ? ( n846 ) : ( pe0_act_output_counter ) ;
assign n848 =  ( n269 ) ? ( bv_8_0_n354 ) : ( n847 ) ;
assign n849 = ~ ( n274 )  ;
assign n850 =  ( n272 ) & (n849 )  ;
assign n851 =  ( pe0_act_output_counter ) + ( bv_8_1_n248 )  ;
assign n852 =  ( n850 ) ? ( n851 ) : ( pe0_act_output_counter ) ;
assign n853 =  ( n275 ) ? ( bv_8_0_n354 ) : ( n852 ) ;
assign n854 = ~ ( n280 )  ;
assign n855 =  ( n278 ) & (n854 )  ;
assign n856 =  ( pe0_act_output_counter ) + ( bv_8_1_n248 )  ;
assign n857 =  ( n855 ) ? ( n856 ) : ( pe0_act_output_counter ) ;
assign n858 =  ( n281 ) ? ( bv_8_0_n354 ) : ( n857 ) ;
assign n859 = ~ ( n286 )  ;
assign n860 =  ( n284 ) & (n859 )  ;
assign n861 =  ( pe0_act_output_counter ) + ( bv_8_1_n248 )  ;
assign n862 =  ( n860 ) ? ( n861 ) : ( pe0_act_output_counter ) ;
assign n863 =  ( n287 ) ? ( bv_8_0_n354 ) : ( n862 ) ;
assign n864 = ~ ( n292 )  ;
assign n865 =  ( n290 ) & (n864 )  ;
assign n866 =  ( pe0_act_output_counter ) + ( bv_8_1_n248 )  ;
assign n867 =  ( n865 ) ? ( n866 ) : ( pe0_act_output_counter ) ;
assign n868 =  ( n293 ) ? ( bv_8_0_n354 ) : ( n867 ) ;
assign n869 = ~ ( n298 )  ;
assign n870 =  ( n296 ) & (n869 )  ;
assign n871 =  ( pe0_act_output_counter ) + ( bv_8_1_n248 )  ;
assign n872 =  ( n870 ) ? ( n871 ) : ( pe0_act_output_counter ) ;
assign n873 =  ( n299 ) ? ( bv_8_0_n354 ) : ( n872 ) ;
assign n874 = ~ ( n304 )  ;
assign n875 =  ( n302 ) & (n874 )  ;
assign n876 =  ( pe0_act_output_counter ) + ( bv_8_1_n248 )  ;
assign n877 =  ( n875 ) ? ( n876 ) : ( pe0_act_output_counter ) ;
assign n878 =  ( n305 ) ? ( bv_8_0_n354 ) : ( n877 ) ;
assign n879 = ~ ( n310 )  ;
assign n880 =  ( n308 ) & (n879 )  ;
assign n881 =  ( pe0_act_output_counter ) + ( bv_8_1_n248 )  ;
assign n882 =  ( n880 ) ? ( n881 ) : ( pe0_act_output_counter ) ;
assign n883 =  ( n311 ) ? ( bv_8_0_n354 ) : ( n882 ) ;
assign n884 = ~ ( n316 )  ;
assign n885 =  ( n314 ) & (n884 )  ;
assign n886 =  ( pe0_act_output_counter ) + ( bv_8_1_n248 )  ;
assign n887 =  ( n885 ) ? ( n886 ) : ( pe0_act_output_counter ) ;
assign n888 =  ( n317 ) ? ( bv_8_0_n354 ) : ( n887 ) ;
assign n889 = ~ ( n43 )  ;
assign n890 =  ( 1'b1 ) & (n889 )  ;
assign n891 =  ( 1'b1 ) & (n43 )  ;
assign n892 =  ( bv_4_15_n401 ) + ( bv_4_0_n402 )  ;
assign n893 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n894 =  ( bv_4_14_n429 ) + ( bv_4_0_n402 )  ;
assign n895 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n896 =  ( bv_4_13_n220 ) + ( bv_4_0_n402 )  ;
assign n897 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n898 =  ( bv_4_12_n214 ) + ( bv_4_0_n402 )  ;
assign n899 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n900 =  ( bv_4_11_n208 ) + ( bv_4_0_n402 )  ;
assign n901 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n902 =  ( bv_4_10_n202 ) + ( bv_4_0_n402 )  ;
assign n903 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n904 =  ( bv_4_9_n196 ) + ( bv_4_0_n402 )  ;
assign n905 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n906 =  ( bv_4_8_n190 ) + ( bv_4_0_n402 )  ;
assign n907 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n908 =  ( bv_4_7_n184 ) + ( bv_4_0_n402 )  ;
assign n909 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n910 =  ( bv_4_6_n630 ) + ( bv_4_0_n402 )  ;
assign n911 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n912 =  ( bv_4_5_n656 ) + ( bv_4_0_n402 )  ;
assign n913 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n914 =  ( bv_4_4_n176 ) + ( bv_4_0_n402 )  ;
assign n915 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n916 =  ( bv_4_3_n166 ) + ( bv_4_0_n402 )  ;
assign n917 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n918 =  ( bv_4_2_n160 ) + ( bv_4_0_n402 )  ;
assign n919 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n920 =  ( bv_4_1_n145 ) + ( bv_4_0_n402 )  ;
assign n921 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n922 =  ( bv_4_0_n402 ) + ( bv_4_0_n402 )  ;
assign n923 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign PE0_act_regs_0_addr0 = n891 ? (n892) : (0) ;
assign PE0_act_regs_0_data0 = n891 ? (n893) : ('d0) ;
assign PE0_act_regs_0_wen0 = (n891) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_0_addr1 = n891 ? (n894) : (0) ;
assign PE0_act_regs_0_data1 = n891 ? (n895) : ('d0) ;
assign PE0_act_regs_0_wen1 = (n891) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_0_addr2 = n891 ? (n896) : (0) ;
assign PE0_act_regs_0_data2 = n891 ? (n897) : ('d0) ;
assign PE0_act_regs_0_wen2 = (n891) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_0_addr3 = n891 ? (n898) : (0) ;
assign PE0_act_regs_0_data3 = n891 ? (n899) : ('d0) ;
assign PE0_act_regs_0_wen3 = (n891) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_0_addr4 = n891 ? (n900) : (0) ;
assign PE0_act_regs_0_data4 = n891 ? (n901) : ('d0) ;
assign PE0_act_regs_0_wen4 = (n891) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_0_addr5 = n891 ? (n902) : (0) ;
assign PE0_act_regs_0_data5 = n891 ? (n903) : ('d0) ;
assign PE0_act_regs_0_wen5 = (n891) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_0_addr6 = n891 ? (n904) : (0) ;
assign PE0_act_regs_0_data6 = n891 ? (n905) : ('d0) ;
assign PE0_act_regs_0_wen6 = (n891) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_0_addr7 = n891 ? (n906) : (0) ;
assign PE0_act_regs_0_data7 = n891 ? (n907) : ('d0) ;
assign PE0_act_regs_0_wen7 = (n891) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_0_addr8 = n891 ? (n908) : (0) ;
assign PE0_act_regs_0_data8 = n891 ? (n909) : ('d0) ;
assign PE0_act_regs_0_wen8 = (n891) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_0_addr9 = n891 ? (n910) : (0) ;
assign PE0_act_regs_0_data9 = n891 ? (n911) : ('d0) ;
assign PE0_act_regs_0_wen9 = (n891) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_0_addr10 = n891 ? (n912) : (0) ;
assign PE0_act_regs_0_data10 = n891 ? (n913) : ('d0) ;
assign PE0_act_regs_0_wen10 = (n891) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_0_addr11 = n891 ? (n914) : (0) ;
assign PE0_act_regs_0_data11 = n891 ? (n915) : ('d0) ;
assign PE0_act_regs_0_wen11 = (n891) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_0_addr12 = n891 ? (n916) : (0) ;
assign PE0_act_regs_0_data12 = n891 ? (n917) : ('d0) ;
assign PE0_act_regs_0_wen12 = (n891) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_0_addr13 = n891 ? (n918) : (0) ;
assign PE0_act_regs_0_data13 = n891 ? (n919) : ('d0) ;
assign PE0_act_regs_0_wen13 = (n891) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_0_addr14 = n891 ? (n920) : (0) ;
assign PE0_act_regs_0_data14 = n891 ? (n921) : ('d0) ;
assign PE0_act_regs_0_wen14 = (n891) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_0_addr15 = n891 ? (n922) : (0) ;
assign PE0_act_regs_0_data15 = n891 ? (n923) : ('d0) ;
assign PE0_act_regs_0_wen15 = (n891) ? ( 1'b1 ) : (1'b0) ;
assign n924 = ~ ( n43 )  ;
assign n925 =  ( 1'b1 ) & (n924 )  ;
assign n926 =  ( 1'b1 ) & (n43 )  ;
assign n927 =  ( bv_4_15_n401 ) + ( bv_4_0_n402 )  ;
assign n928 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n929 =  ( bv_4_14_n429 ) + ( bv_4_0_n402 )  ;
assign n930 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n931 =  ( bv_4_13_n220 ) + ( bv_4_0_n402 )  ;
assign n932 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n933 =  ( bv_4_12_n214 ) + ( bv_4_0_n402 )  ;
assign n934 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n935 =  ( bv_4_11_n208 ) + ( bv_4_0_n402 )  ;
assign n936 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n937 =  ( bv_4_10_n202 ) + ( bv_4_0_n402 )  ;
assign n938 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n939 =  ( bv_4_9_n196 ) + ( bv_4_0_n402 )  ;
assign n940 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n941 =  ( bv_4_8_n190 ) + ( bv_4_0_n402 )  ;
assign n942 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n943 =  ( bv_4_7_n184 ) + ( bv_4_0_n402 )  ;
assign n944 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n945 =  ( bv_4_6_n630 ) + ( bv_4_0_n402 )  ;
assign n946 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n947 =  ( bv_4_5_n656 ) + ( bv_4_0_n402 )  ;
assign n948 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n949 =  ( bv_4_4_n176 ) + ( bv_4_0_n402 )  ;
assign n950 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n951 =  ( bv_4_3_n166 ) + ( bv_4_0_n402 )  ;
assign n952 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n953 =  ( bv_4_2_n160 ) + ( bv_4_0_n402 )  ;
assign n954 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n955 =  ( bv_4_1_n145 ) + ( bv_4_0_n402 )  ;
assign n956 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n957 =  ( bv_4_0_n402 ) + ( bv_4_0_n402 )  ;
assign n958 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign PE0_act_regs_1_addr0 = n926 ? (n927) : (0) ;
assign PE0_act_regs_1_data0 = n926 ? (n928) : ('d0) ;
assign PE0_act_regs_1_wen0 = (n926) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_1_addr1 = n926 ? (n929) : (0) ;
assign PE0_act_regs_1_data1 = n926 ? (n930) : ('d0) ;
assign PE0_act_regs_1_wen1 = (n926) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_1_addr2 = n926 ? (n931) : (0) ;
assign PE0_act_regs_1_data2 = n926 ? (n932) : ('d0) ;
assign PE0_act_regs_1_wen2 = (n926) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_1_addr3 = n926 ? (n933) : (0) ;
assign PE0_act_regs_1_data3 = n926 ? (n934) : ('d0) ;
assign PE0_act_regs_1_wen3 = (n926) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_1_addr4 = n926 ? (n935) : (0) ;
assign PE0_act_regs_1_data4 = n926 ? (n936) : ('d0) ;
assign PE0_act_regs_1_wen4 = (n926) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_1_addr5 = n926 ? (n937) : (0) ;
assign PE0_act_regs_1_data5 = n926 ? (n938) : ('d0) ;
assign PE0_act_regs_1_wen5 = (n926) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_1_addr6 = n926 ? (n939) : (0) ;
assign PE0_act_regs_1_data6 = n926 ? (n940) : ('d0) ;
assign PE0_act_regs_1_wen6 = (n926) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_1_addr7 = n926 ? (n941) : (0) ;
assign PE0_act_regs_1_data7 = n926 ? (n942) : ('d0) ;
assign PE0_act_regs_1_wen7 = (n926) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_1_addr8 = n926 ? (n943) : (0) ;
assign PE0_act_regs_1_data8 = n926 ? (n944) : ('d0) ;
assign PE0_act_regs_1_wen8 = (n926) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_1_addr9 = n926 ? (n945) : (0) ;
assign PE0_act_regs_1_data9 = n926 ? (n946) : ('d0) ;
assign PE0_act_regs_1_wen9 = (n926) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_1_addr10 = n926 ? (n947) : (0) ;
assign PE0_act_regs_1_data10 = n926 ? (n948) : ('d0) ;
assign PE0_act_regs_1_wen10 = (n926) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_1_addr11 = n926 ? (n949) : (0) ;
assign PE0_act_regs_1_data11 = n926 ? (n950) : ('d0) ;
assign PE0_act_regs_1_wen11 = (n926) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_1_addr12 = n926 ? (n951) : (0) ;
assign PE0_act_regs_1_data12 = n926 ? (n952) : ('d0) ;
assign PE0_act_regs_1_wen12 = (n926) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_1_addr13 = n926 ? (n953) : (0) ;
assign PE0_act_regs_1_data13 = n926 ? (n954) : ('d0) ;
assign PE0_act_regs_1_wen13 = (n926) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_1_addr14 = n926 ? (n955) : (0) ;
assign PE0_act_regs_1_data14 = n926 ? (n956) : ('d0) ;
assign PE0_act_regs_1_wen14 = (n926) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_1_addr15 = n926 ? (n957) : (0) ;
assign PE0_act_regs_1_data15 = n926 ? (n958) : ('d0) ;
assign PE0_act_regs_1_wen15 = (n926) ? ( 1'b1 ) : (1'b0) ;
assign n959 = ~ ( n43 )  ;
assign n960 =  ( 1'b1 ) & (n959 )  ;
assign n961 =  ( 1'b1 ) & (n43 )  ;
assign n962 =  ( bv_4_15_n401 ) + ( bv_4_0_n402 )  ;
assign n963 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n964 =  ( bv_4_14_n429 ) + ( bv_4_0_n402 )  ;
assign n965 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n966 =  ( bv_4_13_n220 ) + ( bv_4_0_n402 )  ;
assign n967 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n968 =  ( bv_4_12_n214 ) + ( bv_4_0_n402 )  ;
assign n969 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n970 =  ( bv_4_11_n208 ) + ( bv_4_0_n402 )  ;
assign n971 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n972 =  ( bv_4_10_n202 ) + ( bv_4_0_n402 )  ;
assign n973 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n974 =  ( bv_4_9_n196 ) + ( bv_4_0_n402 )  ;
assign n975 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n976 =  ( bv_4_8_n190 ) + ( bv_4_0_n402 )  ;
assign n977 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n978 =  ( bv_4_7_n184 ) + ( bv_4_0_n402 )  ;
assign n979 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n980 =  ( bv_4_6_n630 ) + ( bv_4_0_n402 )  ;
assign n981 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n982 =  ( bv_4_5_n656 ) + ( bv_4_0_n402 )  ;
assign n983 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n984 =  ( bv_4_4_n176 ) + ( bv_4_0_n402 )  ;
assign n985 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n986 =  ( bv_4_3_n166 ) + ( bv_4_0_n402 )  ;
assign n987 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n988 =  ( bv_4_2_n160 ) + ( bv_4_0_n402 )  ;
assign n989 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n990 =  ( bv_4_1_n145 ) + ( bv_4_0_n402 )  ;
assign n991 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n992 =  ( bv_4_0_n402 ) + ( bv_4_0_n402 )  ;
assign n993 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign PE0_act_regs_2_addr0 = n961 ? (n962) : (0) ;
assign PE0_act_regs_2_data0 = n961 ? (n963) : ('d0) ;
assign PE0_act_regs_2_wen0 = (n961) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_2_addr1 = n961 ? (n964) : (0) ;
assign PE0_act_regs_2_data1 = n961 ? (n965) : ('d0) ;
assign PE0_act_regs_2_wen1 = (n961) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_2_addr2 = n961 ? (n966) : (0) ;
assign PE0_act_regs_2_data2 = n961 ? (n967) : ('d0) ;
assign PE0_act_regs_2_wen2 = (n961) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_2_addr3 = n961 ? (n968) : (0) ;
assign PE0_act_regs_2_data3 = n961 ? (n969) : ('d0) ;
assign PE0_act_regs_2_wen3 = (n961) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_2_addr4 = n961 ? (n970) : (0) ;
assign PE0_act_regs_2_data4 = n961 ? (n971) : ('d0) ;
assign PE0_act_regs_2_wen4 = (n961) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_2_addr5 = n961 ? (n972) : (0) ;
assign PE0_act_regs_2_data5 = n961 ? (n973) : ('d0) ;
assign PE0_act_regs_2_wen5 = (n961) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_2_addr6 = n961 ? (n974) : (0) ;
assign PE0_act_regs_2_data6 = n961 ? (n975) : ('d0) ;
assign PE0_act_regs_2_wen6 = (n961) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_2_addr7 = n961 ? (n976) : (0) ;
assign PE0_act_regs_2_data7 = n961 ? (n977) : ('d0) ;
assign PE0_act_regs_2_wen7 = (n961) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_2_addr8 = n961 ? (n978) : (0) ;
assign PE0_act_regs_2_data8 = n961 ? (n979) : ('d0) ;
assign PE0_act_regs_2_wen8 = (n961) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_2_addr9 = n961 ? (n980) : (0) ;
assign PE0_act_regs_2_data9 = n961 ? (n981) : ('d0) ;
assign PE0_act_regs_2_wen9 = (n961) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_2_addr10 = n961 ? (n982) : (0) ;
assign PE0_act_regs_2_data10 = n961 ? (n983) : ('d0) ;
assign PE0_act_regs_2_wen10 = (n961) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_2_addr11 = n961 ? (n984) : (0) ;
assign PE0_act_regs_2_data11 = n961 ? (n985) : ('d0) ;
assign PE0_act_regs_2_wen11 = (n961) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_2_addr12 = n961 ? (n986) : (0) ;
assign PE0_act_regs_2_data12 = n961 ? (n987) : ('d0) ;
assign PE0_act_regs_2_wen12 = (n961) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_2_addr13 = n961 ? (n988) : (0) ;
assign PE0_act_regs_2_data13 = n961 ? (n989) : ('d0) ;
assign PE0_act_regs_2_wen13 = (n961) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_2_addr14 = n961 ? (n990) : (0) ;
assign PE0_act_regs_2_data14 = n961 ? (n991) : ('d0) ;
assign PE0_act_regs_2_wen14 = (n961) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_2_addr15 = n961 ? (n992) : (0) ;
assign PE0_act_regs_2_data15 = n961 ? (n993) : ('d0) ;
assign PE0_act_regs_2_wen15 = (n961) ? ( 1'b1 ) : (1'b0) ;
assign n994 = ~ ( n43 )  ;
assign n995 =  ( 1'b1 ) & (n994 )  ;
assign n996 =  ( 1'b1 ) & (n43 )  ;
assign n997 =  ( bv_4_15_n401 ) + ( bv_4_0_n402 )  ;
assign n998 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n999 =  ( bv_4_14_n429 ) + ( bv_4_0_n402 )  ;
assign n1000 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n1001 =  ( bv_4_13_n220 ) + ( bv_4_0_n402 )  ;
assign n1002 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n1003 =  ( bv_4_12_n214 ) + ( bv_4_0_n402 )  ;
assign n1004 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n1005 =  ( bv_4_11_n208 ) + ( bv_4_0_n402 )  ;
assign n1006 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n1007 =  ( bv_4_10_n202 ) + ( bv_4_0_n402 )  ;
assign n1008 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n1009 =  ( bv_4_9_n196 ) + ( bv_4_0_n402 )  ;
assign n1010 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n1011 =  ( bv_4_8_n190 ) + ( bv_4_0_n402 )  ;
assign n1012 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n1013 =  ( bv_4_7_n184 ) + ( bv_4_0_n402 )  ;
assign n1014 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n1015 =  ( bv_4_6_n630 ) + ( bv_4_0_n402 )  ;
assign n1016 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n1017 =  ( bv_4_5_n656 ) + ( bv_4_0_n402 )  ;
assign n1018 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n1019 =  ( bv_4_4_n176 ) + ( bv_4_0_n402 )  ;
assign n1020 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n1021 =  ( bv_4_3_n166 ) + ( bv_4_0_n402 )  ;
assign n1022 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n1023 =  ( bv_4_2_n160 ) + ( bv_4_0_n402 )  ;
assign n1024 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n1025 =  ( bv_4_1_n145 ) + ( bv_4_0_n402 )  ;
assign n1026 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n1027 =  ( bv_4_0_n402 ) + ( bv_4_0_n402 )  ;
assign n1028 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign PE0_act_regs_3_addr0 = n996 ? (n997) : (0) ;
assign PE0_act_regs_3_data0 = n996 ? (n998) : ('d0) ;
assign PE0_act_regs_3_wen0 = (n996) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_3_addr1 = n996 ? (n999) : (0) ;
assign PE0_act_regs_3_data1 = n996 ? (n1000) : ('d0) ;
assign PE0_act_regs_3_wen1 = (n996) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_3_addr2 = n996 ? (n1001) : (0) ;
assign PE0_act_regs_3_data2 = n996 ? (n1002) : ('d0) ;
assign PE0_act_regs_3_wen2 = (n996) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_3_addr3 = n996 ? (n1003) : (0) ;
assign PE0_act_regs_3_data3 = n996 ? (n1004) : ('d0) ;
assign PE0_act_regs_3_wen3 = (n996) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_3_addr4 = n996 ? (n1005) : (0) ;
assign PE0_act_regs_3_data4 = n996 ? (n1006) : ('d0) ;
assign PE0_act_regs_3_wen4 = (n996) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_3_addr5 = n996 ? (n1007) : (0) ;
assign PE0_act_regs_3_data5 = n996 ? (n1008) : ('d0) ;
assign PE0_act_regs_3_wen5 = (n996) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_3_addr6 = n996 ? (n1009) : (0) ;
assign PE0_act_regs_3_data6 = n996 ? (n1010) : ('d0) ;
assign PE0_act_regs_3_wen6 = (n996) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_3_addr7 = n996 ? (n1011) : (0) ;
assign PE0_act_regs_3_data7 = n996 ? (n1012) : ('d0) ;
assign PE0_act_regs_3_wen7 = (n996) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_3_addr8 = n996 ? (n1013) : (0) ;
assign PE0_act_regs_3_data8 = n996 ? (n1014) : ('d0) ;
assign PE0_act_regs_3_wen8 = (n996) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_3_addr9 = n996 ? (n1015) : (0) ;
assign PE0_act_regs_3_data9 = n996 ? (n1016) : ('d0) ;
assign PE0_act_regs_3_wen9 = (n996) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_3_addr10 = n996 ? (n1017) : (0) ;
assign PE0_act_regs_3_data10 = n996 ? (n1018) : ('d0) ;
assign PE0_act_regs_3_wen10 = (n996) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_3_addr11 = n996 ? (n1019) : (0) ;
assign PE0_act_regs_3_data11 = n996 ? (n1020) : ('d0) ;
assign PE0_act_regs_3_wen11 = (n996) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_3_addr12 = n996 ? (n1021) : (0) ;
assign PE0_act_regs_3_data12 = n996 ? (n1022) : ('d0) ;
assign PE0_act_regs_3_wen12 = (n996) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_3_addr13 = n996 ? (n1023) : (0) ;
assign PE0_act_regs_3_data13 = n996 ? (n1024) : ('d0) ;
assign PE0_act_regs_3_wen13 = (n996) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_3_addr14 = n996 ? (n1025) : (0) ;
assign PE0_act_regs_3_data14 = n996 ? (n1026) : ('d0) ;
assign PE0_act_regs_3_wen14 = (n996) ? ( 1'b1 ) : (1'b0) ;
assign PE0_act_regs_3_addr15 = n996 ? (n1027) : (0) ;
assign PE0_act_regs_3_data15 = n996 ? (n1028) : ('d0) ;
assign PE0_act_regs_3_wen15 = (n996) ? ( 1'b1 ) : (1'b0) ;
assign n1029 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n1030 =  { ( bv_24_0_n391 ) , ( pe0_act_output_counter ) }  ;
assign n1031 =  { ( bv_27_0_n393 ) , ( pe0_act_mngr_buffer_addr_base ) }  ;
assign n1032 =  ( n1030 ) + ( n1031 )  ;
assign n1033 =  ( n1032 ) << ( bv_32_4_n380 )  ;
assign n1034 =  ( n1033 ) + ( bv_32_0_n388 )  ;
assign pe0_act_buffer_addr_n1035 = n1034 ;
assign n1037 = pe0_act_buffer_data_n1036 ;
fun_Adptfloat2Fixed  applyFunc_n1039(
    .arg0( n1037 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n1038 )
);
assign n1040 = n1038 ;
assign n1041 = n143[1:0] ;
assign n1042 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n1043 =  ( bv_4_0_n402 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1044 = n1043 ;
assign n1046 = PE0_act_regs_3_data_n1045 ;
assign n1047 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1048 = n1043 ;
assign n1050 = PE0_act_regs_2_data_n1049 ;
assign n1051 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1052 = n1043 ;
assign n1054 = PE0_act_regs_1_data_n1053 ;
assign n1055 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1056 = n1043 ;
assign n1058 = PE0_act_regs_0_data_n1057 ;
assign n1059 =  ( n1055 ) ? ( n1058 ) : ( bv_20_0_n419 ) ;
assign n1060 =  ( n1051 ) ? ( n1054 ) : ( n1059 ) ;
assign n1061 =  ( n1047 ) ? ( n1050 ) : ( n1060 ) ;
assign n1062 =  ( n1042 ) ? ( n1046 ) : ( n1061 ) ;
assign n1063 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n1064 =  ( bv_4_0_n402 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1065 = n1064 ;
assign n1067 = PE0_act_regs_3_data_n1066 ;
assign n1068 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1069 = n1064 ;
assign n1071 = PE0_act_regs_2_data_n1070 ;
assign n1072 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1073 = n1064 ;
assign n1075 = PE0_act_regs_1_data_n1074 ;
assign n1076 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1077 = n1064 ;
assign n1079 = PE0_act_regs_0_data_n1078 ;
assign n1080 =  ( n1076 ) ? ( n1079 ) : ( bv_20_0_n419 ) ;
assign n1081 =  ( n1072 ) ? ( n1075 ) : ( n1080 ) ;
assign n1082 =  ( n1068 ) ? ( n1071 ) : ( n1081 ) ;
assign n1083 =  ( n1063 ) ? ( n1067 ) : ( n1082 ) ;
assign n1084 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n1085 = n1064 ;
assign n1087 = PE0_act_regs_3_data_n1086 ;
assign n1088 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1089 = n1064 ;
assign n1091 = PE0_act_regs_2_data_n1090 ;
assign n1092 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1093 = n1064 ;
assign n1095 = PE0_act_regs_1_data_n1094 ;
assign n1096 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1097 = n1064 ;
assign n1099 = PE0_act_regs_0_data_n1098 ;
assign n1100 =  ( n1096 ) ? ( n1099 ) : ( bv_20_0_n419 ) ;
assign n1101 =  ( n1092 ) ? ( n1095 ) : ( n1100 ) ;
assign n1102 =  ( n1088 ) ? ( n1091 ) : ( n1101 ) ;
assign n1103 =  ( n1084 ) ? ( n1087 ) : ( n1102 ) ;
fun_PEActEadd  applyFunc_n1105(
    .arg0( n1083 ),
    .arg1( n1103 ),
    .result( n1104 )
);
assign n1106 = n1104 ;
assign n1107 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n1108 =  ( bv_4_0_n402 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1109 = n1108 ;
assign n1111 = PE0_act_regs_3_data_n1110 ;
assign n1112 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1113 = n1108 ;
assign n1115 = PE0_act_regs_2_data_n1114 ;
assign n1116 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1117 = n1108 ;
assign n1119 = PE0_act_regs_1_data_n1118 ;
assign n1120 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1121 = n1108 ;
assign n1123 = PE0_act_regs_0_data_n1122 ;
assign n1124 =  ( n1120 ) ? ( n1123 ) : ( bv_20_0_n419 ) ;
assign n1125 =  ( n1116 ) ? ( n1119 ) : ( n1124 ) ;
assign n1126 =  ( n1112 ) ? ( n1115 ) : ( n1125 ) ;
assign n1127 =  ( n1107 ) ? ( n1111 ) : ( n1126 ) ;
assign n1128 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n1129 = n1108 ;
assign n1131 = PE0_act_regs_3_data_n1130 ;
assign n1132 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1133 = n1108 ;
assign n1135 = PE0_act_regs_2_data_n1134 ;
assign n1136 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1137 = n1108 ;
assign n1139 = PE0_act_regs_1_data_n1138 ;
assign n1140 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1141 = n1108 ;
assign n1143 = PE0_act_regs_0_data_n1142 ;
assign n1144 =  ( n1140 ) ? ( n1143 ) : ( bv_20_0_n419 ) ;
assign n1145 =  ( n1136 ) ? ( n1139 ) : ( n1144 ) ;
assign n1146 =  ( n1132 ) ? ( n1135 ) : ( n1145 ) ;
assign n1147 =  ( n1128 ) ? ( n1131 ) : ( n1146 ) ;
fun_PEActEmul  applyFunc_n1149(
    .arg0( n1127 ),
    .arg1( n1147 ),
    .result( n1148 )
);
assign n1150 = n1148 ;
assign n1151 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n1152 =  ( bv_4_0_n402 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1153 = n1152 ;
assign n1155 = PE0_act_regs_3_data_n1154 ;
assign n1156 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1157 = n1152 ;
assign n1159 = PE0_act_regs_2_data_n1158 ;
assign n1160 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1161 = n1152 ;
assign n1163 = PE0_act_regs_1_data_n1162 ;
assign n1164 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1165 = n1152 ;
assign n1167 = PE0_act_regs_0_data_n1166 ;
assign n1168 =  ( n1164 ) ? ( n1167 ) : ( bv_20_0_n419 ) ;
assign n1169 =  ( n1160 ) ? ( n1163 ) : ( n1168 ) ;
assign n1170 =  ( n1156 ) ? ( n1159 ) : ( n1169 ) ;
assign n1171 =  ( n1151 ) ? ( n1155 ) : ( n1170 ) ;
fun_PEActSigmoid  applyFunc_n1173(
    .arg0( n1171 ),
    .result( n1172 )
);
assign n1174 = n1172 ;
assign n1175 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n1176 =  ( bv_4_0_n402 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1177 = n1176 ;
assign n1179 = PE0_act_regs_3_data_n1178 ;
assign n1180 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1181 = n1176 ;
assign n1183 = PE0_act_regs_2_data_n1182 ;
assign n1184 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1185 = n1176 ;
assign n1187 = PE0_act_regs_1_data_n1186 ;
assign n1188 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1189 = n1176 ;
assign n1191 = PE0_act_regs_0_data_n1190 ;
assign n1192 =  ( n1188 ) ? ( n1191 ) : ( bv_20_0_n419 ) ;
assign n1193 =  ( n1184 ) ? ( n1187 ) : ( n1192 ) ;
assign n1194 =  ( n1180 ) ? ( n1183 ) : ( n1193 ) ;
assign n1195 =  ( n1175 ) ? ( n1179 ) : ( n1194 ) ;
fun_PEActTanh  applyFunc_n1197(
    .arg0( n1195 ),
    .result( n1196 )
);
assign n1198 = n1196 ;
assign n1199 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n1200 =  ( bv_4_0_n402 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1201 = n1200 ;
assign n1203 = PE0_act_regs_3_data_n1202 ;
assign n1204 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1205 = n1200 ;
assign n1207 = PE0_act_regs_2_data_n1206 ;
assign n1208 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1209 = n1200 ;
assign n1211 = PE0_act_regs_1_data_n1210 ;
assign n1212 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1213 = n1200 ;
assign n1215 = PE0_act_regs_0_data_n1214 ;
assign n1216 =  ( n1212 ) ? ( n1215 ) : ( bv_20_0_n419 ) ;
assign n1217 =  ( n1208 ) ? ( n1211 ) : ( n1216 ) ;
assign n1218 =  ( n1204 ) ? ( n1207 ) : ( n1217 ) ;
assign n1219 =  ( n1199 ) ? ( n1203 ) : ( n1218 ) ;
fun_PEActRelu  applyFunc_n1221(
    .arg0( n1219 ),
    .result( n1220 )
);
assign n1222 = n1220 ;
assign n1223 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n1224 =  ( bv_4_0_n402 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1225 = n1224 ;
assign n1227 = PE0_act_regs_3_data_n1226 ;
assign n1228 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1229 = n1224 ;
assign n1231 = PE0_act_regs_2_data_n1230 ;
assign n1232 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1233 = n1224 ;
assign n1235 = PE0_act_regs_1_data_n1234 ;
assign n1236 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1237 = n1224 ;
assign n1239 = PE0_act_regs_0_data_n1238 ;
assign n1240 =  ( n1236 ) ? ( n1239 ) : ( bv_20_0_n419 ) ;
assign n1241 =  ( n1232 ) ? ( n1235 ) : ( n1240 ) ;
assign n1242 =  ( n1228 ) ? ( n1231 ) : ( n1241 ) ;
assign n1243 =  ( n1223 ) ? ( n1227 ) : ( n1242 ) ;
fun_PEActOnex  applyFunc_n1245(
    .arg0( n1243 ),
    .result( n1244 )
);
assign n1246 = n1244 ;
assign n1247 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n1248 =  ( n1033 ) + ( bv_32_1_n386 )  ;
assign pe0_act_buffer_addr_n1249 = n1248 ;
assign n1251 = pe0_act_buffer_data_n1250 ;
fun_Adptfloat2Fixed  applyFunc_n1253(
    .arg0( n1251 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n1252 )
);
assign n1254 = n1252 ;
assign n1255 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n1256 =  ( bv_4_1_n145 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1257 = n1256 ;
assign n1259 = PE0_act_regs_3_data_n1258 ;
assign n1260 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1261 = n1256 ;
assign n1263 = PE0_act_regs_2_data_n1262 ;
assign n1264 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1265 = n1256 ;
assign n1267 = PE0_act_regs_1_data_n1266 ;
assign n1268 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1269 = n1256 ;
assign n1271 = PE0_act_regs_0_data_n1270 ;
assign n1272 =  ( n1268 ) ? ( n1271 ) : ( bv_20_0_n419 ) ;
assign n1273 =  ( n1264 ) ? ( n1267 ) : ( n1272 ) ;
assign n1274 =  ( n1260 ) ? ( n1263 ) : ( n1273 ) ;
assign n1275 =  ( n1255 ) ? ( n1259 ) : ( n1274 ) ;
assign n1276 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n1277 =  ( bv_4_1_n145 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1278 = n1277 ;
assign n1280 = PE0_act_regs_3_data_n1279 ;
assign n1281 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1282 = n1277 ;
assign n1284 = PE0_act_regs_2_data_n1283 ;
assign n1285 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1286 = n1277 ;
assign n1288 = PE0_act_regs_1_data_n1287 ;
assign n1289 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1290 = n1277 ;
assign n1292 = PE0_act_regs_0_data_n1291 ;
assign n1293 =  ( n1289 ) ? ( n1292 ) : ( bv_20_0_n419 ) ;
assign n1294 =  ( n1285 ) ? ( n1288 ) : ( n1293 ) ;
assign n1295 =  ( n1281 ) ? ( n1284 ) : ( n1294 ) ;
assign n1296 =  ( n1276 ) ? ( n1280 ) : ( n1295 ) ;
assign n1297 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n1298 = n1277 ;
assign n1300 = PE0_act_regs_3_data_n1299 ;
assign n1301 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1302 = n1277 ;
assign n1304 = PE0_act_regs_2_data_n1303 ;
assign n1305 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1306 = n1277 ;
assign n1308 = PE0_act_regs_1_data_n1307 ;
assign n1309 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1310 = n1277 ;
assign n1312 = PE0_act_regs_0_data_n1311 ;
assign n1313 =  ( n1309 ) ? ( n1312 ) : ( bv_20_0_n419 ) ;
assign n1314 =  ( n1305 ) ? ( n1308 ) : ( n1313 ) ;
assign n1315 =  ( n1301 ) ? ( n1304 ) : ( n1314 ) ;
assign n1316 =  ( n1297 ) ? ( n1300 ) : ( n1315 ) ;
fun_PEActEadd  applyFunc_n1318(
    .arg0( n1296 ),
    .arg1( n1316 ),
    .result( n1317 )
);
assign n1319 = n1317 ;
assign n1320 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n1321 =  ( bv_4_1_n145 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1322 = n1321 ;
assign n1324 = PE0_act_regs_3_data_n1323 ;
assign n1325 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1326 = n1321 ;
assign n1328 = PE0_act_regs_2_data_n1327 ;
assign n1329 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1330 = n1321 ;
assign n1332 = PE0_act_regs_1_data_n1331 ;
assign n1333 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1334 = n1321 ;
assign n1336 = PE0_act_regs_0_data_n1335 ;
assign n1337 =  ( n1333 ) ? ( n1336 ) : ( bv_20_0_n419 ) ;
assign n1338 =  ( n1329 ) ? ( n1332 ) : ( n1337 ) ;
assign n1339 =  ( n1325 ) ? ( n1328 ) : ( n1338 ) ;
assign n1340 =  ( n1320 ) ? ( n1324 ) : ( n1339 ) ;
assign n1341 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n1342 = n1321 ;
assign n1344 = PE0_act_regs_3_data_n1343 ;
assign n1345 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1346 = n1321 ;
assign n1348 = PE0_act_regs_2_data_n1347 ;
assign n1349 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1350 = n1321 ;
assign n1352 = PE0_act_regs_1_data_n1351 ;
assign n1353 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1354 = n1321 ;
assign n1356 = PE0_act_regs_0_data_n1355 ;
assign n1357 =  ( n1353 ) ? ( n1356 ) : ( bv_20_0_n419 ) ;
assign n1358 =  ( n1349 ) ? ( n1352 ) : ( n1357 ) ;
assign n1359 =  ( n1345 ) ? ( n1348 ) : ( n1358 ) ;
assign n1360 =  ( n1341 ) ? ( n1344 ) : ( n1359 ) ;
fun_PEActEmul  applyFunc_n1362(
    .arg0( n1340 ),
    .arg1( n1360 ),
    .result( n1361 )
);
assign n1363 = n1361 ;
assign n1364 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n1365 =  ( bv_4_1_n145 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1366 = n1365 ;
assign n1368 = PE0_act_regs_3_data_n1367 ;
assign n1369 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1370 = n1365 ;
assign n1372 = PE0_act_regs_2_data_n1371 ;
assign n1373 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1374 = n1365 ;
assign n1376 = PE0_act_regs_1_data_n1375 ;
assign n1377 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1378 = n1365 ;
assign n1380 = PE0_act_regs_0_data_n1379 ;
assign n1381 =  ( n1377 ) ? ( n1380 ) : ( bv_20_0_n419 ) ;
assign n1382 =  ( n1373 ) ? ( n1376 ) : ( n1381 ) ;
assign n1383 =  ( n1369 ) ? ( n1372 ) : ( n1382 ) ;
assign n1384 =  ( n1364 ) ? ( n1368 ) : ( n1383 ) ;
fun_PEActSigmoid  applyFunc_n1386(
    .arg0( n1384 ),
    .result( n1385 )
);
assign n1387 = n1385 ;
assign n1388 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n1389 =  ( bv_4_1_n145 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1390 = n1389 ;
assign n1392 = PE0_act_regs_3_data_n1391 ;
assign n1393 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1394 = n1389 ;
assign n1396 = PE0_act_regs_2_data_n1395 ;
assign n1397 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1398 = n1389 ;
assign n1400 = PE0_act_regs_1_data_n1399 ;
assign n1401 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1402 = n1389 ;
assign n1404 = PE0_act_regs_0_data_n1403 ;
assign n1405 =  ( n1401 ) ? ( n1404 ) : ( bv_20_0_n419 ) ;
assign n1406 =  ( n1397 ) ? ( n1400 ) : ( n1405 ) ;
assign n1407 =  ( n1393 ) ? ( n1396 ) : ( n1406 ) ;
assign n1408 =  ( n1388 ) ? ( n1392 ) : ( n1407 ) ;
fun_PEActTanh  applyFunc_n1410(
    .arg0( n1408 ),
    .result( n1409 )
);
assign n1411 = n1409 ;
assign n1412 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n1413 =  ( bv_4_1_n145 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1414 = n1413 ;
assign n1416 = PE0_act_regs_3_data_n1415 ;
assign n1417 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1418 = n1413 ;
assign n1420 = PE0_act_regs_2_data_n1419 ;
assign n1421 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1422 = n1413 ;
assign n1424 = PE0_act_regs_1_data_n1423 ;
assign n1425 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1426 = n1413 ;
assign n1428 = PE0_act_regs_0_data_n1427 ;
assign n1429 =  ( n1425 ) ? ( n1428 ) : ( bv_20_0_n419 ) ;
assign n1430 =  ( n1421 ) ? ( n1424 ) : ( n1429 ) ;
assign n1431 =  ( n1417 ) ? ( n1420 ) : ( n1430 ) ;
assign n1432 =  ( n1412 ) ? ( n1416 ) : ( n1431 ) ;
fun_PEActRelu  applyFunc_n1434(
    .arg0( n1432 ),
    .result( n1433 )
);
assign n1435 = n1433 ;
assign n1436 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n1437 =  ( bv_4_1_n145 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1438 = n1437 ;
assign n1440 = PE0_act_regs_3_data_n1439 ;
assign n1441 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1442 = n1437 ;
assign n1444 = PE0_act_regs_2_data_n1443 ;
assign n1445 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1446 = n1437 ;
assign n1448 = PE0_act_regs_1_data_n1447 ;
assign n1449 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1450 = n1437 ;
assign n1452 = PE0_act_regs_0_data_n1451 ;
assign n1453 =  ( n1449 ) ? ( n1452 ) : ( bv_20_0_n419 ) ;
assign n1454 =  ( n1445 ) ? ( n1448 ) : ( n1453 ) ;
assign n1455 =  ( n1441 ) ? ( n1444 ) : ( n1454 ) ;
assign n1456 =  ( n1436 ) ? ( n1440 ) : ( n1455 ) ;
fun_PEActOnex  applyFunc_n1458(
    .arg0( n1456 ),
    .result( n1457 )
);
assign n1459 = n1457 ;
assign n1460 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n1461 =  ( n1033 ) + ( bv_32_2_n384 )  ;
assign pe0_act_buffer_addr_n1462 = n1461 ;
assign n1464 = pe0_act_buffer_data_n1463 ;
fun_Adptfloat2Fixed  applyFunc_n1466(
    .arg0( n1464 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n1465 )
);
assign n1467 = n1465 ;
assign n1468 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n1469 =  ( bv_4_2_n160 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1470 = n1469 ;
assign n1472 = PE0_act_regs_3_data_n1471 ;
assign n1473 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1474 = n1469 ;
assign n1476 = PE0_act_regs_2_data_n1475 ;
assign n1477 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1478 = n1469 ;
assign n1480 = PE0_act_regs_1_data_n1479 ;
assign n1481 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1482 = n1469 ;
assign n1484 = PE0_act_regs_0_data_n1483 ;
assign n1485 =  ( n1481 ) ? ( n1484 ) : ( bv_20_0_n419 ) ;
assign n1486 =  ( n1477 ) ? ( n1480 ) : ( n1485 ) ;
assign n1487 =  ( n1473 ) ? ( n1476 ) : ( n1486 ) ;
assign n1488 =  ( n1468 ) ? ( n1472 ) : ( n1487 ) ;
assign n1489 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n1490 =  ( bv_4_2_n160 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1491 = n1490 ;
assign n1493 = PE0_act_regs_3_data_n1492 ;
assign n1494 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1495 = n1490 ;
assign n1497 = PE0_act_regs_2_data_n1496 ;
assign n1498 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1499 = n1490 ;
assign n1501 = PE0_act_regs_1_data_n1500 ;
assign n1502 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1503 = n1490 ;
assign n1505 = PE0_act_regs_0_data_n1504 ;
assign n1506 =  ( n1502 ) ? ( n1505 ) : ( bv_20_0_n419 ) ;
assign n1507 =  ( n1498 ) ? ( n1501 ) : ( n1506 ) ;
assign n1508 =  ( n1494 ) ? ( n1497 ) : ( n1507 ) ;
assign n1509 =  ( n1489 ) ? ( n1493 ) : ( n1508 ) ;
assign n1510 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n1511 = n1490 ;
assign n1513 = PE0_act_regs_3_data_n1512 ;
assign n1514 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1515 = n1490 ;
assign n1517 = PE0_act_regs_2_data_n1516 ;
assign n1518 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1519 = n1490 ;
assign n1521 = PE0_act_regs_1_data_n1520 ;
assign n1522 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1523 = n1490 ;
assign n1525 = PE0_act_regs_0_data_n1524 ;
assign n1526 =  ( n1522 ) ? ( n1525 ) : ( bv_20_0_n419 ) ;
assign n1527 =  ( n1518 ) ? ( n1521 ) : ( n1526 ) ;
assign n1528 =  ( n1514 ) ? ( n1517 ) : ( n1527 ) ;
assign n1529 =  ( n1510 ) ? ( n1513 ) : ( n1528 ) ;
fun_PEActEadd  applyFunc_n1531(
    .arg0( n1509 ),
    .arg1( n1529 ),
    .result( n1530 )
);
assign n1532 = n1530 ;
assign n1533 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n1534 =  ( bv_4_2_n160 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1535 = n1534 ;
assign n1537 = PE0_act_regs_3_data_n1536 ;
assign n1538 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1539 = n1534 ;
assign n1541 = PE0_act_regs_2_data_n1540 ;
assign n1542 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1543 = n1534 ;
assign n1545 = PE0_act_regs_1_data_n1544 ;
assign n1546 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1547 = n1534 ;
assign n1549 = PE0_act_regs_0_data_n1548 ;
assign n1550 =  ( n1546 ) ? ( n1549 ) : ( bv_20_0_n419 ) ;
assign n1551 =  ( n1542 ) ? ( n1545 ) : ( n1550 ) ;
assign n1552 =  ( n1538 ) ? ( n1541 ) : ( n1551 ) ;
assign n1553 =  ( n1533 ) ? ( n1537 ) : ( n1552 ) ;
assign n1554 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n1555 = n1534 ;
assign n1557 = PE0_act_regs_3_data_n1556 ;
assign n1558 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1559 = n1534 ;
assign n1561 = PE0_act_regs_2_data_n1560 ;
assign n1562 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1563 = n1534 ;
assign n1565 = PE0_act_regs_1_data_n1564 ;
assign n1566 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1567 = n1534 ;
assign n1569 = PE0_act_regs_0_data_n1568 ;
assign n1570 =  ( n1566 ) ? ( n1569 ) : ( bv_20_0_n419 ) ;
assign n1571 =  ( n1562 ) ? ( n1565 ) : ( n1570 ) ;
assign n1572 =  ( n1558 ) ? ( n1561 ) : ( n1571 ) ;
assign n1573 =  ( n1554 ) ? ( n1557 ) : ( n1572 ) ;
fun_PEActEmul  applyFunc_n1575(
    .arg0( n1553 ),
    .arg1( n1573 ),
    .result( n1574 )
);
assign n1576 = n1574 ;
assign n1577 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n1578 =  ( bv_4_2_n160 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1579 = n1578 ;
assign n1581 = PE0_act_regs_3_data_n1580 ;
assign n1582 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1583 = n1578 ;
assign n1585 = PE0_act_regs_2_data_n1584 ;
assign n1586 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1587 = n1578 ;
assign n1589 = PE0_act_regs_1_data_n1588 ;
assign n1590 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1591 = n1578 ;
assign n1593 = PE0_act_regs_0_data_n1592 ;
assign n1594 =  ( n1590 ) ? ( n1593 ) : ( bv_20_0_n419 ) ;
assign n1595 =  ( n1586 ) ? ( n1589 ) : ( n1594 ) ;
assign n1596 =  ( n1582 ) ? ( n1585 ) : ( n1595 ) ;
assign n1597 =  ( n1577 ) ? ( n1581 ) : ( n1596 ) ;
fun_PEActSigmoid  applyFunc_n1599(
    .arg0( n1597 ),
    .result( n1598 )
);
assign n1600 = n1598 ;
assign n1601 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n1602 =  ( bv_4_2_n160 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1603 = n1602 ;
assign n1605 = PE0_act_regs_3_data_n1604 ;
assign n1606 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1607 = n1602 ;
assign n1609 = PE0_act_regs_2_data_n1608 ;
assign n1610 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1611 = n1602 ;
assign n1613 = PE0_act_regs_1_data_n1612 ;
assign n1614 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1615 = n1602 ;
assign n1617 = PE0_act_regs_0_data_n1616 ;
assign n1618 =  ( n1614 ) ? ( n1617 ) : ( bv_20_0_n419 ) ;
assign n1619 =  ( n1610 ) ? ( n1613 ) : ( n1618 ) ;
assign n1620 =  ( n1606 ) ? ( n1609 ) : ( n1619 ) ;
assign n1621 =  ( n1601 ) ? ( n1605 ) : ( n1620 ) ;
fun_PEActTanh  applyFunc_n1623(
    .arg0( n1621 ),
    .result( n1622 )
);
assign n1624 = n1622 ;
assign n1625 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n1626 =  ( bv_4_2_n160 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1627 = n1626 ;
assign n1629 = PE0_act_regs_3_data_n1628 ;
assign n1630 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1631 = n1626 ;
assign n1633 = PE0_act_regs_2_data_n1632 ;
assign n1634 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1635 = n1626 ;
assign n1637 = PE0_act_regs_1_data_n1636 ;
assign n1638 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1639 = n1626 ;
assign n1641 = PE0_act_regs_0_data_n1640 ;
assign n1642 =  ( n1638 ) ? ( n1641 ) : ( bv_20_0_n419 ) ;
assign n1643 =  ( n1634 ) ? ( n1637 ) : ( n1642 ) ;
assign n1644 =  ( n1630 ) ? ( n1633 ) : ( n1643 ) ;
assign n1645 =  ( n1625 ) ? ( n1629 ) : ( n1644 ) ;
fun_PEActRelu  applyFunc_n1647(
    .arg0( n1645 ),
    .result( n1646 )
);
assign n1648 = n1646 ;
assign n1649 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n1650 =  ( bv_4_2_n160 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1651 = n1650 ;
assign n1653 = PE0_act_regs_3_data_n1652 ;
assign n1654 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1655 = n1650 ;
assign n1657 = PE0_act_regs_2_data_n1656 ;
assign n1658 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1659 = n1650 ;
assign n1661 = PE0_act_regs_1_data_n1660 ;
assign n1662 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1663 = n1650 ;
assign n1665 = PE0_act_regs_0_data_n1664 ;
assign n1666 =  ( n1662 ) ? ( n1665 ) : ( bv_20_0_n419 ) ;
assign n1667 =  ( n1658 ) ? ( n1661 ) : ( n1666 ) ;
assign n1668 =  ( n1654 ) ? ( n1657 ) : ( n1667 ) ;
assign n1669 =  ( n1649 ) ? ( n1653 ) : ( n1668 ) ;
fun_PEActOnex  applyFunc_n1671(
    .arg0( n1669 ),
    .result( n1670 )
);
assign n1672 = n1670 ;
assign n1673 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n1674 =  ( n1033 ) + ( bv_32_3_n382 )  ;
assign pe0_act_buffer_addr_n1675 = n1674 ;
assign n1677 = pe0_act_buffer_data_n1676 ;
fun_Adptfloat2Fixed  applyFunc_n1679(
    .arg0( n1677 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n1678 )
);
assign n1680 = n1678 ;
assign n1681 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n1682 =  ( bv_4_3_n166 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1683 = n1682 ;
assign n1685 = PE0_act_regs_3_data_n1684 ;
assign n1686 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1687 = n1682 ;
assign n1689 = PE0_act_regs_2_data_n1688 ;
assign n1690 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1691 = n1682 ;
assign n1693 = PE0_act_regs_1_data_n1692 ;
assign n1694 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1695 = n1682 ;
assign n1697 = PE0_act_regs_0_data_n1696 ;
assign n1698 =  ( n1694 ) ? ( n1697 ) : ( bv_20_0_n419 ) ;
assign n1699 =  ( n1690 ) ? ( n1693 ) : ( n1698 ) ;
assign n1700 =  ( n1686 ) ? ( n1689 ) : ( n1699 ) ;
assign n1701 =  ( n1681 ) ? ( n1685 ) : ( n1700 ) ;
assign n1702 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n1703 =  ( bv_4_3_n166 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1704 = n1703 ;
assign n1706 = PE0_act_regs_3_data_n1705 ;
assign n1707 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1708 = n1703 ;
assign n1710 = PE0_act_regs_2_data_n1709 ;
assign n1711 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1712 = n1703 ;
assign n1714 = PE0_act_regs_1_data_n1713 ;
assign n1715 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1716 = n1703 ;
assign n1718 = PE0_act_regs_0_data_n1717 ;
assign n1719 =  ( n1715 ) ? ( n1718 ) : ( bv_20_0_n419 ) ;
assign n1720 =  ( n1711 ) ? ( n1714 ) : ( n1719 ) ;
assign n1721 =  ( n1707 ) ? ( n1710 ) : ( n1720 ) ;
assign n1722 =  ( n1702 ) ? ( n1706 ) : ( n1721 ) ;
assign n1723 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n1724 = n1703 ;
assign n1726 = PE0_act_regs_3_data_n1725 ;
assign n1727 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1728 = n1703 ;
assign n1730 = PE0_act_regs_2_data_n1729 ;
assign n1731 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1732 = n1703 ;
assign n1734 = PE0_act_regs_1_data_n1733 ;
assign n1735 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1736 = n1703 ;
assign n1738 = PE0_act_regs_0_data_n1737 ;
assign n1739 =  ( n1735 ) ? ( n1738 ) : ( bv_20_0_n419 ) ;
assign n1740 =  ( n1731 ) ? ( n1734 ) : ( n1739 ) ;
assign n1741 =  ( n1727 ) ? ( n1730 ) : ( n1740 ) ;
assign n1742 =  ( n1723 ) ? ( n1726 ) : ( n1741 ) ;
fun_PEActEadd  applyFunc_n1744(
    .arg0( n1722 ),
    .arg1( n1742 ),
    .result( n1743 )
);
assign n1745 = n1743 ;
assign n1746 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n1747 =  ( bv_4_3_n166 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1748 = n1747 ;
assign n1750 = PE0_act_regs_3_data_n1749 ;
assign n1751 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1752 = n1747 ;
assign n1754 = PE0_act_regs_2_data_n1753 ;
assign n1755 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1756 = n1747 ;
assign n1758 = PE0_act_regs_1_data_n1757 ;
assign n1759 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1760 = n1747 ;
assign n1762 = PE0_act_regs_0_data_n1761 ;
assign n1763 =  ( n1759 ) ? ( n1762 ) : ( bv_20_0_n419 ) ;
assign n1764 =  ( n1755 ) ? ( n1758 ) : ( n1763 ) ;
assign n1765 =  ( n1751 ) ? ( n1754 ) : ( n1764 ) ;
assign n1766 =  ( n1746 ) ? ( n1750 ) : ( n1765 ) ;
assign n1767 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n1768 = n1747 ;
assign n1770 = PE0_act_regs_3_data_n1769 ;
assign n1771 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1772 = n1747 ;
assign n1774 = PE0_act_regs_2_data_n1773 ;
assign n1775 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1776 = n1747 ;
assign n1778 = PE0_act_regs_1_data_n1777 ;
assign n1779 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1780 = n1747 ;
assign n1782 = PE0_act_regs_0_data_n1781 ;
assign n1783 =  ( n1779 ) ? ( n1782 ) : ( bv_20_0_n419 ) ;
assign n1784 =  ( n1775 ) ? ( n1778 ) : ( n1783 ) ;
assign n1785 =  ( n1771 ) ? ( n1774 ) : ( n1784 ) ;
assign n1786 =  ( n1767 ) ? ( n1770 ) : ( n1785 ) ;
fun_PEActEmul  applyFunc_n1788(
    .arg0( n1766 ),
    .arg1( n1786 ),
    .result( n1787 )
);
assign n1789 = n1787 ;
assign n1790 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n1791 =  ( bv_4_3_n166 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1792 = n1791 ;
assign n1794 = PE0_act_regs_3_data_n1793 ;
assign n1795 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1796 = n1791 ;
assign n1798 = PE0_act_regs_2_data_n1797 ;
assign n1799 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1800 = n1791 ;
assign n1802 = PE0_act_regs_1_data_n1801 ;
assign n1803 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1804 = n1791 ;
assign n1806 = PE0_act_regs_0_data_n1805 ;
assign n1807 =  ( n1803 ) ? ( n1806 ) : ( bv_20_0_n419 ) ;
assign n1808 =  ( n1799 ) ? ( n1802 ) : ( n1807 ) ;
assign n1809 =  ( n1795 ) ? ( n1798 ) : ( n1808 ) ;
assign n1810 =  ( n1790 ) ? ( n1794 ) : ( n1809 ) ;
fun_PEActSigmoid  applyFunc_n1812(
    .arg0( n1810 ),
    .result( n1811 )
);
assign n1813 = n1811 ;
assign n1814 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n1815 =  ( bv_4_3_n166 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1816 = n1815 ;
assign n1818 = PE0_act_regs_3_data_n1817 ;
assign n1819 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1820 = n1815 ;
assign n1822 = PE0_act_regs_2_data_n1821 ;
assign n1823 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1824 = n1815 ;
assign n1826 = PE0_act_regs_1_data_n1825 ;
assign n1827 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1828 = n1815 ;
assign n1830 = PE0_act_regs_0_data_n1829 ;
assign n1831 =  ( n1827 ) ? ( n1830 ) : ( bv_20_0_n419 ) ;
assign n1832 =  ( n1823 ) ? ( n1826 ) : ( n1831 ) ;
assign n1833 =  ( n1819 ) ? ( n1822 ) : ( n1832 ) ;
assign n1834 =  ( n1814 ) ? ( n1818 ) : ( n1833 ) ;
fun_PEActTanh  applyFunc_n1836(
    .arg0( n1834 ),
    .result( n1835 )
);
assign n1837 = n1835 ;
assign n1838 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n1839 =  ( bv_4_3_n166 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1840 = n1839 ;
assign n1842 = PE0_act_regs_3_data_n1841 ;
assign n1843 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1844 = n1839 ;
assign n1846 = PE0_act_regs_2_data_n1845 ;
assign n1847 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1848 = n1839 ;
assign n1850 = PE0_act_regs_1_data_n1849 ;
assign n1851 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1852 = n1839 ;
assign n1854 = PE0_act_regs_0_data_n1853 ;
assign n1855 =  ( n1851 ) ? ( n1854 ) : ( bv_20_0_n419 ) ;
assign n1856 =  ( n1847 ) ? ( n1850 ) : ( n1855 ) ;
assign n1857 =  ( n1843 ) ? ( n1846 ) : ( n1856 ) ;
assign n1858 =  ( n1838 ) ? ( n1842 ) : ( n1857 ) ;
fun_PEActRelu  applyFunc_n1860(
    .arg0( n1858 ),
    .result( n1859 )
);
assign n1861 = n1859 ;
assign n1862 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n1863 =  ( bv_4_3_n166 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1864 = n1863 ;
assign n1866 = PE0_act_regs_3_data_n1865 ;
assign n1867 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1868 = n1863 ;
assign n1870 = PE0_act_regs_2_data_n1869 ;
assign n1871 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1872 = n1863 ;
assign n1874 = PE0_act_regs_1_data_n1873 ;
assign n1875 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1876 = n1863 ;
assign n1878 = PE0_act_regs_0_data_n1877 ;
assign n1879 =  ( n1875 ) ? ( n1878 ) : ( bv_20_0_n419 ) ;
assign n1880 =  ( n1871 ) ? ( n1874 ) : ( n1879 ) ;
assign n1881 =  ( n1867 ) ? ( n1870 ) : ( n1880 ) ;
assign n1882 =  ( n1862 ) ? ( n1866 ) : ( n1881 ) ;
fun_PEActOnex  applyFunc_n1884(
    .arg0( n1882 ),
    .result( n1883 )
);
assign n1885 = n1883 ;
assign n1886 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n1887 =  ( n1033 ) + ( bv_32_4_n380 )  ;
assign pe0_act_buffer_addr_n1888 = n1887 ;
assign n1890 = pe0_act_buffer_data_n1889 ;
fun_Adptfloat2Fixed  applyFunc_n1892(
    .arg0( n1890 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n1891 )
);
assign n1893 = n1891 ;
assign n1894 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n1895 =  ( bv_4_4_n176 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1896 = n1895 ;
assign n1898 = PE0_act_regs_3_data_n1897 ;
assign n1899 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1900 = n1895 ;
assign n1902 = PE0_act_regs_2_data_n1901 ;
assign n1903 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1904 = n1895 ;
assign n1906 = PE0_act_regs_1_data_n1905 ;
assign n1907 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1908 = n1895 ;
assign n1910 = PE0_act_regs_0_data_n1909 ;
assign n1911 =  ( n1907 ) ? ( n1910 ) : ( bv_20_0_n419 ) ;
assign n1912 =  ( n1903 ) ? ( n1906 ) : ( n1911 ) ;
assign n1913 =  ( n1899 ) ? ( n1902 ) : ( n1912 ) ;
assign n1914 =  ( n1894 ) ? ( n1898 ) : ( n1913 ) ;
assign n1915 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n1916 =  ( bv_4_4_n176 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1917 = n1916 ;
assign n1919 = PE0_act_regs_3_data_n1918 ;
assign n1920 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1921 = n1916 ;
assign n1923 = PE0_act_regs_2_data_n1922 ;
assign n1924 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1925 = n1916 ;
assign n1927 = PE0_act_regs_1_data_n1926 ;
assign n1928 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1929 = n1916 ;
assign n1931 = PE0_act_regs_0_data_n1930 ;
assign n1932 =  ( n1928 ) ? ( n1931 ) : ( bv_20_0_n419 ) ;
assign n1933 =  ( n1924 ) ? ( n1927 ) : ( n1932 ) ;
assign n1934 =  ( n1920 ) ? ( n1923 ) : ( n1933 ) ;
assign n1935 =  ( n1915 ) ? ( n1919 ) : ( n1934 ) ;
assign n1936 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n1937 = n1916 ;
assign n1939 = PE0_act_regs_3_data_n1938 ;
assign n1940 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1941 = n1916 ;
assign n1943 = PE0_act_regs_2_data_n1942 ;
assign n1944 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1945 = n1916 ;
assign n1947 = PE0_act_regs_1_data_n1946 ;
assign n1948 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1949 = n1916 ;
assign n1951 = PE0_act_regs_0_data_n1950 ;
assign n1952 =  ( n1948 ) ? ( n1951 ) : ( bv_20_0_n419 ) ;
assign n1953 =  ( n1944 ) ? ( n1947 ) : ( n1952 ) ;
assign n1954 =  ( n1940 ) ? ( n1943 ) : ( n1953 ) ;
assign n1955 =  ( n1936 ) ? ( n1939 ) : ( n1954 ) ;
fun_PEActEadd  applyFunc_n1957(
    .arg0( n1935 ),
    .arg1( n1955 ),
    .result( n1956 )
);
assign n1958 = n1956 ;
assign n1959 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n1960 =  ( bv_4_4_n176 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n1961 = n1960 ;
assign n1963 = PE0_act_regs_3_data_n1962 ;
assign n1964 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1965 = n1960 ;
assign n1967 = PE0_act_regs_2_data_n1966 ;
assign n1968 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1969 = n1960 ;
assign n1971 = PE0_act_regs_1_data_n1970 ;
assign n1972 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1973 = n1960 ;
assign n1975 = PE0_act_regs_0_data_n1974 ;
assign n1976 =  ( n1972 ) ? ( n1975 ) : ( bv_20_0_n419 ) ;
assign n1977 =  ( n1968 ) ? ( n1971 ) : ( n1976 ) ;
assign n1978 =  ( n1964 ) ? ( n1967 ) : ( n1977 ) ;
assign n1979 =  ( n1959 ) ? ( n1963 ) : ( n1978 ) ;
assign n1980 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n1981 = n1960 ;
assign n1983 = PE0_act_regs_3_data_n1982 ;
assign n1984 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n1985 = n1960 ;
assign n1987 = PE0_act_regs_2_data_n1986 ;
assign n1988 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n1989 = n1960 ;
assign n1991 = PE0_act_regs_1_data_n1990 ;
assign n1992 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n1993 = n1960 ;
assign n1995 = PE0_act_regs_0_data_n1994 ;
assign n1996 =  ( n1992 ) ? ( n1995 ) : ( bv_20_0_n419 ) ;
assign n1997 =  ( n1988 ) ? ( n1991 ) : ( n1996 ) ;
assign n1998 =  ( n1984 ) ? ( n1987 ) : ( n1997 ) ;
assign n1999 =  ( n1980 ) ? ( n1983 ) : ( n1998 ) ;
fun_PEActEmul  applyFunc_n2001(
    .arg0( n1979 ),
    .arg1( n1999 ),
    .result( n2000 )
);
assign n2002 = n2000 ;
assign n2003 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n2004 =  ( bv_4_4_n176 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2005 = n2004 ;
assign n2007 = PE0_act_regs_3_data_n2006 ;
assign n2008 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2009 = n2004 ;
assign n2011 = PE0_act_regs_2_data_n2010 ;
assign n2012 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2013 = n2004 ;
assign n2015 = PE0_act_regs_1_data_n2014 ;
assign n2016 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2017 = n2004 ;
assign n2019 = PE0_act_regs_0_data_n2018 ;
assign n2020 =  ( n2016 ) ? ( n2019 ) : ( bv_20_0_n419 ) ;
assign n2021 =  ( n2012 ) ? ( n2015 ) : ( n2020 ) ;
assign n2022 =  ( n2008 ) ? ( n2011 ) : ( n2021 ) ;
assign n2023 =  ( n2003 ) ? ( n2007 ) : ( n2022 ) ;
fun_PEActSigmoid  applyFunc_n2025(
    .arg0( n2023 ),
    .result( n2024 )
);
assign n2026 = n2024 ;
assign n2027 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n2028 =  ( bv_4_4_n176 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2029 = n2028 ;
assign n2031 = PE0_act_regs_3_data_n2030 ;
assign n2032 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2033 = n2028 ;
assign n2035 = PE0_act_regs_2_data_n2034 ;
assign n2036 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2037 = n2028 ;
assign n2039 = PE0_act_regs_1_data_n2038 ;
assign n2040 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2041 = n2028 ;
assign n2043 = PE0_act_regs_0_data_n2042 ;
assign n2044 =  ( n2040 ) ? ( n2043 ) : ( bv_20_0_n419 ) ;
assign n2045 =  ( n2036 ) ? ( n2039 ) : ( n2044 ) ;
assign n2046 =  ( n2032 ) ? ( n2035 ) : ( n2045 ) ;
assign n2047 =  ( n2027 ) ? ( n2031 ) : ( n2046 ) ;
fun_PEActTanh  applyFunc_n2049(
    .arg0( n2047 ),
    .result( n2048 )
);
assign n2050 = n2048 ;
assign n2051 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n2052 =  ( bv_4_4_n176 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2053 = n2052 ;
assign n2055 = PE0_act_regs_3_data_n2054 ;
assign n2056 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2057 = n2052 ;
assign n2059 = PE0_act_regs_2_data_n2058 ;
assign n2060 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2061 = n2052 ;
assign n2063 = PE0_act_regs_1_data_n2062 ;
assign n2064 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2065 = n2052 ;
assign n2067 = PE0_act_regs_0_data_n2066 ;
assign n2068 =  ( n2064 ) ? ( n2067 ) : ( bv_20_0_n419 ) ;
assign n2069 =  ( n2060 ) ? ( n2063 ) : ( n2068 ) ;
assign n2070 =  ( n2056 ) ? ( n2059 ) : ( n2069 ) ;
assign n2071 =  ( n2051 ) ? ( n2055 ) : ( n2070 ) ;
fun_PEActRelu  applyFunc_n2073(
    .arg0( n2071 ),
    .result( n2072 )
);
assign n2074 = n2072 ;
assign n2075 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n2076 =  ( bv_4_4_n176 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2077 = n2076 ;
assign n2079 = PE0_act_regs_3_data_n2078 ;
assign n2080 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2081 = n2076 ;
assign n2083 = PE0_act_regs_2_data_n2082 ;
assign n2084 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2085 = n2076 ;
assign n2087 = PE0_act_regs_1_data_n2086 ;
assign n2088 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2089 = n2076 ;
assign n2091 = PE0_act_regs_0_data_n2090 ;
assign n2092 =  ( n2088 ) ? ( n2091 ) : ( bv_20_0_n419 ) ;
assign n2093 =  ( n2084 ) ? ( n2087 ) : ( n2092 ) ;
assign n2094 =  ( n2080 ) ? ( n2083 ) : ( n2093 ) ;
assign n2095 =  ( n2075 ) ? ( n2079 ) : ( n2094 ) ;
fun_PEActOnex  applyFunc_n2097(
    .arg0( n2095 ),
    .result( n2096 )
);
assign n2098 = n2096 ;
assign n2099 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n2100 =  ( n1033 ) + ( bv_32_5_n378 )  ;
assign pe0_act_buffer_addr_n2101 = n2100 ;
assign n2103 = pe0_act_buffer_data_n2102 ;
fun_Adptfloat2Fixed  applyFunc_n2105(
    .arg0( n2103 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n2104 )
);
assign n2106 = n2104 ;
assign n2107 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n2108 =  ( bv_4_5_n656 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2109 = n2108 ;
assign n2111 = PE0_act_regs_3_data_n2110 ;
assign n2112 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2113 = n2108 ;
assign n2115 = PE0_act_regs_2_data_n2114 ;
assign n2116 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2117 = n2108 ;
assign n2119 = PE0_act_regs_1_data_n2118 ;
assign n2120 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2121 = n2108 ;
assign n2123 = PE0_act_regs_0_data_n2122 ;
assign n2124 =  ( n2120 ) ? ( n2123 ) : ( bv_20_0_n419 ) ;
assign n2125 =  ( n2116 ) ? ( n2119 ) : ( n2124 ) ;
assign n2126 =  ( n2112 ) ? ( n2115 ) : ( n2125 ) ;
assign n2127 =  ( n2107 ) ? ( n2111 ) : ( n2126 ) ;
assign n2128 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n2129 =  ( bv_4_5_n656 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2130 = n2129 ;
assign n2132 = PE0_act_regs_3_data_n2131 ;
assign n2133 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2134 = n2129 ;
assign n2136 = PE0_act_regs_2_data_n2135 ;
assign n2137 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2138 = n2129 ;
assign n2140 = PE0_act_regs_1_data_n2139 ;
assign n2141 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2142 = n2129 ;
assign n2144 = PE0_act_regs_0_data_n2143 ;
assign n2145 =  ( n2141 ) ? ( n2144 ) : ( bv_20_0_n419 ) ;
assign n2146 =  ( n2137 ) ? ( n2140 ) : ( n2145 ) ;
assign n2147 =  ( n2133 ) ? ( n2136 ) : ( n2146 ) ;
assign n2148 =  ( n2128 ) ? ( n2132 ) : ( n2147 ) ;
assign n2149 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n2150 = n2129 ;
assign n2152 = PE0_act_regs_3_data_n2151 ;
assign n2153 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2154 = n2129 ;
assign n2156 = PE0_act_regs_2_data_n2155 ;
assign n2157 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2158 = n2129 ;
assign n2160 = PE0_act_regs_1_data_n2159 ;
assign n2161 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2162 = n2129 ;
assign n2164 = PE0_act_regs_0_data_n2163 ;
assign n2165 =  ( n2161 ) ? ( n2164 ) : ( bv_20_0_n419 ) ;
assign n2166 =  ( n2157 ) ? ( n2160 ) : ( n2165 ) ;
assign n2167 =  ( n2153 ) ? ( n2156 ) : ( n2166 ) ;
assign n2168 =  ( n2149 ) ? ( n2152 ) : ( n2167 ) ;
fun_PEActEadd  applyFunc_n2170(
    .arg0( n2148 ),
    .arg1( n2168 ),
    .result( n2169 )
);
assign n2171 = n2169 ;
assign n2172 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n2173 =  ( bv_4_5_n656 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2174 = n2173 ;
assign n2176 = PE0_act_regs_3_data_n2175 ;
assign n2177 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2178 = n2173 ;
assign n2180 = PE0_act_regs_2_data_n2179 ;
assign n2181 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2182 = n2173 ;
assign n2184 = PE0_act_regs_1_data_n2183 ;
assign n2185 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2186 = n2173 ;
assign n2188 = PE0_act_regs_0_data_n2187 ;
assign n2189 =  ( n2185 ) ? ( n2188 ) : ( bv_20_0_n419 ) ;
assign n2190 =  ( n2181 ) ? ( n2184 ) : ( n2189 ) ;
assign n2191 =  ( n2177 ) ? ( n2180 ) : ( n2190 ) ;
assign n2192 =  ( n2172 ) ? ( n2176 ) : ( n2191 ) ;
assign n2193 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n2194 = n2173 ;
assign n2196 = PE0_act_regs_3_data_n2195 ;
assign n2197 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2198 = n2173 ;
assign n2200 = PE0_act_regs_2_data_n2199 ;
assign n2201 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2202 = n2173 ;
assign n2204 = PE0_act_regs_1_data_n2203 ;
assign n2205 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2206 = n2173 ;
assign n2208 = PE0_act_regs_0_data_n2207 ;
assign n2209 =  ( n2205 ) ? ( n2208 ) : ( bv_20_0_n419 ) ;
assign n2210 =  ( n2201 ) ? ( n2204 ) : ( n2209 ) ;
assign n2211 =  ( n2197 ) ? ( n2200 ) : ( n2210 ) ;
assign n2212 =  ( n2193 ) ? ( n2196 ) : ( n2211 ) ;
fun_PEActEmul  applyFunc_n2214(
    .arg0( n2192 ),
    .arg1( n2212 ),
    .result( n2213 )
);
assign n2215 = n2213 ;
assign n2216 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n2217 =  ( bv_4_5_n656 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2218 = n2217 ;
assign n2220 = PE0_act_regs_3_data_n2219 ;
assign n2221 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2222 = n2217 ;
assign n2224 = PE0_act_regs_2_data_n2223 ;
assign n2225 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2226 = n2217 ;
assign n2228 = PE0_act_regs_1_data_n2227 ;
assign n2229 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2230 = n2217 ;
assign n2232 = PE0_act_regs_0_data_n2231 ;
assign n2233 =  ( n2229 ) ? ( n2232 ) : ( bv_20_0_n419 ) ;
assign n2234 =  ( n2225 ) ? ( n2228 ) : ( n2233 ) ;
assign n2235 =  ( n2221 ) ? ( n2224 ) : ( n2234 ) ;
assign n2236 =  ( n2216 ) ? ( n2220 ) : ( n2235 ) ;
fun_PEActSigmoid  applyFunc_n2238(
    .arg0( n2236 ),
    .result( n2237 )
);
assign n2239 = n2237 ;
assign n2240 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n2241 =  ( bv_4_5_n656 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2242 = n2241 ;
assign n2244 = PE0_act_regs_3_data_n2243 ;
assign n2245 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2246 = n2241 ;
assign n2248 = PE0_act_regs_2_data_n2247 ;
assign n2249 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2250 = n2241 ;
assign n2252 = PE0_act_regs_1_data_n2251 ;
assign n2253 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2254 = n2241 ;
assign n2256 = PE0_act_regs_0_data_n2255 ;
assign n2257 =  ( n2253 ) ? ( n2256 ) : ( bv_20_0_n419 ) ;
assign n2258 =  ( n2249 ) ? ( n2252 ) : ( n2257 ) ;
assign n2259 =  ( n2245 ) ? ( n2248 ) : ( n2258 ) ;
assign n2260 =  ( n2240 ) ? ( n2244 ) : ( n2259 ) ;
fun_PEActTanh  applyFunc_n2262(
    .arg0( n2260 ),
    .result( n2261 )
);
assign n2263 = n2261 ;
assign n2264 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n2265 =  ( bv_4_5_n656 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2266 = n2265 ;
assign n2268 = PE0_act_regs_3_data_n2267 ;
assign n2269 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2270 = n2265 ;
assign n2272 = PE0_act_regs_2_data_n2271 ;
assign n2273 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2274 = n2265 ;
assign n2276 = PE0_act_regs_1_data_n2275 ;
assign n2277 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2278 = n2265 ;
assign n2280 = PE0_act_regs_0_data_n2279 ;
assign n2281 =  ( n2277 ) ? ( n2280 ) : ( bv_20_0_n419 ) ;
assign n2282 =  ( n2273 ) ? ( n2276 ) : ( n2281 ) ;
assign n2283 =  ( n2269 ) ? ( n2272 ) : ( n2282 ) ;
assign n2284 =  ( n2264 ) ? ( n2268 ) : ( n2283 ) ;
fun_PEActRelu  applyFunc_n2286(
    .arg0( n2284 ),
    .result( n2285 )
);
assign n2287 = n2285 ;
assign n2288 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n2289 =  ( bv_4_5_n656 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2290 = n2289 ;
assign n2292 = PE0_act_regs_3_data_n2291 ;
assign n2293 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2294 = n2289 ;
assign n2296 = PE0_act_regs_2_data_n2295 ;
assign n2297 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2298 = n2289 ;
assign n2300 = PE0_act_regs_1_data_n2299 ;
assign n2301 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2302 = n2289 ;
assign n2304 = PE0_act_regs_0_data_n2303 ;
assign n2305 =  ( n2301 ) ? ( n2304 ) : ( bv_20_0_n419 ) ;
assign n2306 =  ( n2297 ) ? ( n2300 ) : ( n2305 ) ;
assign n2307 =  ( n2293 ) ? ( n2296 ) : ( n2306 ) ;
assign n2308 =  ( n2288 ) ? ( n2292 ) : ( n2307 ) ;
fun_PEActOnex  applyFunc_n2310(
    .arg0( n2308 ),
    .result( n2309 )
);
assign n2311 = n2309 ;
assign n2312 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n2313 =  ( n1033 ) + ( bv_32_6_n376 )  ;
assign pe0_act_buffer_addr_n2314 = n2313 ;
assign n2316 = pe0_act_buffer_data_n2315 ;
fun_Adptfloat2Fixed  applyFunc_n2318(
    .arg0( n2316 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n2317 )
);
assign n2319 = n2317 ;
assign n2320 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n2321 =  ( bv_4_6_n630 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2322 = n2321 ;
assign n2324 = PE0_act_regs_3_data_n2323 ;
assign n2325 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2326 = n2321 ;
assign n2328 = PE0_act_regs_2_data_n2327 ;
assign n2329 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2330 = n2321 ;
assign n2332 = PE0_act_regs_1_data_n2331 ;
assign n2333 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2334 = n2321 ;
assign n2336 = PE0_act_regs_0_data_n2335 ;
assign n2337 =  ( n2333 ) ? ( n2336 ) : ( bv_20_0_n419 ) ;
assign n2338 =  ( n2329 ) ? ( n2332 ) : ( n2337 ) ;
assign n2339 =  ( n2325 ) ? ( n2328 ) : ( n2338 ) ;
assign n2340 =  ( n2320 ) ? ( n2324 ) : ( n2339 ) ;
assign n2341 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n2342 =  ( bv_4_6_n630 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2343 = n2342 ;
assign n2345 = PE0_act_regs_3_data_n2344 ;
assign n2346 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2347 = n2342 ;
assign n2349 = PE0_act_regs_2_data_n2348 ;
assign n2350 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2351 = n2342 ;
assign n2353 = PE0_act_regs_1_data_n2352 ;
assign n2354 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2355 = n2342 ;
assign n2357 = PE0_act_regs_0_data_n2356 ;
assign n2358 =  ( n2354 ) ? ( n2357 ) : ( bv_20_0_n419 ) ;
assign n2359 =  ( n2350 ) ? ( n2353 ) : ( n2358 ) ;
assign n2360 =  ( n2346 ) ? ( n2349 ) : ( n2359 ) ;
assign n2361 =  ( n2341 ) ? ( n2345 ) : ( n2360 ) ;
assign n2362 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n2363 = n2342 ;
assign n2365 = PE0_act_regs_3_data_n2364 ;
assign n2366 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2367 = n2342 ;
assign n2369 = PE0_act_regs_2_data_n2368 ;
assign n2370 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2371 = n2342 ;
assign n2373 = PE0_act_regs_1_data_n2372 ;
assign n2374 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2375 = n2342 ;
assign n2377 = PE0_act_regs_0_data_n2376 ;
assign n2378 =  ( n2374 ) ? ( n2377 ) : ( bv_20_0_n419 ) ;
assign n2379 =  ( n2370 ) ? ( n2373 ) : ( n2378 ) ;
assign n2380 =  ( n2366 ) ? ( n2369 ) : ( n2379 ) ;
assign n2381 =  ( n2362 ) ? ( n2365 ) : ( n2380 ) ;
fun_PEActEadd  applyFunc_n2383(
    .arg0( n2361 ),
    .arg1( n2381 ),
    .result( n2382 )
);
assign n2384 = n2382 ;
assign n2385 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n2386 =  ( bv_4_6_n630 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2387 = n2386 ;
assign n2389 = PE0_act_regs_3_data_n2388 ;
assign n2390 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2391 = n2386 ;
assign n2393 = PE0_act_regs_2_data_n2392 ;
assign n2394 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2395 = n2386 ;
assign n2397 = PE0_act_regs_1_data_n2396 ;
assign n2398 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2399 = n2386 ;
assign n2401 = PE0_act_regs_0_data_n2400 ;
assign n2402 =  ( n2398 ) ? ( n2401 ) : ( bv_20_0_n419 ) ;
assign n2403 =  ( n2394 ) ? ( n2397 ) : ( n2402 ) ;
assign n2404 =  ( n2390 ) ? ( n2393 ) : ( n2403 ) ;
assign n2405 =  ( n2385 ) ? ( n2389 ) : ( n2404 ) ;
assign n2406 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n2407 = n2386 ;
assign n2409 = PE0_act_regs_3_data_n2408 ;
assign n2410 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2411 = n2386 ;
assign n2413 = PE0_act_regs_2_data_n2412 ;
assign n2414 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2415 = n2386 ;
assign n2417 = PE0_act_regs_1_data_n2416 ;
assign n2418 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2419 = n2386 ;
assign n2421 = PE0_act_regs_0_data_n2420 ;
assign n2422 =  ( n2418 ) ? ( n2421 ) : ( bv_20_0_n419 ) ;
assign n2423 =  ( n2414 ) ? ( n2417 ) : ( n2422 ) ;
assign n2424 =  ( n2410 ) ? ( n2413 ) : ( n2423 ) ;
assign n2425 =  ( n2406 ) ? ( n2409 ) : ( n2424 ) ;
fun_PEActEmul  applyFunc_n2427(
    .arg0( n2405 ),
    .arg1( n2425 ),
    .result( n2426 )
);
assign n2428 = n2426 ;
assign n2429 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n2430 =  ( bv_4_6_n630 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2431 = n2430 ;
assign n2433 = PE0_act_regs_3_data_n2432 ;
assign n2434 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2435 = n2430 ;
assign n2437 = PE0_act_regs_2_data_n2436 ;
assign n2438 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2439 = n2430 ;
assign n2441 = PE0_act_regs_1_data_n2440 ;
assign n2442 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2443 = n2430 ;
assign n2445 = PE0_act_regs_0_data_n2444 ;
assign n2446 =  ( n2442 ) ? ( n2445 ) : ( bv_20_0_n419 ) ;
assign n2447 =  ( n2438 ) ? ( n2441 ) : ( n2446 ) ;
assign n2448 =  ( n2434 ) ? ( n2437 ) : ( n2447 ) ;
assign n2449 =  ( n2429 ) ? ( n2433 ) : ( n2448 ) ;
fun_PEActSigmoid  applyFunc_n2451(
    .arg0( n2449 ),
    .result( n2450 )
);
assign n2452 = n2450 ;
assign n2453 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n2454 =  ( bv_4_6_n630 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2455 = n2454 ;
assign n2457 = PE0_act_regs_3_data_n2456 ;
assign n2458 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2459 = n2454 ;
assign n2461 = PE0_act_regs_2_data_n2460 ;
assign n2462 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2463 = n2454 ;
assign n2465 = PE0_act_regs_1_data_n2464 ;
assign n2466 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2467 = n2454 ;
assign n2469 = PE0_act_regs_0_data_n2468 ;
assign n2470 =  ( n2466 ) ? ( n2469 ) : ( bv_20_0_n419 ) ;
assign n2471 =  ( n2462 ) ? ( n2465 ) : ( n2470 ) ;
assign n2472 =  ( n2458 ) ? ( n2461 ) : ( n2471 ) ;
assign n2473 =  ( n2453 ) ? ( n2457 ) : ( n2472 ) ;
fun_PEActTanh  applyFunc_n2475(
    .arg0( n2473 ),
    .result( n2474 )
);
assign n2476 = n2474 ;
assign n2477 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n2478 =  ( bv_4_6_n630 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2479 = n2478 ;
assign n2481 = PE0_act_regs_3_data_n2480 ;
assign n2482 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2483 = n2478 ;
assign n2485 = PE0_act_regs_2_data_n2484 ;
assign n2486 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2487 = n2478 ;
assign n2489 = PE0_act_regs_1_data_n2488 ;
assign n2490 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2491 = n2478 ;
assign n2493 = PE0_act_regs_0_data_n2492 ;
assign n2494 =  ( n2490 ) ? ( n2493 ) : ( bv_20_0_n419 ) ;
assign n2495 =  ( n2486 ) ? ( n2489 ) : ( n2494 ) ;
assign n2496 =  ( n2482 ) ? ( n2485 ) : ( n2495 ) ;
assign n2497 =  ( n2477 ) ? ( n2481 ) : ( n2496 ) ;
fun_PEActRelu  applyFunc_n2499(
    .arg0( n2497 ),
    .result( n2498 )
);
assign n2500 = n2498 ;
assign n2501 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n2502 =  ( bv_4_6_n630 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2503 = n2502 ;
assign n2505 = PE0_act_regs_3_data_n2504 ;
assign n2506 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2507 = n2502 ;
assign n2509 = PE0_act_regs_2_data_n2508 ;
assign n2510 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2511 = n2502 ;
assign n2513 = PE0_act_regs_1_data_n2512 ;
assign n2514 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2515 = n2502 ;
assign n2517 = PE0_act_regs_0_data_n2516 ;
assign n2518 =  ( n2514 ) ? ( n2517 ) : ( bv_20_0_n419 ) ;
assign n2519 =  ( n2510 ) ? ( n2513 ) : ( n2518 ) ;
assign n2520 =  ( n2506 ) ? ( n2509 ) : ( n2519 ) ;
assign n2521 =  ( n2501 ) ? ( n2505 ) : ( n2520 ) ;
fun_PEActOnex  applyFunc_n2523(
    .arg0( n2521 ),
    .result( n2522 )
);
assign n2524 = n2522 ;
assign n2525 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n2526 =  ( n1033 ) + ( bv_32_7_n374 )  ;
assign pe0_act_buffer_addr_n2527 = n2526 ;
assign n2529 = pe0_act_buffer_data_n2528 ;
fun_Adptfloat2Fixed  applyFunc_n2531(
    .arg0( n2529 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n2530 )
);
assign n2532 = n2530 ;
assign n2533 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n2534 =  ( bv_4_7_n184 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2535 = n2534 ;
assign n2537 = PE0_act_regs_3_data_n2536 ;
assign n2538 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2539 = n2534 ;
assign n2541 = PE0_act_regs_2_data_n2540 ;
assign n2542 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2543 = n2534 ;
assign n2545 = PE0_act_regs_1_data_n2544 ;
assign n2546 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2547 = n2534 ;
assign n2549 = PE0_act_regs_0_data_n2548 ;
assign n2550 =  ( n2546 ) ? ( n2549 ) : ( bv_20_0_n419 ) ;
assign n2551 =  ( n2542 ) ? ( n2545 ) : ( n2550 ) ;
assign n2552 =  ( n2538 ) ? ( n2541 ) : ( n2551 ) ;
assign n2553 =  ( n2533 ) ? ( n2537 ) : ( n2552 ) ;
assign n2554 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n2555 =  ( bv_4_7_n184 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2556 = n2555 ;
assign n2558 = PE0_act_regs_3_data_n2557 ;
assign n2559 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2560 = n2555 ;
assign n2562 = PE0_act_regs_2_data_n2561 ;
assign n2563 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2564 = n2555 ;
assign n2566 = PE0_act_regs_1_data_n2565 ;
assign n2567 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2568 = n2555 ;
assign n2570 = PE0_act_regs_0_data_n2569 ;
assign n2571 =  ( n2567 ) ? ( n2570 ) : ( bv_20_0_n419 ) ;
assign n2572 =  ( n2563 ) ? ( n2566 ) : ( n2571 ) ;
assign n2573 =  ( n2559 ) ? ( n2562 ) : ( n2572 ) ;
assign n2574 =  ( n2554 ) ? ( n2558 ) : ( n2573 ) ;
assign n2575 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n2576 = n2555 ;
assign n2578 = PE0_act_regs_3_data_n2577 ;
assign n2579 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2580 = n2555 ;
assign n2582 = PE0_act_regs_2_data_n2581 ;
assign n2583 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2584 = n2555 ;
assign n2586 = PE0_act_regs_1_data_n2585 ;
assign n2587 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2588 = n2555 ;
assign n2590 = PE0_act_regs_0_data_n2589 ;
assign n2591 =  ( n2587 ) ? ( n2590 ) : ( bv_20_0_n419 ) ;
assign n2592 =  ( n2583 ) ? ( n2586 ) : ( n2591 ) ;
assign n2593 =  ( n2579 ) ? ( n2582 ) : ( n2592 ) ;
assign n2594 =  ( n2575 ) ? ( n2578 ) : ( n2593 ) ;
fun_PEActEadd  applyFunc_n2596(
    .arg0( n2574 ),
    .arg1( n2594 ),
    .result( n2595 )
);
assign n2597 = n2595 ;
assign n2598 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n2599 =  ( bv_4_7_n184 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2600 = n2599 ;
assign n2602 = PE0_act_regs_3_data_n2601 ;
assign n2603 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2604 = n2599 ;
assign n2606 = PE0_act_regs_2_data_n2605 ;
assign n2607 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2608 = n2599 ;
assign n2610 = PE0_act_regs_1_data_n2609 ;
assign n2611 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2612 = n2599 ;
assign n2614 = PE0_act_regs_0_data_n2613 ;
assign n2615 =  ( n2611 ) ? ( n2614 ) : ( bv_20_0_n419 ) ;
assign n2616 =  ( n2607 ) ? ( n2610 ) : ( n2615 ) ;
assign n2617 =  ( n2603 ) ? ( n2606 ) : ( n2616 ) ;
assign n2618 =  ( n2598 ) ? ( n2602 ) : ( n2617 ) ;
assign n2619 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n2620 = n2599 ;
assign n2622 = PE0_act_regs_3_data_n2621 ;
assign n2623 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2624 = n2599 ;
assign n2626 = PE0_act_regs_2_data_n2625 ;
assign n2627 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2628 = n2599 ;
assign n2630 = PE0_act_regs_1_data_n2629 ;
assign n2631 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2632 = n2599 ;
assign n2634 = PE0_act_regs_0_data_n2633 ;
assign n2635 =  ( n2631 ) ? ( n2634 ) : ( bv_20_0_n419 ) ;
assign n2636 =  ( n2627 ) ? ( n2630 ) : ( n2635 ) ;
assign n2637 =  ( n2623 ) ? ( n2626 ) : ( n2636 ) ;
assign n2638 =  ( n2619 ) ? ( n2622 ) : ( n2637 ) ;
fun_PEActEmul  applyFunc_n2640(
    .arg0( n2618 ),
    .arg1( n2638 ),
    .result( n2639 )
);
assign n2641 = n2639 ;
assign n2642 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n2643 =  ( bv_4_7_n184 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2644 = n2643 ;
assign n2646 = PE0_act_regs_3_data_n2645 ;
assign n2647 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2648 = n2643 ;
assign n2650 = PE0_act_regs_2_data_n2649 ;
assign n2651 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2652 = n2643 ;
assign n2654 = PE0_act_regs_1_data_n2653 ;
assign n2655 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2656 = n2643 ;
assign n2658 = PE0_act_regs_0_data_n2657 ;
assign n2659 =  ( n2655 ) ? ( n2658 ) : ( bv_20_0_n419 ) ;
assign n2660 =  ( n2651 ) ? ( n2654 ) : ( n2659 ) ;
assign n2661 =  ( n2647 ) ? ( n2650 ) : ( n2660 ) ;
assign n2662 =  ( n2642 ) ? ( n2646 ) : ( n2661 ) ;
fun_PEActSigmoid  applyFunc_n2664(
    .arg0( n2662 ),
    .result( n2663 )
);
assign n2665 = n2663 ;
assign n2666 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n2667 =  ( bv_4_7_n184 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2668 = n2667 ;
assign n2670 = PE0_act_regs_3_data_n2669 ;
assign n2671 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2672 = n2667 ;
assign n2674 = PE0_act_regs_2_data_n2673 ;
assign n2675 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2676 = n2667 ;
assign n2678 = PE0_act_regs_1_data_n2677 ;
assign n2679 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2680 = n2667 ;
assign n2682 = PE0_act_regs_0_data_n2681 ;
assign n2683 =  ( n2679 ) ? ( n2682 ) : ( bv_20_0_n419 ) ;
assign n2684 =  ( n2675 ) ? ( n2678 ) : ( n2683 ) ;
assign n2685 =  ( n2671 ) ? ( n2674 ) : ( n2684 ) ;
assign n2686 =  ( n2666 ) ? ( n2670 ) : ( n2685 ) ;
fun_PEActTanh  applyFunc_n2688(
    .arg0( n2686 ),
    .result( n2687 )
);
assign n2689 = n2687 ;
assign n2690 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n2691 =  ( bv_4_7_n184 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2692 = n2691 ;
assign n2694 = PE0_act_regs_3_data_n2693 ;
assign n2695 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2696 = n2691 ;
assign n2698 = PE0_act_regs_2_data_n2697 ;
assign n2699 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2700 = n2691 ;
assign n2702 = PE0_act_regs_1_data_n2701 ;
assign n2703 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2704 = n2691 ;
assign n2706 = PE0_act_regs_0_data_n2705 ;
assign n2707 =  ( n2703 ) ? ( n2706 ) : ( bv_20_0_n419 ) ;
assign n2708 =  ( n2699 ) ? ( n2702 ) : ( n2707 ) ;
assign n2709 =  ( n2695 ) ? ( n2698 ) : ( n2708 ) ;
assign n2710 =  ( n2690 ) ? ( n2694 ) : ( n2709 ) ;
fun_PEActRelu  applyFunc_n2712(
    .arg0( n2710 ),
    .result( n2711 )
);
assign n2713 = n2711 ;
assign n2714 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n2715 =  ( bv_4_7_n184 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2716 = n2715 ;
assign n2718 = PE0_act_regs_3_data_n2717 ;
assign n2719 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2720 = n2715 ;
assign n2722 = PE0_act_regs_2_data_n2721 ;
assign n2723 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2724 = n2715 ;
assign n2726 = PE0_act_regs_1_data_n2725 ;
assign n2727 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2728 = n2715 ;
assign n2730 = PE0_act_regs_0_data_n2729 ;
assign n2731 =  ( n2727 ) ? ( n2730 ) : ( bv_20_0_n419 ) ;
assign n2732 =  ( n2723 ) ? ( n2726 ) : ( n2731 ) ;
assign n2733 =  ( n2719 ) ? ( n2722 ) : ( n2732 ) ;
assign n2734 =  ( n2714 ) ? ( n2718 ) : ( n2733 ) ;
fun_PEActOnex  applyFunc_n2736(
    .arg0( n2734 ),
    .result( n2735 )
);
assign n2737 = n2735 ;
assign n2738 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n2739 =  ( n1033 ) + ( bv_32_8_n372 )  ;
assign pe0_act_buffer_addr_n2740 = n2739 ;
assign n2742 = pe0_act_buffer_data_n2741 ;
fun_Adptfloat2Fixed  applyFunc_n2744(
    .arg0( n2742 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n2743 )
);
assign n2745 = n2743 ;
assign n2746 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n2747 =  ( bv_4_8_n190 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2748 = n2747 ;
assign n2750 = PE0_act_regs_3_data_n2749 ;
assign n2751 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2752 = n2747 ;
assign n2754 = PE0_act_regs_2_data_n2753 ;
assign n2755 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2756 = n2747 ;
assign n2758 = PE0_act_regs_1_data_n2757 ;
assign n2759 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2760 = n2747 ;
assign n2762 = PE0_act_regs_0_data_n2761 ;
assign n2763 =  ( n2759 ) ? ( n2762 ) : ( bv_20_0_n419 ) ;
assign n2764 =  ( n2755 ) ? ( n2758 ) : ( n2763 ) ;
assign n2765 =  ( n2751 ) ? ( n2754 ) : ( n2764 ) ;
assign n2766 =  ( n2746 ) ? ( n2750 ) : ( n2765 ) ;
assign n2767 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n2768 =  ( bv_4_8_n190 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2769 = n2768 ;
assign n2771 = PE0_act_regs_3_data_n2770 ;
assign n2772 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2773 = n2768 ;
assign n2775 = PE0_act_regs_2_data_n2774 ;
assign n2776 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2777 = n2768 ;
assign n2779 = PE0_act_regs_1_data_n2778 ;
assign n2780 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2781 = n2768 ;
assign n2783 = PE0_act_regs_0_data_n2782 ;
assign n2784 =  ( n2780 ) ? ( n2783 ) : ( bv_20_0_n419 ) ;
assign n2785 =  ( n2776 ) ? ( n2779 ) : ( n2784 ) ;
assign n2786 =  ( n2772 ) ? ( n2775 ) : ( n2785 ) ;
assign n2787 =  ( n2767 ) ? ( n2771 ) : ( n2786 ) ;
assign n2788 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n2789 = n2768 ;
assign n2791 = PE0_act_regs_3_data_n2790 ;
assign n2792 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2793 = n2768 ;
assign n2795 = PE0_act_regs_2_data_n2794 ;
assign n2796 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2797 = n2768 ;
assign n2799 = PE0_act_regs_1_data_n2798 ;
assign n2800 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2801 = n2768 ;
assign n2803 = PE0_act_regs_0_data_n2802 ;
assign n2804 =  ( n2800 ) ? ( n2803 ) : ( bv_20_0_n419 ) ;
assign n2805 =  ( n2796 ) ? ( n2799 ) : ( n2804 ) ;
assign n2806 =  ( n2792 ) ? ( n2795 ) : ( n2805 ) ;
assign n2807 =  ( n2788 ) ? ( n2791 ) : ( n2806 ) ;
fun_PEActEadd  applyFunc_n2809(
    .arg0( n2787 ),
    .arg1( n2807 ),
    .result( n2808 )
);
assign n2810 = n2808 ;
assign n2811 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n2812 =  ( bv_4_8_n190 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2813 = n2812 ;
assign n2815 = PE0_act_regs_3_data_n2814 ;
assign n2816 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2817 = n2812 ;
assign n2819 = PE0_act_regs_2_data_n2818 ;
assign n2820 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2821 = n2812 ;
assign n2823 = PE0_act_regs_1_data_n2822 ;
assign n2824 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2825 = n2812 ;
assign n2827 = PE0_act_regs_0_data_n2826 ;
assign n2828 =  ( n2824 ) ? ( n2827 ) : ( bv_20_0_n419 ) ;
assign n2829 =  ( n2820 ) ? ( n2823 ) : ( n2828 ) ;
assign n2830 =  ( n2816 ) ? ( n2819 ) : ( n2829 ) ;
assign n2831 =  ( n2811 ) ? ( n2815 ) : ( n2830 ) ;
assign n2832 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n2833 = n2812 ;
assign n2835 = PE0_act_regs_3_data_n2834 ;
assign n2836 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2837 = n2812 ;
assign n2839 = PE0_act_regs_2_data_n2838 ;
assign n2840 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2841 = n2812 ;
assign n2843 = PE0_act_regs_1_data_n2842 ;
assign n2844 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2845 = n2812 ;
assign n2847 = PE0_act_regs_0_data_n2846 ;
assign n2848 =  ( n2844 ) ? ( n2847 ) : ( bv_20_0_n419 ) ;
assign n2849 =  ( n2840 ) ? ( n2843 ) : ( n2848 ) ;
assign n2850 =  ( n2836 ) ? ( n2839 ) : ( n2849 ) ;
assign n2851 =  ( n2832 ) ? ( n2835 ) : ( n2850 ) ;
fun_PEActEmul  applyFunc_n2853(
    .arg0( n2831 ),
    .arg1( n2851 ),
    .result( n2852 )
);
assign n2854 = n2852 ;
assign n2855 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n2856 =  ( bv_4_8_n190 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2857 = n2856 ;
assign n2859 = PE0_act_regs_3_data_n2858 ;
assign n2860 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2861 = n2856 ;
assign n2863 = PE0_act_regs_2_data_n2862 ;
assign n2864 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2865 = n2856 ;
assign n2867 = PE0_act_regs_1_data_n2866 ;
assign n2868 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2869 = n2856 ;
assign n2871 = PE0_act_regs_0_data_n2870 ;
assign n2872 =  ( n2868 ) ? ( n2871 ) : ( bv_20_0_n419 ) ;
assign n2873 =  ( n2864 ) ? ( n2867 ) : ( n2872 ) ;
assign n2874 =  ( n2860 ) ? ( n2863 ) : ( n2873 ) ;
assign n2875 =  ( n2855 ) ? ( n2859 ) : ( n2874 ) ;
fun_PEActSigmoid  applyFunc_n2877(
    .arg0( n2875 ),
    .result( n2876 )
);
assign n2878 = n2876 ;
assign n2879 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n2880 =  ( bv_4_8_n190 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2881 = n2880 ;
assign n2883 = PE0_act_regs_3_data_n2882 ;
assign n2884 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2885 = n2880 ;
assign n2887 = PE0_act_regs_2_data_n2886 ;
assign n2888 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2889 = n2880 ;
assign n2891 = PE0_act_regs_1_data_n2890 ;
assign n2892 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2893 = n2880 ;
assign n2895 = PE0_act_regs_0_data_n2894 ;
assign n2896 =  ( n2892 ) ? ( n2895 ) : ( bv_20_0_n419 ) ;
assign n2897 =  ( n2888 ) ? ( n2891 ) : ( n2896 ) ;
assign n2898 =  ( n2884 ) ? ( n2887 ) : ( n2897 ) ;
assign n2899 =  ( n2879 ) ? ( n2883 ) : ( n2898 ) ;
fun_PEActTanh  applyFunc_n2901(
    .arg0( n2899 ),
    .result( n2900 )
);
assign n2902 = n2900 ;
assign n2903 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n2904 =  ( bv_4_8_n190 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2905 = n2904 ;
assign n2907 = PE0_act_regs_3_data_n2906 ;
assign n2908 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2909 = n2904 ;
assign n2911 = PE0_act_regs_2_data_n2910 ;
assign n2912 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2913 = n2904 ;
assign n2915 = PE0_act_regs_1_data_n2914 ;
assign n2916 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2917 = n2904 ;
assign n2919 = PE0_act_regs_0_data_n2918 ;
assign n2920 =  ( n2916 ) ? ( n2919 ) : ( bv_20_0_n419 ) ;
assign n2921 =  ( n2912 ) ? ( n2915 ) : ( n2920 ) ;
assign n2922 =  ( n2908 ) ? ( n2911 ) : ( n2921 ) ;
assign n2923 =  ( n2903 ) ? ( n2907 ) : ( n2922 ) ;
fun_PEActRelu  applyFunc_n2925(
    .arg0( n2923 ),
    .result( n2924 )
);
assign n2926 = n2924 ;
assign n2927 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n2928 =  ( bv_4_8_n190 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2929 = n2928 ;
assign n2931 = PE0_act_regs_3_data_n2930 ;
assign n2932 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2933 = n2928 ;
assign n2935 = PE0_act_regs_2_data_n2934 ;
assign n2936 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2937 = n2928 ;
assign n2939 = PE0_act_regs_1_data_n2938 ;
assign n2940 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2941 = n2928 ;
assign n2943 = PE0_act_regs_0_data_n2942 ;
assign n2944 =  ( n2940 ) ? ( n2943 ) : ( bv_20_0_n419 ) ;
assign n2945 =  ( n2936 ) ? ( n2939 ) : ( n2944 ) ;
assign n2946 =  ( n2932 ) ? ( n2935 ) : ( n2945 ) ;
assign n2947 =  ( n2927 ) ? ( n2931 ) : ( n2946 ) ;
fun_PEActOnex  applyFunc_n2949(
    .arg0( n2947 ),
    .result( n2948 )
);
assign n2950 = n2948 ;
assign n2951 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n2952 =  ( n1033 ) + ( bv_32_9_n370 )  ;
assign pe0_act_buffer_addr_n2953 = n2952 ;
assign n2955 = pe0_act_buffer_data_n2954 ;
fun_Adptfloat2Fixed  applyFunc_n2957(
    .arg0( n2955 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n2956 )
);
assign n2958 = n2956 ;
assign n2959 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n2960 =  ( bv_4_9_n196 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2961 = n2960 ;
assign n2963 = PE0_act_regs_3_data_n2962 ;
assign n2964 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2965 = n2960 ;
assign n2967 = PE0_act_regs_2_data_n2966 ;
assign n2968 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2969 = n2960 ;
assign n2971 = PE0_act_regs_1_data_n2970 ;
assign n2972 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2973 = n2960 ;
assign n2975 = PE0_act_regs_0_data_n2974 ;
assign n2976 =  ( n2972 ) ? ( n2975 ) : ( bv_20_0_n419 ) ;
assign n2977 =  ( n2968 ) ? ( n2971 ) : ( n2976 ) ;
assign n2978 =  ( n2964 ) ? ( n2967 ) : ( n2977 ) ;
assign n2979 =  ( n2959 ) ? ( n2963 ) : ( n2978 ) ;
assign n2980 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n2981 =  ( bv_4_9_n196 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n2982 = n2981 ;
assign n2984 = PE0_act_regs_3_data_n2983 ;
assign n2985 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n2986 = n2981 ;
assign n2988 = PE0_act_regs_2_data_n2987 ;
assign n2989 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n2990 = n2981 ;
assign n2992 = PE0_act_regs_1_data_n2991 ;
assign n2993 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n2994 = n2981 ;
assign n2996 = PE0_act_regs_0_data_n2995 ;
assign n2997 =  ( n2993 ) ? ( n2996 ) : ( bv_20_0_n419 ) ;
assign n2998 =  ( n2989 ) ? ( n2992 ) : ( n2997 ) ;
assign n2999 =  ( n2985 ) ? ( n2988 ) : ( n2998 ) ;
assign n3000 =  ( n2980 ) ? ( n2984 ) : ( n2999 ) ;
assign n3001 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n3002 = n2981 ;
assign n3004 = PE0_act_regs_3_data_n3003 ;
assign n3005 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3006 = n2981 ;
assign n3008 = PE0_act_regs_2_data_n3007 ;
assign n3009 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3010 = n2981 ;
assign n3012 = PE0_act_regs_1_data_n3011 ;
assign n3013 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3014 = n2981 ;
assign n3016 = PE0_act_regs_0_data_n3015 ;
assign n3017 =  ( n3013 ) ? ( n3016 ) : ( bv_20_0_n419 ) ;
assign n3018 =  ( n3009 ) ? ( n3012 ) : ( n3017 ) ;
assign n3019 =  ( n3005 ) ? ( n3008 ) : ( n3018 ) ;
assign n3020 =  ( n3001 ) ? ( n3004 ) : ( n3019 ) ;
fun_PEActEadd  applyFunc_n3022(
    .arg0( n3000 ),
    .arg1( n3020 ),
    .result( n3021 )
);
assign n3023 = n3021 ;
assign n3024 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n3025 =  ( bv_4_9_n196 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3026 = n3025 ;
assign n3028 = PE0_act_regs_3_data_n3027 ;
assign n3029 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3030 = n3025 ;
assign n3032 = PE0_act_regs_2_data_n3031 ;
assign n3033 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3034 = n3025 ;
assign n3036 = PE0_act_regs_1_data_n3035 ;
assign n3037 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3038 = n3025 ;
assign n3040 = PE0_act_regs_0_data_n3039 ;
assign n3041 =  ( n3037 ) ? ( n3040 ) : ( bv_20_0_n419 ) ;
assign n3042 =  ( n3033 ) ? ( n3036 ) : ( n3041 ) ;
assign n3043 =  ( n3029 ) ? ( n3032 ) : ( n3042 ) ;
assign n3044 =  ( n3024 ) ? ( n3028 ) : ( n3043 ) ;
assign n3045 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n3046 = n3025 ;
assign n3048 = PE0_act_regs_3_data_n3047 ;
assign n3049 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3050 = n3025 ;
assign n3052 = PE0_act_regs_2_data_n3051 ;
assign n3053 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3054 = n3025 ;
assign n3056 = PE0_act_regs_1_data_n3055 ;
assign n3057 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3058 = n3025 ;
assign n3060 = PE0_act_regs_0_data_n3059 ;
assign n3061 =  ( n3057 ) ? ( n3060 ) : ( bv_20_0_n419 ) ;
assign n3062 =  ( n3053 ) ? ( n3056 ) : ( n3061 ) ;
assign n3063 =  ( n3049 ) ? ( n3052 ) : ( n3062 ) ;
assign n3064 =  ( n3045 ) ? ( n3048 ) : ( n3063 ) ;
fun_PEActEmul  applyFunc_n3066(
    .arg0( n3044 ),
    .arg1( n3064 ),
    .result( n3065 )
);
assign n3067 = n3065 ;
assign n3068 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n3069 =  ( bv_4_9_n196 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3070 = n3069 ;
assign n3072 = PE0_act_regs_3_data_n3071 ;
assign n3073 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3074 = n3069 ;
assign n3076 = PE0_act_regs_2_data_n3075 ;
assign n3077 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3078 = n3069 ;
assign n3080 = PE0_act_regs_1_data_n3079 ;
assign n3081 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3082 = n3069 ;
assign n3084 = PE0_act_regs_0_data_n3083 ;
assign n3085 =  ( n3081 ) ? ( n3084 ) : ( bv_20_0_n419 ) ;
assign n3086 =  ( n3077 ) ? ( n3080 ) : ( n3085 ) ;
assign n3087 =  ( n3073 ) ? ( n3076 ) : ( n3086 ) ;
assign n3088 =  ( n3068 ) ? ( n3072 ) : ( n3087 ) ;
fun_PEActSigmoid  applyFunc_n3090(
    .arg0( n3088 ),
    .result( n3089 )
);
assign n3091 = n3089 ;
assign n3092 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n3093 =  ( bv_4_9_n196 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3094 = n3093 ;
assign n3096 = PE0_act_regs_3_data_n3095 ;
assign n3097 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3098 = n3093 ;
assign n3100 = PE0_act_regs_2_data_n3099 ;
assign n3101 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3102 = n3093 ;
assign n3104 = PE0_act_regs_1_data_n3103 ;
assign n3105 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3106 = n3093 ;
assign n3108 = PE0_act_regs_0_data_n3107 ;
assign n3109 =  ( n3105 ) ? ( n3108 ) : ( bv_20_0_n419 ) ;
assign n3110 =  ( n3101 ) ? ( n3104 ) : ( n3109 ) ;
assign n3111 =  ( n3097 ) ? ( n3100 ) : ( n3110 ) ;
assign n3112 =  ( n3092 ) ? ( n3096 ) : ( n3111 ) ;
fun_PEActTanh  applyFunc_n3114(
    .arg0( n3112 ),
    .result( n3113 )
);
assign n3115 = n3113 ;
assign n3116 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n3117 =  ( bv_4_9_n196 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3118 = n3117 ;
assign n3120 = PE0_act_regs_3_data_n3119 ;
assign n3121 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3122 = n3117 ;
assign n3124 = PE0_act_regs_2_data_n3123 ;
assign n3125 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3126 = n3117 ;
assign n3128 = PE0_act_regs_1_data_n3127 ;
assign n3129 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3130 = n3117 ;
assign n3132 = PE0_act_regs_0_data_n3131 ;
assign n3133 =  ( n3129 ) ? ( n3132 ) : ( bv_20_0_n419 ) ;
assign n3134 =  ( n3125 ) ? ( n3128 ) : ( n3133 ) ;
assign n3135 =  ( n3121 ) ? ( n3124 ) : ( n3134 ) ;
assign n3136 =  ( n3116 ) ? ( n3120 ) : ( n3135 ) ;
fun_PEActRelu  applyFunc_n3138(
    .arg0( n3136 ),
    .result( n3137 )
);
assign n3139 = n3137 ;
assign n3140 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n3141 =  ( bv_4_9_n196 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3142 = n3141 ;
assign n3144 = PE0_act_regs_3_data_n3143 ;
assign n3145 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3146 = n3141 ;
assign n3148 = PE0_act_regs_2_data_n3147 ;
assign n3149 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3150 = n3141 ;
assign n3152 = PE0_act_regs_1_data_n3151 ;
assign n3153 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3154 = n3141 ;
assign n3156 = PE0_act_regs_0_data_n3155 ;
assign n3157 =  ( n3153 ) ? ( n3156 ) : ( bv_20_0_n419 ) ;
assign n3158 =  ( n3149 ) ? ( n3152 ) : ( n3157 ) ;
assign n3159 =  ( n3145 ) ? ( n3148 ) : ( n3158 ) ;
assign n3160 =  ( n3140 ) ? ( n3144 ) : ( n3159 ) ;
fun_PEActOnex  applyFunc_n3162(
    .arg0( n3160 ),
    .result( n3161 )
);
assign n3163 = n3161 ;
assign n3164 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n3165 =  ( n1033 ) + ( bv_32_10_n368 )  ;
assign pe0_act_buffer_addr_n3166 = n3165 ;
assign n3168 = pe0_act_buffer_data_n3167 ;
fun_Adptfloat2Fixed  applyFunc_n3170(
    .arg0( n3168 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n3169 )
);
assign n3171 = n3169 ;
assign n3172 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n3173 =  ( bv_4_10_n202 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3174 = n3173 ;
assign n3176 = PE0_act_regs_3_data_n3175 ;
assign n3177 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3178 = n3173 ;
assign n3180 = PE0_act_regs_2_data_n3179 ;
assign n3181 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3182 = n3173 ;
assign n3184 = PE0_act_regs_1_data_n3183 ;
assign n3185 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3186 = n3173 ;
assign n3188 = PE0_act_regs_0_data_n3187 ;
assign n3189 =  ( n3185 ) ? ( n3188 ) : ( bv_20_0_n419 ) ;
assign n3190 =  ( n3181 ) ? ( n3184 ) : ( n3189 ) ;
assign n3191 =  ( n3177 ) ? ( n3180 ) : ( n3190 ) ;
assign n3192 =  ( n3172 ) ? ( n3176 ) : ( n3191 ) ;
assign n3193 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n3194 =  ( bv_4_10_n202 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3195 = n3194 ;
assign n3197 = PE0_act_regs_3_data_n3196 ;
assign n3198 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3199 = n3194 ;
assign n3201 = PE0_act_regs_2_data_n3200 ;
assign n3202 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3203 = n3194 ;
assign n3205 = PE0_act_regs_1_data_n3204 ;
assign n3206 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3207 = n3194 ;
assign n3209 = PE0_act_regs_0_data_n3208 ;
assign n3210 =  ( n3206 ) ? ( n3209 ) : ( bv_20_0_n419 ) ;
assign n3211 =  ( n3202 ) ? ( n3205 ) : ( n3210 ) ;
assign n3212 =  ( n3198 ) ? ( n3201 ) : ( n3211 ) ;
assign n3213 =  ( n3193 ) ? ( n3197 ) : ( n3212 ) ;
assign n3214 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n3215 = n3194 ;
assign n3217 = PE0_act_regs_3_data_n3216 ;
assign n3218 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3219 = n3194 ;
assign n3221 = PE0_act_regs_2_data_n3220 ;
assign n3222 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3223 = n3194 ;
assign n3225 = PE0_act_regs_1_data_n3224 ;
assign n3226 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3227 = n3194 ;
assign n3229 = PE0_act_regs_0_data_n3228 ;
assign n3230 =  ( n3226 ) ? ( n3229 ) : ( bv_20_0_n419 ) ;
assign n3231 =  ( n3222 ) ? ( n3225 ) : ( n3230 ) ;
assign n3232 =  ( n3218 ) ? ( n3221 ) : ( n3231 ) ;
assign n3233 =  ( n3214 ) ? ( n3217 ) : ( n3232 ) ;
fun_PEActEadd  applyFunc_n3235(
    .arg0( n3213 ),
    .arg1( n3233 ),
    .result( n3234 )
);
assign n3236 = n3234 ;
assign n3237 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n3238 =  ( bv_4_10_n202 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3239 = n3238 ;
assign n3241 = PE0_act_regs_3_data_n3240 ;
assign n3242 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3243 = n3238 ;
assign n3245 = PE0_act_regs_2_data_n3244 ;
assign n3246 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3247 = n3238 ;
assign n3249 = PE0_act_regs_1_data_n3248 ;
assign n3250 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3251 = n3238 ;
assign n3253 = PE0_act_regs_0_data_n3252 ;
assign n3254 =  ( n3250 ) ? ( n3253 ) : ( bv_20_0_n419 ) ;
assign n3255 =  ( n3246 ) ? ( n3249 ) : ( n3254 ) ;
assign n3256 =  ( n3242 ) ? ( n3245 ) : ( n3255 ) ;
assign n3257 =  ( n3237 ) ? ( n3241 ) : ( n3256 ) ;
assign n3258 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n3259 = n3238 ;
assign n3261 = PE0_act_regs_3_data_n3260 ;
assign n3262 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3263 = n3238 ;
assign n3265 = PE0_act_regs_2_data_n3264 ;
assign n3266 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3267 = n3238 ;
assign n3269 = PE0_act_regs_1_data_n3268 ;
assign n3270 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3271 = n3238 ;
assign n3273 = PE0_act_regs_0_data_n3272 ;
assign n3274 =  ( n3270 ) ? ( n3273 ) : ( bv_20_0_n419 ) ;
assign n3275 =  ( n3266 ) ? ( n3269 ) : ( n3274 ) ;
assign n3276 =  ( n3262 ) ? ( n3265 ) : ( n3275 ) ;
assign n3277 =  ( n3258 ) ? ( n3261 ) : ( n3276 ) ;
fun_PEActEmul  applyFunc_n3279(
    .arg0( n3257 ),
    .arg1( n3277 ),
    .result( n3278 )
);
assign n3280 = n3278 ;
assign n3281 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n3282 =  ( bv_4_10_n202 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3283 = n3282 ;
assign n3285 = PE0_act_regs_3_data_n3284 ;
assign n3286 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3287 = n3282 ;
assign n3289 = PE0_act_regs_2_data_n3288 ;
assign n3290 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3291 = n3282 ;
assign n3293 = PE0_act_regs_1_data_n3292 ;
assign n3294 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3295 = n3282 ;
assign n3297 = PE0_act_regs_0_data_n3296 ;
assign n3298 =  ( n3294 ) ? ( n3297 ) : ( bv_20_0_n419 ) ;
assign n3299 =  ( n3290 ) ? ( n3293 ) : ( n3298 ) ;
assign n3300 =  ( n3286 ) ? ( n3289 ) : ( n3299 ) ;
assign n3301 =  ( n3281 ) ? ( n3285 ) : ( n3300 ) ;
fun_PEActSigmoid  applyFunc_n3303(
    .arg0( n3301 ),
    .result( n3302 )
);
assign n3304 = n3302 ;
assign n3305 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n3306 =  ( bv_4_10_n202 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3307 = n3306 ;
assign n3309 = PE0_act_regs_3_data_n3308 ;
assign n3310 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3311 = n3306 ;
assign n3313 = PE0_act_regs_2_data_n3312 ;
assign n3314 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3315 = n3306 ;
assign n3317 = PE0_act_regs_1_data_n3316 ;
assign n3318 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3319 = n3306 ;
assign n3321 = PE0_act_regs_0_data_n3320 ;
assign n3322 =  ( n3318 ) ? ( n3321 ) : ( bv_20_0_n419 ) ;
assign n3323 =  ( n3314 ) ? ( n3317 ) : ( n3322 ) ;
assign n3324 =  ( n3310 ) ? ( n3313 ) : ( n3323 ) ;
assign n3325 =  ( n3305 ) ? ( n3309 ) : ( n3324 ) ;
fun_PEActTanh  applyFunc_n3327(
    .arg0( n3325 ),
    .result( n3326 )
);
assign n3328 = n3326 ;
assign n3329 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n3330 =  ( bv_4_10_n202 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3331 = n3330 ;
assign n3333 = PE0_act_regs_3_data_n3332 ;
assign n3334 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3335 = n3330 ;
assign n3337 = PE0_act_regs_2_data_n3336 ;
assign n3338 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3339 = n3330 ;
assign n3341 = PE0_act_regs_1_data_n3340 ;
assign n3342 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3343 = n3330 ;
assign n3345 = PE0_act_regs_0_data_n3344 ;
assign n3346 =  ( n3342 ) ? ( n3345 ) : ( bv_20_0_n419 ) ;
assign n3347 =  ( n3338 ) ? ( n3341 ) : ( n3346 ) ;
assign n3348 =  ( n3334 ) ? ( n3337 ) : ( n3347 ) ;
assign n3349 =  ( n3329 ) ? ( n3333 ) : ( n3348 ) ;
fun_PEActRelu  applyFunc_n3351(
    .arg0( n3349 ),
    .result( n3350 )
);
assign n3352 = n3350 ;
assign n3353 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n3354 =  ( bv_4_10_n202 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3355 = n3354 ;
assign n3357 = PE0_act_regs_3_data_n3356 ;
assign n3358 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3359 = n3354 ;
assign n3361 = PE0_act_regs_2_data_n3360 ;
assign n3362 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3363 = n3354 ;
assign n3365 = PE0_act_regs_1_data_n3364 ;
assign n3366 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3367 = n3354 ;
assign n3369 = PE0_act_regs_0_data_n3368 ;
assign n3370 =  ( n3366 ) ? ( n3369 ) : ( bv_20_0_n419 ) ;
assign n3371 =  ( n3362 ) ? ( n3365 ) : ( n3370 ) ;
assign n3372 =  ( n3358 ) ? ( n3361 ) : ( n3371 ) ;
assign n3373 =  ( n3353 ) ? ( n3357 ) : ( n3372 ) ;
fun_PEActOnex  applyFunc_n3375(
    .arg0( n3373 ),
    .result( n3374 )
);
assign n3376 = n3374 ;
assign n3377 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n3378 =  ( n1033 ) + ( bv_32_11_n366 )  ;
assign pe0_act_buffer_addr_n3379 = n3378 ;
assign n3381 = pe0_act_buffer_data_n3380 ;
fun_Adptfloat2Fixed  applyFunc_n3383(
    .arg0( n3381 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n3382 )
);
assign n3384 = n3382 ;
assign n3385 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n3386 =  ( bv_4_11_n208 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3387 = n3386 ;
assign n3389 = PE0_act_regs_3_data_n3388 ;
assign n3390 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3391 = n3386 ;
assign n3393 = PE0_act_regs_2_data_n3392 ;
assign n3394 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3395 = n3386 ;
assign n3397 = PE0_act_regs_1_data_n3396 ;
assign n3398 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3399 = n3386 ;
assign n3401 = PE0_act_regs_0_data_n3400 ;
assign n3402 =  ( n3398 ) ? ( n3401 ) : ( bv_20_0_n419 ) ;
assign n3403 =  ( n3394 ) ? ( n3397 ) : ( n3402 ) ;
assign n3404 =  ( n3390 ) ? ( n3393 ) : ( n3403 ) ;
assign n3405 =  ( n3385 ) ? ( n3389 ) : ( n3404 ) ;
assign n3406 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n3407 =  ( bv_4_11_n208 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3408 = n3407 ;
assign n3410 = PE0_act_regs_3_data_n3409 ;
assign n3411 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3412 = n3407 ;
assign n3414 = PE0_act_regs_2_data_n3413 ;
assign n3415 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3416 = n3407 ;
assign n3418 = PE0_act_regs_1_data_n3417 ;
assign n3419 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3420 = n3407 ;
assign n3422 = PE0_act_regs_0_data_n3421 ;
assign n3423 =  ( n3419 ) ? ( n3422 ) : ( bv_20_0_n419 ) ;
assign n3424 =  ( n3415 ) ? ( n3418 ) : ( n3423 ) ;
assign n3425 =  ( n3411 ) ? ( n3414 ) : ( n3424 ) ;
assign n3426 =  ( n3406 ) ? ( n3410 ) : ( n3425 ) ;
assign n3427 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n3428 = n3407 ;
assign n3430 = PE0_act_regs_3_data_n3429 ;
assign n3431 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3432 = n3407 ;
assign n3434 = PE0_act_regs_2_data_n3433 ;
assign n3435 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3436 = n3407 ;
assign n3438 = PE0_act_regs_1_data_n3437 ;
assign n3439 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3440 = n3407 ;
assign n3442 = PE0_act_regs_0_data_n3441 ;
assign n3443 =  ( n3439 ) ? ( n3442 ) : ( bv_20_0_n419 ) ;
assign n3444 =  ( n3435 ) ? ( n3438 ) : ( n3443 ) ;
assign n3445 =  ( n3431 ) ? ( n3434 ) : ( n3444 ) ;
assign n3446 =  ( n3427 ) ? ( n3430 ) : ( n3445 ) ;
fun_PEActEadd  applyFunc_n3448(
    .arg0( n3426 ),
    .arg1( n3446 ),
    .result( n3447 )
);
assign n3449 = n3447 ;
assign n3450 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n3451 =  ( bv_4_11_n208 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3452 = n3451 ;
assign n3454 = PE0_act_regs_3_data_n3453 ;
assign n3455 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3456 = n3451 ;
assign n3458 = PE0_act_regs_2_data_n3457 ;
assign n3459 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3460 = n3451 ;
assign n3462 = PE0_act_regs_1_data_n3461 ;
assign n3463 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3464 = n3451 ;
assign n3466 = PE0_act_regs_0_data_n3465 ;
assign n3467 =  ( n3463 ) ? ( n3466 ) : ( bv_20_0_n419 ) ;
assign n3468 =  ( n3459 ) ? ( n3462 ) : ( n3467 ) ;
assign n3469 =  ( n3455 ) ? ( n3458 ) : ( n3468 ) ;
assign n3470 =  ( n3450 ) ? ( n3454 ) : ( n3469 ) ;
assign n3471 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n3472 = n3451 ;
assign n3474 = PE0_act_regs_3_data_n3473 ;
assign n3475 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3476 = n3451 ;
assign n3478 = PE0_act_regs_2_data_n3477 ;
assign n3479 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3480 = n3451 ;
assign n3482 = PE0_act_regs_1_data_n3481 ;
assign n3483 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3484 = n3451 ;
assign n3486 = PE0_act_regs_0_data_n3485 ;
assign n3487 =  ( n3483 ) ? ( n3486 ) : ( bv_20_0_n419 ) ;
assign n3488 =  ( n3479 ) ? ( n3482 ) : ( n3487 ) ;
assign n3489 =  ( n3475 ) ? ( n3478 ) : ( n3488 ) ;
assign n3490 =  ( n3471 ) ? ( n3474 ) : ( n3489 ) ;
fun_PEActEmul  applyFunc_n3492(
    .arg0( n3470 ),
    .arg1( n3490 ),
    .result( n3491 )
);
assign n3493 = n3491 ;
assign n3494 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n3495 =  ( bv_4_11_n208 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3496 = n3495 ;
assign n3498 = PE0_act_regs_3_data_n3497 ;
assign n3499 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3500 = n3495 ;
assign n3502 = PE0_act_regs_2_data_n3501 ;
assign n3503 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3504 = n3495 ;
assign n3506 = PE0_act_regs_1_data_n3505 ;
assign n3507 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3508 = n3495 ;
assign n3510 = PE0_act_regs_0_data_n3509 ;
assign n3511 =  ( n3507 ) ? ( n3510 ) : ( bv_20_0_n419 ) ;
assign n3512 =  ( n3503 ) ? ( n3506 ) : ( n3511 ) ;
assign n3513 =  ( n3499 ) ? ( n3502 ) : ( n3512 ) ;
assign n3514 =  ( n3494 ) ? ( n3498 ) : ( n3513 ) ;
fun_PEActSigmoid  applyFunc_n3516(
    .arg0( n3514 ),
    .result( n3515 )
);
assign n3517 = n3515 ;
assign n3518 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n3519 =  ( bv_4_11_n208 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3520 = n3519 ;
assign n3522 = PE0_act_regs_3_data_n3521 ;
assign n3523 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3524 = n3519 ;
assign n3526 = PE0_act_regs_2_data_n3525 ;
assign n3527 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3528 = n3519 ;
assign n3530 = PE0_act_regs_1_data_n3529 ;
assign n3531 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3532 = n3519 ;
assign n3534 = PE0_act_regs_0_data_n3533 ;
assign n3535 =  ( n3531 ) ? ( n3534 ) : ( bv_20_0_n419 ) ;
assign n3536 =  ( n3527 ) ? ( n3530 ) : ( n3535 ) ;
assign n3537 =  ( n3523 ) ? ( n3526 ) : ( n3536 ) ;
assign n3538 =  ( n3518 ) ? ( n3522 ) : ( n3537 ) ;
fun_PEActTanh  applyFunc_n3540(
    .arg0( n3538 ),
    .result( n3539 )
);
assign n3541 = n3539 ;
assign n3542 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n3543 =  ( bv_4_11_n208 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3544 = n3543 ;
assign n3546 = PE0_act_regs_3_data_n3545 ;
assign n3547 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3548 = n3543 ;
assign n3550 = PE0_act_regs_2_data_n3549 ;
assign n3551 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3552 = n3543 ;
assign n3554 = PE0_act_regs_1_data_n3553 ;
assign n3555 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3556 = n3543 ;
assign n3558 = PE0_act_regs_0_data_n3557 ;
assign n3559 =  ( n3555 ) ? ( n3558 ) : ( bv_20_0_n419 ) ;
assign n3560 =  ( n3551 ) ? ( n3554 ) : ( n3559 ) ;
assign n3561 =  ( n3547 ) ? ( n3550 ) : ( n3560 ) ;
assign n3562 =  ( n3542 ) ? ( n3546 ) : ( n3561 ) ;
fun_PEActRelu  applyFunc_n3564(
    .arg0( n3562 ),
    .result( n3563 )
);
assign n3565 = n3563 ;
assign n3566 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n3567 =  ( bv_4_11_n208 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3568 = n3567 ;
assign n3570 = PE0_act_regs_3_data_n3569 ;
assign n3571 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3572 = n3567 ;
assign n3574 = PE0_act_regs_2_data_n3573 ;
assign n3575 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3576 = n3567 ;
assign n3578 = PE0_act_regs_1_data_n3577 ;
assign n3579 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3580 = n3567 ;
assign n3582 = PE0_act_regs_0_data_n3581 ;
assign n3583 =  ( n3579 ) ? ( n3582 ) : ( bv_20_0_n419 ) ;
assign n3584 =  ( n3575 ) ? ( n3578 ) : ( n3583 ) ;
assign n3585 =  ( n3571 ) ? ( n3574 ) : ( n3584 ) ;
assign n3586 =  ( n3566 ) ? ( n3570 ) : ( n3585 ) ;
fun_PEActOnex  applyFunc_n3588(
    .arg0( n3586 ),
    .result( n3587 )
);
assign n3589 = n3587 ;
assign n3590 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n3591 =  ( n1033 ) + ( bv_32_12_n364 )  ;
assign pe0_act_buffer_addr_n3592 = n3591 ;
assign n3594 = pe0_act_buffer_data_n3593 ;
fun_Adptfloat2Fixed  applyFunc_n3596(
    .arg0( n3594 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n3595 )
);
assign n3597 = n3595 ;
assign n3598 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n3599 =  ( bv_4_12_n214 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3600 = n3599 ;
assign n3602 = PE0_act_regs_3_data_n3601 ;
assign n3603 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3604 = n3599 ;
assign n3606 = PE0_act_regs_2_data_n3605 ;
assign n3607 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3608 = n3599 ;
assign n3610 = PE0_act_regs_1_data_n3609 ;
assign n3611 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3612 = n3599 ;
assign n3614 = PE0_act_regs_0_data_n3613 ;
assign n3615 =  ( n3611 ) ? ( n3614 ) : ( bv_20_0_n419 ) ;
assign n3616 =  ( n3607 ) ? ( n3610 ) : ( n3615 ) ;
assign n3617 =  ( n3603 ) ? ( n3606 ) : ( n3616 ) ;
assign n3618 =  ( n3598 ) ? ( n3602 ) : ( n3617 ) ;
assign n3619 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n3620 =  ( bv_4_12_n214 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3621 = n3620 ;
assign n3623 = PE0_act_regs_3_data_n3622 ;
assign n3624 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3625 = n3620 ;
assign n3627 = PE0_act_regs_2_data_n3626 ;
assign n3628 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3629 = n3620 ;
assign n3631 = PE0_act_regs_1_data_n3630 ;
assign n3632 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3633 = n3620 ;
assign n3635 = PE0_act_regs_0_data_n3634 ;
assign n3636 =  ( n3632 ) ? ( n3635 ) : ( bv_20_0_n419 ) ;
assign n3637 =  ( n3628 ) ? ( n3631 ) : ( n3636 ) ;
assign n3638 =  ( n3624 ) ? ( n3627 ) : ( n3637 ) ;
assign n3639 =  ( n3619 ) ? ( n3623 ) : ( n3638 ) ;
assign n3640 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n3641 = n3620 ;
assign n3643 = PE0_act_regs_3_data_n3642 ;
assign n3644 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3645 = n3620 ;
assign n3647 = PE0_act_regs_2_data_n3646 ;
assign n3648 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3649 = n3620 ;
assign n3651 = PE0_act_regs_1_data_n3650 ;
assign n3652 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3653 = n3620 ;
assign n3655 = PE0_act_regs_0_data_n3654 ;
assign n3656 =  ( n3652 ) ? ( n3655 ) : ( bv_20_0_n419 ) ;
assign n3657 =  ( n3648 ) ? ( n3651 ) : ( n3656 ) ;
assign n3658 =  ( n3644 ) ? ( n3647 ) : ( n3657 ) ;
assign n3659 =  ( n3640 ) ? ( n3643 ) : ( n3658 ) ;
fun_PEActEadd  applyFunc_n3661(
    .arg0( n3639 ),
    .arg1( n3659 ),
    .result( n3660 )
);
assign n3662 = n3660 ;
assign n3663 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n3664 =  ( bv_4_12_n214 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3665 = n3664 ;
assign n3667 = PE0_act_regs_3_data_n3666 ;
assign n3668 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3669 = n3664 ;
assign n3671 = PE0_act_regs_2_data_n3670 ;
assign n3672 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3673 = n3664 ;
assign n3675 = PE0_act_regs_1_data_n3674 ;
assign n3676 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3677 = n3664 ;
assign n3679 = PE0_act_regs_0_data_n3678 ;
assign n3680 =  ( n3676 ) ? ( n3679 ) : ( bv_20_0_n419 ) ;
assign n3681 =  ( n3672 ) ? ( n3675 ) : ( n3680 ) ;
assign n3682 =  ( n3668 ) ? ( n3671 ) : ( n3681 ) ;
assign n3683 =  ( n3663 ) ? ( n3667 ) : ( n3682 ) ;
assign n3684 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n3685 = n3664 ;
assign n3687 = PE0_act_regs_3_data_n3686 ;
assign n3688 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3689 = n3664 ;
assign n3691 = PE0_act_regs_2_data_n3690 ;
assign n3692 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3693 = n3664 ;
assign n3695 = PE0_act_regs_1_data_n3694 ;
assign n3696 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3697 = n3664 ;
assign n3699 = PE0_act_regs_0_data_n3698 ;
assign n3700 =  ( n3696 ) ? ( n3699 ) : ( bv_20_0_n419 ) ;
assign n3701 =  ( n3692 ) ? ( n3695 ) : ( n3700 ) ;
assign n3702 =  ( n3688 ) ? ( n3691 ) : ( n3701 ) ;
assign n3703 =  ( n3684 ) ? ( n3687 ) : ( n3702 ) ;
fun_PEActEmul  applyFunc_n3705(
    .arg0( n3683 ),
    .arg1( n3703 ),
    .result( n3704 )
);
assign n3706 = n3704 ;
assign n3707 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n3708 =  ( bv_4_12_n214 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3709 = n3708 ;
assign n3711 = PE0_act_regs_3_data_n3710 ;
assign n3712 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3713 = n3708 ;
assign n3715 = PE0_act_regs_2_data_n3714 ;
assign n3716 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3717 = n3708 ;
assign n3719 = PE0_act_regs_1_data_n3718 ;
assign n3720 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3721 = n3708 ;
assign n3723 = PE0_act_regs_0_data_n3722 ;
assign n3724 =  ( n3720 ) ? ( n3723 ) : ( bv_20_0_n419 ) ;
assign n3725 =  ( n3716 ) ? ( n3719 ) : ( n3724 ) ;
assign n3726 =  ( n3712 ) ? ( n3715 ) : ( n3725 ) ;
assign n3727 =  ( n3707 ) ? ( n3711 ) : ( n3726 ) ;
fun_PEActSigmoid  applyFunc_n3729(
    .arg0( n3727 ),
    .result( n3728 )
);
assign n3730 = n3728 ;
assign n3731 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n3732 =  ( bv_4_12_n214 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3733 = n3732 ;
assign n3735 = PE0_act_regs_3_data_n3734 ;
assign n3736 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3737 = n3732 ;
assign n3739 = PE0_act_regs_2_data_n3738 ;
assign n3740 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3741 = n3732 ;
assign n3743 = PE0_act_regs_1_data_n3742 ;
assign n3744 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3745 = n3732 ;
assign n3747 = PE0_act_regs_0_data_n3746 ;
assign n3748 =  ( n3744 ) ? ( n3747 ) : ( bv_20_0_n419 ) ;
assign n3749 =  ( n3740 ) ? ( n3743 ) : ( n3748 ) ;
assign n3750 =  ( n3736 ) ? ( n3739 ) : ( n3749 ) ;
assign n3751 =  ( n3731 ) ? ( n3735 ) : ( n3750 ) ;
fun_PEActTanh  applyFunc_n3753(
    .arg0( n3751 ),
    .result( n3752 )
);
assign n3754 = n3752 ;
assign n3755 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n3756 =  ( bv_4_12_n214 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3757 = n3756 ;
assign n3759 = PE0_act_regs_3_data_n3758 ;
assign n3760 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3761 = n3756 ;
assign n3763 = PE0_act_regs_2_data_n3762 ;
assign n3764 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3765 = n3756 ;
assign n3767 = PE0_act_regs_1_data_n3766 ;
assign n3768 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3769 = n3756 ;
assign n3771 = PE0_act_regs_0_data_n3770 ;
assign n3772 =  ( n3768 ) ? ( n3771 ) : ( bv_20_0_n419 ) ;
assign n3773 =  ( n3764 ) ? ( n3767 ) : ( n3772 ) ;
assign n3774 =  ( n3760 ) ? ( n3763 ) : ( n3773 ) ;
assign n3775 =  ( n3755 ) ? ( n3759 ) : ( n3774 ) ;
fun_PEActRelu  applyFunc_n3777(
    .arg0( n3775 ),
    .result( n3776 )
);
assign n3778 = n3776 ;
assign n3779 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n3780 =  ( bv_4_12_n214 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3781 = n3780 ;
assign n3783 = PE0_act_regs_3_data_n3782 ;
assign n3784 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3785 = n3780 ;
assign n3787 = PE0_act_regs_2_data_n3786 ;
assign n3788 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3789 = n3780 ;
assign n3791 = PE0_act_regs_1_data_n3790 ;
assign n3792 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3793 = n3780 ;
assign n3795 = PE0_act_regs_0_data_n3794 ;
assign n3796 =  ( n3792 ) ? ( n3795 ) : ( bv_20_0_n419 ) ;
assign n3797 =  ( n3788 ) ? ( n3791 ) : ( n3796 ) ;
assign n3798 =  ( n3784 ) ? ( n3787 ) : ( n3797 ) ;
assign n3799 =  ( n3779 ) ? ( n3783 ) : ( n3798 ) ;
fun_PEActOnex  applyFunc_n3801(
    .arg0( n3799 ),
    .result( n3800 )
);
assign n3802 = n3800 ;
assign n3803 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n3804 =  ( n1033 ) + ( bv_32_13_n362 )  ;
assign pe0_act_buffer_addr_n3805 = n3804 ;
assign n3807 = pe0_act_buffer_data_n3806 ;
fun_Adptfloat2Fixed  applyFunc_n3809(
    .arg0( n3807 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n3808 )
);
assign n3810 = n3808 ;
assign n3811 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n3812 =  ( bv_4_13_n220 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3813 = n3812 ;
assign n3815 = PE0_act_regs_3_data_n3814 ;
assign n3816 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3817 = n3812 ;
assign n3819 = PE0_act_regs_2_data_n3818 ;
assign n3820 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3821 = n3812 ;
assign n3823 = PE0_act_regs_1_data_n3822 ;
assign n3824 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3825 = n3812 ;
assign n3827 = PE0_act_regs_0_data_n3826 ;
assign n3828 =  ( n3824 ) ? ( n3827 ) : ( bv_20_0_n419 ) ;
assign n3829 =  ( n3820 ) ? ( n3823 ) : ( n3828 ) ;
assign n3830 =  ( n3816 ) ? ( n3819 ) : ( n3829 ) ;
assign n3831 =  ( n3811 ) ? ( n3815 ) : ( n3830 ) ;
assign n3832 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n3833 =  ( bv_4_13_n220 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3834 = n3833 ;
assign n3836 = PE0_act_regs_3_data_n3835 ;
assign n3837 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3838 = n3833 ;
assign n3840 = PE0_act_regs_2_data_n3839 ;
assign n3841 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3842 = n3833 ;
assign n3844 = PE0_act_regs_1_data_n3843 ;
assign n3845 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3846 = n3833 ;
assign n3848 = PE0_act_regs_0_data_n3847 ;
assign n3849 =  ( n3845 ) ? ( n3848 ) : ( bv_20_0_n419 ) ;
assign n3850 =  ( n3841 ) ? ( n3844 ) : ( n3849 ) ;
assign n3851 =  ( n3837 ) ? ( n3840 ) : ( n3850 ) ;
assign n3852 =  ( n3832 ) ? ( n3836 ) : ( n3851 ) ;
assign n3853 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n3854 = n3833 ;
assign n3856 = PE0_act_regs_3_data_n3855 ;
assign n3857 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3858 = n3833 ;
assign n3860 = PE0_act_regs_2_data_n3859 ;
assign n3861 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3862 = n3833 ;
assign n3864 = PE0_act_regs_1_data_n3863 ;
assign n3865 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3866 = n3833 ;
assign n3868 = PE0_act_regs_0_data_n3867 ;
assign n3869 =  ( n3865 ) ? ( n3868 ) : ( bv_20_0_n419 ) ;
assign n3870 =  ( n3861 ) ? ( n3864 ) : ( n3869 ) ;
assign n3871 =  ( n3857 ) ? ( n3860 ) : ( n3870 ) ;
assign n3872 =  ( n3853 ) ? ( n3856 ) : ( n3871 ) ;
fun_PEActEadd  applyFunc_n3874(
    .arg0( n3852 ),
    .arg1( n3872 ),
    .result( n3873 )
);
assign n3875 = n3873 ;
assign n3876 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n3877 =  ( bv_4_13_n220 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3878 = n3877 ;
assign n3880 = PE0_act_regs_3_data_n3879 ;
assign n3881 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3882 = n3877 ;
assign n3884 = PE0_act_regs_2_data_n3883 ;
assign n3885 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3886 = n3877 ;
assign n3888 = PE0_act_regs_1_data_n3887 ;
assign n3889 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3890 = n3877 ;
assign n3892 = PE0_act_regs_0_data_n3891 ;
assign n3893 =  ( n3889 ) ? ( n3892 ) : ( bv_20_0_n419 ) ;
assign n3894 =  ( n3885 ) ? ( n3888 ) : ( n3893 ) ;
assign n3895 =  ( n3881 ) ? ( n3884 ) : ( n3894 ) ;
assign n3896 =  ( n3876 ) ? ( n3880 ) : ( n3895 ) ;
assign n3897 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n3898 = n3877 ;
assign n3900 = PE0_act_regs_3_data_n3899 ;
assign n3901 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3902 = n3877 ;
assign n3904 = PE0_act_regs_2_data_n3903 ;
assign n3905 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3906 = n3877 ;
assign n3908 = PE0_act_regs_1_data_n3907 ;
assign n3909 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3910 = n3877 ;
assign n3912 = PE0_act_regs_0_data_n3911 ;
assign n3913 =  ( n3909 ) ? ( n3912 ) : ( bv_20_0_n419 ) ;
assign n3914 =  ( n3905 ) ? ( n3908 ) : ( n3913 ) ;
assign n3915 =  ( n3901 ) ? ( n3904 ) : ( n3914 ) ;
assign n3916 =  ( n3897 ) ? ( n3900 ) : ( n3915 ) ;
fun_PEActEmul  applyFunc_n3918(
    .arg0( n3896 ),
    .arg1( n3916 ),
    .result( n3917 )
);
assign n3919 = n3917 ;
assign n3920 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n3921 =  ( bv_4_13_n220 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3922 = n3921 ;
assign n3924 = PE0_act_regs_3_data_n3923 ;
assign n3925 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3926 = n3921 ;
assign n3928 = PE0_act_regs_2_data_n3927 ;
assign n3929 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3930 = n3921 ;
assign n3932 = PE0_act_regs_1_data_n3931 ;
assign n3933 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3934 = n3921 ;
assign n3936 = PE0_act_regs_0_data_n3935 ;
assign n3937 =  ( n3933 ) ? ( n3936 ) : ( bv_20_0_n419 ) ;
assign n3938 =  ( n3929 ) ? ( n3932 ) : ( n3937 ) ;
assign n3939 =  ( n3925 ) ? ( n3928 ) : ( n3938 ) ;
assign n3940 =  ( n3920 ) ? ( n3924 ) : ( n3939 ) ;
fun_PEActSigmoid  applyFunc_n3942(
    .arg0( n3940 ),
    .result( n3941 )
);
assign n3943 = n3941 ;
assign n3944 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n3945 =  ( bv_4_13_n220 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3946 = n3945 ;
assign n3948 = PE0_act_regs_3_data_n3947 ;
assign n3949 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3950 = n3945 ;
assign n3952 = PE0_act_regs_2_data_n3951 ;
assign n3953 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3954 = n3945 ;
assign n3956 = PE0_act_regs_1_data_n3955 ;
assign n3957 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3958 = n3945 ;
assign n3960 = PE0_act_regs_0_data_n3959 ;
assign n3961 =  ( n3957 ) ? ( n3960 ) : ( bv_20_0_n419 ) ;
assign n3962 =  ( n3953 ) ? ( n3956 ) : ( n3961 ) ;
assign n3963 =  ( n3949 ) ? ( n3952 ) : ( n3962 ) ;
assign n3964 =  ( n3944 ) ? ( n3948 ) : ( n3963 ) ;
fun_PEActTanh  applyFunc_n3966(
    .arg0( n3964 ),
    .result( n3965 )
);
assign n3967 = n3965 ;
assign n3968 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n3969 =  ( bv_4_13_n220 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3970 = n3969 ;
assign n3972 = PE0_act_regs_3_data_n3971 ;
assign n3973 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3974 = n3969 ;
assign n3976 = PE0_act_regs_2_data_n3975 ;
assign n3977 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n3978 = n3969 ;
assign n3980 = PE0_act_regs_1_data_n3979 ;
assign n3981 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n3982 = n3969 ;
assign n3984 = PE0_act_regs_0_data_n3983 ;
assign n3985 =  ( n3981 ) ? ( n3984 ) : ( bv_20_0_n419 ) ;
assign n3986 =  ( n3977 ) ? ( n3980 ) : ( n3985 ) ;
assign n3987 =  ( n3973 ) ? ( n3976 ) : ( n3986 ) ;
assign n3988 =  ( n3968 ) ? ( n3972 ) : ( n3987 ) ;
fun_PEActRelu  applyFunc_n3990(
    .arg0( n3988 ),
    .result( n3989 )
);
assign n3991 = n3989 ;
assign n3992 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n3993 =  ( bv_4_13_n220 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n3994 = n3993 ;
assign n3996 = PE0_act_regs_3_data_n3995 ;
assign n3997 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n3998 = n3993 ;
assign n4000 = PE0_act_regs_2_data_n3999 ;
assign n4001 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n4002 = n3993 ;
assign n4004 = PE0_act_regs_1_data_n4003 ;
assign n4005 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n4006 = n3993 ;
assign n4008 = PE0_act_regs_0_data_n4007 ;
assign n4009 =  ( n4005 ) ? ( n4008 ) : ( bv_20_0_n419 ) ;
assign n4010 =  ( n4001 ) ? ( n4004 ) : ( n4009 ) ;
assign n4011 =  ( n3997 ) ? ( n4000 ) : ( n4010 ) ;
assign n4012 =  ( n3992 ) ? ( n3996 ) : ( n4011 ) ;
fun_PEActOnex  applyFunc_n4014(
    .arg0( n4012 ),
    .result( n4013 )
);
assign n4015 = n4013 ;
assign n4016 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n4017 =  ( n1033 ) + ( bv_32_14_n360 )  ;
assign pe0_act_buffer_addr_n4018 = n4017 ;
assign n4020 = pe0_act_buffer_data_n4019 ;
fun_Adptfloat2Fixed  applyFunc_n4022(
    .arg0( n4020 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n4021 )
);
assign n4023 = n4021 ;
assign n4024 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n4025 =  ( bv_4_14_n429 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n4026 = n4025 ;
assign n4028 = PE0_act_regs_3_data_n4027 ;
assign n4029 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n4030 = n4025 ;
assign n4032 = PE0_act_regs_2_data_n4031 ;
assign n4033 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n4034 = n4025 ;
assign n4036 = PE0_act_regs_1_data_n4035 ;
assign n4037 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n4038 = n4025 ;
assign n4040 = PE0_act_regs_0_data_n4039 ;
assign n4041 =  ( n4037 ) ? ( n4040 ) : ( bv_20_0_n419 ) ;
assign n4042 =  ( n4033 ) ? ( n4036 ) : ( n4041 ) ;
assign n4043 =  ( n4029 ) ? ( n4032 ) : ( n4042 ) ;
assign n4044 =  ( n4024 ) ? ( n4028 ) : ( n4043 ) ;
assign n4045 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n4046 =  ( bv_4_14_n429 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n4047 = n4046 ;
assign n4049 = PE0_act_regs_3_data_n4048 ;
assign n4050 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n4051 = n4046 ;
assign n4053 = PE0_act_regs_2_data_n4052 ;
assign n4054 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n4055 = n4046 ;
assign n4057 = PE0_act_regs_1_data_n4056 ;
assign n4058 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n4059 = n4046 ;
assign n4061 = PE0_act_regs_0_data_n4060 ;
assign n4062 =  ( n4058 ) ? ( n4061 ) : ( bv_20_0_n419 ) ;
assign n4063 =  ( n4054 ) ? ( n4057 ) : ( n4062 ) ;
assign n4064 =  ( n4050 ) ? ( n4053 ) : ( n4063 ) ;
assign n4065 =  ( n4045 ) ? ( n4049 ) : ( n4064 ) ;
assign n4066 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n4067 = n4046 ;
assign n4069 = PE0_act_regs_3_data_n4068 ;
assign n4070 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n4071 = n4046 ;
assign n4073 = PE0_act_regs_2_data_n4072 ;
assign n4074 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n4075 = n4046 ;
assign n4077 = PE0_act_regs_1_data_n4076 ;
assign n4078 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n4079 = n4046 ;
assign n4081 = PE0_act_regs_0_data_n4080 ;
assign n4082 =  ( n4078 ) ? ( n4081 ) : ( bv_20_0_n419 ) ;
assign n4083 =  ( n4074 ) ? ( n4077 ) : ( n4082 ) ;
assign n4084 =  ( n4070 ) ? ( n4073 ) : ( n4083 ) ;
assign n4085 =  ( n4066 ) ? ( n4069 ) : ( n4084 ) ;
fun_PEActEadd  applyFunc_n4087(
    .arg0( n4065 ),
    .arg1( n4085 ),
    .result( n4086 )
);
assign n4088 = n4086 ;
assign n4089 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n4090 =  ( bv_4_14_n429 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n4091 = n4090 ;
assign n4093 = PE0_act_regs_3_data_n4092 ;
assign n4094 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n4095 = n4090 ;
assign n4097 = PE0_act_regs_2_data_n4096 ;
assign n4098 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n4099 = n4090 ;
assign n4101 = PE0_act_regs_1_data_n4100 ;
assign n4102 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n4103 = n4090 ;
assign n4105 = PE0_act_regs_0_data_n4104 ;
assign n4106 =  ( n4102 ) ? ( n4105 ) : ( bv_20_0_n419 ) ;
assign n4107 =  ( n4098 ) ? ( n4101 ) : ( n4106 ) ;
assign n4108 =  ( n4094 ) ? ( n4097 ) : ( n4107 ) ;
assign n4109 =  ( n4089 ) ? ( n4093 ) : ( n4108 ) ;
assign n4110 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n4111 = n4090 ;
assign n4113 = PE0_act_regs_3_data_n4112 ;
assign n4114 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n4115 = n4090 ;
assign n4117 = PE0_act_regs_2_data_n4116 ;
assign n4118 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n4119 = n4090 ;
assign n4121 = PE0_act_regs_1_data_n4120 ;
assign n4122 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n4123 = n4090 ;
assign n4125 = PE0_act_regs_0_data_n4124 ;
assign n4126 =  ( n4122 ) ? ( n4125 ) : ( bv_20_0_n419 ) ;
assign n4127 =  ( n4118 ) ? ( n4121 ) : ( n4126 ) ;
assign n4128 =  ( n4114 ) ? ( n4117 ) : ( n4127 ) ;
assign n4129 =  ( n4110 ) ? ( n4113 ) : ( n4128 ) ;
fun_PEActEmul  applyFunc_n4131(
    .arg0( n4109 ),
    .arg1( n4129 ),
    .result( n4130 )
);
assign n4132 = n4130 ;
assign n4133 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n4134 =  ( bv_4_14_n429 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n4135 = n4134 ;
assign n4137 = PE0_act_regs_3_data_n4136 ;
assign n4138 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n4139 = n4134 ;
assign n4141 = PE0_act_regs_2_data_n4140 ;
assign n4142 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n4143 = n4134 ;
assign n4145 = PE0_act_regs_1_data_n4144 ;
assign n4146 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n4147 = n4134 ;
assign n4149 = PE0_act_regs_0_data_n4148 ;
assign n4150 =  ( n4146 ) ? ( n4149 ) : ( bv_20_0_n419 ) ;
assign n4151 =  ( n4142 ) ? ( n4145 ) : ( n4150 ) ;
assign n4152 =  ( n4138 ) ? ( n4141 ) : ( n4151 ) ;
assign n4153 =  ( n4133 ) ? ( n4137 ) : ( n4152 ) ;
fun_PEActSigmoid  applyFunc_n4155(
    .arg0( n4153 ),
    .result( n4154 )
);
assign n4156 = n4154 ;
assign n4157 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n4158 =  ( bv_4_14_n429 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n4159 = n4158 ;
assign n4161 = PE0_act_regs_3_data_n4160 ;
assign n4162 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n4163 = n4158 ;
assign n4165 = PE0_act_regs_2_data_n4164 ;
assign n4166 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n4167 = n4158 ;
assign n4169 = PE0_act_regs_1_data_n4168 ;
assign n4170 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n4171 = n4158 ;
assign n4173 = PE0_act_regs_0_data_n4172 ;
assign n4174 =  ( n4170 ) ? ( n4173 ) : ( bv_20_0_n419 ) ;
assign n4175 =  ( n4166 ) ? ( n4169 ) : ( n4174 ) ;
assign n4176 =  ( n4162 ) ? ( n4165 ) : ( n4175 ) ;
assign n4177 =  ( n4157 ) ? ( n4161 ) : ( n4176 ) ;
fun_PEActTanh  applyFunc_n4179(
    .arg0( n4177 ),
    .result( n4178 )
);
assign n4180 = n4178 ;
assign n4181 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n4182 =  ( bv_4_14_n429 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n4183 = n4182 ;
assign n4185 = PE0_act_regs_3_data_n4184 ;
assign n4186 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n4187 = n4182 ;
assign n4189 = PE0_act_regs_2_data_n4188 ;
assign n4190 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n4191 = n4182 ;
assign n4193 = PE0_act_regs_1_data_n4192 ;
assign n4194 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n4195 = n4182 ;
assign n4197 = PE0_act_regs_0_data_n4196 ;
assign n4198 =  ( n4194 ) ? ( n4197 ) : ( bv_20_0_n419 ) ;
assign n4199 =  ( n4190 ) ? ( n4193 ) : ( n4198 ) ;
assign n4200 =  ( n4186 ) ? ( n4189 ) : ( n4199 ) ;
assign n4201 =  ( n4181 ) ? ( n4185 ) : ( n4200 ) ;
fun_PEActRelu  applyFunc_n4203(
    .arg0( n4201 ),
    .result( n4202 )
);
assign n4204 = n4202 ;
assign n4205 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n4206 =  ( bv_4_14_n429 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n4207 = n4206 ;
assign n4209 = PE0_act_regs_3_data_n4208 ;
assign n4210 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n4211 = n4206 ;
assign n4213 = PE0_act_regs_2_data_n4212 ;
assign n4214 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n4215 = n4206 ;
assign n4217 = PE0_act_regs_1_data_n4216 ;
assign n4218 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n4219 = n4206 ;
assign n4221 = PE0_act_regs_0_data_n4220 ;
assign n4222 =  ( n4218 ) ? ( n4221 ) : ( bv_20_0_n419 ) ;
assign n4223 =  ( n4214 ) ? ( n4217 ) : ( n4222 ) ;
assign n4224 =  ( n4210 ) ? ( n4213 ) : ( n4223 ) ;
assign n4225 =  ( n4205 ) ? ( n4209 ) : ( n4224 ) ;
fun_PEActOnex  applyFunc_n4227(
    .arg0( n4225 ),
    .result( n4226 )
);
assign n4228 = n4226 ;
assign n4229 =  ( bv_20_0_n419 ) + ( bv_20_0_n419 )  ;
assign n4230 =  ( n1033 ) + ( bv_32_15_n358 )  ;
assign pe0_act_buffer_addr_n4231 = n4230 ;
assign n4233 = pe0_act_buffer_data_n4232 ;
fun_Adptfloat2Fixed  applyFunc_n4235(
    .arg0( n4233 ),
    .arg1( pe0_act_mngr_adpfloat_bias ),
    .result( n4234 )
);
assign n4236 = n4234 ;
assign n4237 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n4238 =  ( bv_4_15_n401 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n4239 = n4238 ;
assign n4241 = PE0_act_regs_3_data_n4240 ;
assign n4242 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n4243 = n4238 ;
assign n4245 = PE0_act_regs_2_data_n4244 ;
assign n4246 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n4247 = n4238 ;
assign n4249 = PE0_act_regs_1_data_n4248 ;
assign n4250 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n4251 = n4238 ;
assign n4253 = PE0_act_regs_0_data_n4252 ;
assign n4254 =  ( n4250 ) ? ( n4253 ) : ( bv_20_0_n419 ) ;
assign n4255 =  ( n4246 ) ? ( n4249 ) : ( n4254 ) ;
assign n4256 =  ( n4242 ) ? ( n4245 ) : ( n4255 ) ;
assign n4257 =  ( n4237 ) ? ( n4241 ) : ( n4256 ) ;
assign n4258 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n4259 =  ( bv_4_15_n401 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n4260 = n4259 ;
assign n4262 = PE0_act_regs_3_data_n4261 ;
assign n4263 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n4264 = n4259 ;
assign n4266 = PE0_act_regs_2_data_n4265 ;
assign n4267 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n4268 = n4259 ;
assign n4270 = PE0_act_regs_1_data_n4269 ;
assign n4271 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n4272 = n4259 ;
assign n4274 = PE0_act_regs_0_data_n4273 ;
assign n4275 =  ( n4271 ) ? ( n4274 ) : ( bv_20_0_n419 ) ;
assign n4276 =  ( n4267 ) ? ( n4270 ) : ( n4275 ) ;
assign n4277 =  ( n4263 ) ? ( n4266 ) : ( n4276 ) ;
assign n4278 =  ( n4258 ) ? ( n4262 ) : ( n4277 ) ;
assign n4279 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n4280 = n4259 ;
assign n4282 = PE0_act_regs_3_data_n4281 ;
assign n4283 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n4284 = n4259 ;
assign n4286 = PE0_act_regs_2_data_n4285 ;
assign n4287 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n4288 = n4259 ;
assign n4290 = PE0_act_regs_1_data_n4289 ;
assign n4291 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n4292 = n4259 ;
assign n4294 = PE0_act_regs_0_data_n4293 ;
assign n4295 =  ( n4291 ) ? ( n4294 ) : ( bv_20_0_n419 ) ;
assign n4296 =  ( n4287 ) ? ( n4290 ) : ( n4295 ) ;
assign n4297 =  ( n4283 ) ? ( n4286 ) : ( n4296 ) ;
assign n4298 =  ( n4279 ) ? ( n4282 ) : ( n4297 ) ;
fun_PEActEadd  applyFunc_n4300(
    .arg0( n4278 ),
    .arg1( n4298 ),
    .result( n4299 )
);
assign n4301 = n4299 ;
assign n4302 =  ( n1041 ) == ( bv_2_3_n399 )  ;
assign n4303 =  ( bv_4_15_n401 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n4304 = n4303 ;
assign n4306 = PE0_act_regs_3_data_n4305 ;
assign n4307 =  ( n1041 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n4308 = n4303 ;
assign n4310 = PE0_act_regs_2_data_n4309 ;
assign n4311 =  ( n1041 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n4312 = n4303 ;
assign n4314 = PE0_act_regs_1_data_n4313 ;
assign n4315 =  ( n1041 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n4316 = n4303 ;
assign n4318 = PE0_act_regs_0_data_n4317 ;
assign n4319 =  ( n4315 ) ? ( n4318 ) : ( bv_20_0_n419 ) ;
assign n4320 =  ( n4311 ) ? ( n4314 ) : ( n4319 ) ;
assign n4321 =  ( n4307 ) ? ( n4310 ) : ( n4320 ) ;
assign n4322 =  ( n4302 ) ? ( n4306 ) : ( n4321 ) ;
assign n4323 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign PE0_act_regs_3_addr_n4324 = n4303 ;
assign n4326 = PE0_act_regs_3_data_n4325 ;
assign n4327 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n4328 = n4303 ;
assign n4330 = PE0_act_regs_2_data_n4329 ;
assign n4331 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n4332 = n4303 ;
assign n4334 = PE0_act_regs_1_data_n4333 ;
assign n4335 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n4336 = n4303 ;
assign n4338 = PE0_act_regs_0_data_n4337 ;
assign n4339 =  ( n4335 ) ? ( n4338 ) : ( bv_20_0_n419 ) ;
assign n4340 =  ( n4331 ) ? ( n4334 ) : ( n4339 ) ;
assign n4341 =  ( n4327 ) ? ( n4330 ) : ( n4340 ) ;
assign n4342 =  ( n4323 ) ? ( n4326 ) : ( n4341 ) ;
fun_PEActEmul  applyFunc_n4344(
    .arg0( n4322 ),
    .arg1( n4342 ),
    .result( n4343 )
);
assign n4345 = n4343 ;
assign n4346 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n4347 =  ( bv_4_15_n401 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n4348 = n4347 ;
assign n4350 = PE0_act_regs_3_data_n4349 ;
assign n4351 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n4352 = n4347 ;
assign n4354 = PE0_act_regs_2_data_n4353 ;
assign n4355 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n4356 = n4347 ;
assign n4358 = PE0_act_regs_1_data_n4357 ;
assign n4359 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n4360 = n4347 ;
assign n4362 = PE0_act_regs_0_data_n4361 ;
assign n4363 =  ( n4359 ) ? ( n4362 ) : ( bv_20_0_n419 ) ;
assign n4364 =  ( n4355 ) ? ( n4358 ) : ( n4363 ) ;
assign n4365 =  ( n4351 ) ? ( n4354 ) : ( n4364 ) ;
assign n4366 =  ( n4346 ) ? ( n4350 ) : ( n4365 ) ;
fun_PEActSigmoid  applyFunc_n4368(
    .arg0( n4366 ),
    .result( n4367 )
);
assign n4369 = n4367 ;
assign n4370 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n4371 =  ( bv_4_15_n401 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n4372 = n4371 ;
assign n4374 = PE0_act_regs_3_data_n4373 ;
assign n4375 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n4376 = n4371 ;
assign n4378 = PE0_act_regs_2_data_n4377 ;
assign n4379 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n4380 = n4371 ;
assign n4382 = PE0_act_regs_1_data_n4381 ;
assign n4383 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n4384 = n4371 ;
assign n4386 = PE0_act_regs_0_data_n4385 ;
assign n4387 =  ( n4383 ) ? ( n4386 ) : ( bv_20_0_n419 ) ;
assign n4388 =  ( n4379 ) ? ( n4382 ) : ( n4387 ) ;
assign n4389 =  ( n4375 ) ? ( n4378 ) : ( n4388 ) ;
assign n4390 =  ( n4370 ) ? ( n4374 ) : ( n4389 ) ;
fun_PEActTanh  applyFunc_n4392(
    .arg0( n4390 ),
    .result( n4391 )
);
assign n4393 = n4391 ;
assign n4394 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n4395 =  ( bv_4_15_n401 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n4396 = n4395 ;
assign n4398 = PE0_act_regs_3_data_n4397 ;
assign n4399 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n4400 = n4395 ;
assign n4402 = PE0_act_regs_2_data_n4401 ;
assign n4403 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n4404 = n4395 ;
assign n4406 = PE0_act_regs_1_data_n4405 ;
assign n4407 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n4408 = n4395 ;
assign n4410 = PE0_act_regs_0_data_n4409 ;
assign n4411 =  ( n4407 ) ? ( n4410 ) : ( bv_20_0_n419 ) ;
assign n4412 =  ( n4403 ) ? ( n4406 ) : ( n4411 ) ;
assign n4413 =  ( n4399 ) ? ( n4402 ) : ( n4412 ) ;
assign n4414 =  ( n4394 ) ? ( n4398 ) : ( n4413 ) ;
fun_PEActRelu  applyFunc_n4416(
    .arg0( n4414 ),
    .result( n4415 )
);
assign n4417 = n4415 ;
assign n4418 =  ( n398 ) == ( bv_2_3_n399 )  ;
assign n4419 =  ( bv_4_15_n401 ) + ( bv_4_0_n402 )  ;
assign PE0_act_regs_3_addr_n4420 = n4419 ;
assign n4422 = PE0_act_regs_3_data_n4421 ;
assign n4423 =  ( n398 ) == ( bv_2_2_n224 )  ;
assign PE0_act_regs_2_addr_n4424 = n4419 ;
assign n4426 = PE0_act_regs_2_data_n4425 ;
assign n4427 =  ( n398 ) == ( bv_2_1_n45 )  ;
assign PE0_act_regs_1_addr_n4428 = n4419 ;
assign n4430 = PE0_act_regs_1_data_n4429 ;
assign n4431 =  ( n398 ) == ( bv_2_0_n41 )  ;
assign PE0_act_regs_0_addr_n4432 = n4419 ;
assign n4434 = PE0_act_regs_0_data_n4433 ;
assign n4435 =  ( n4431 ) ? ( n4434 ) : ( bv_20_0_n419 ) ;
assign n4436 =  ( n4427 ) ? ( n4430 ) : ( n4435 ) ;
assign n4437 =  ( n4423 ) ? ( n4426 ) : ( n4436 ) ;
assign n4438 =  ( n4418 ) ? ( n4422 ) : ( n4437 ) ;
fun_PEActOnex  applyFunc_n4440(
    .arg0( n4438 ),
    .result( n4439 )
);
assign n4441 = n4439 ;
always @(posedge clk) begin
   if(rst) begin
   end
   else if(__ILA_pe_act_valid__) begin
       if ( __ILA_pe_act_decode_of_PE0_act_child_op_inpe__ && __ILA_pe_act_grant__[8] ) begin
           act_port_ready <= bv_1_0_n32;
       end
       if ( __ILA_pe_act_decode_of_PE0_act_child_op_outgb__ && __ILA_pe_act_grant__[9] ) begin
           output_port_addr <= n245;
       end
       if ( __ILA_pe_act_decode_of_PE0_act_child_op_outgb__ && __ILA_pe_act_grant__[9] ) begin
           output_port_valid <= bv_1_1_n0;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_out_sent__ && __ILA_pe_act_grant__[18] ) begin
           output_port_valid <= bv_1_0_n32;
       end
       if ( __ILA_pe_act_decode_of_PE0_act_child_op_load_zero__ && __ILA_pe_act_grant__[5] ) begin
           done <= n252;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_load__ && __ILA_pe_act_grant__[6] ) begin
           done <= n258;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_store__ && __ILA_pe_act_grant__[7] ) begin
           done <= n264;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_inpe__ && __ILA_pe_act_grant__[8] ) begin
           done <= n270;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_outgb__ && __ILA_pe_act_grant__[9] ) begin
           done <= n276;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_copy__ && __ILA_pe_act_grant__[10] ) begin
           done <= n282;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_eadd__ && __ILA_pe_act_grant__[11] ) begin
           done <= n288;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_emul__ && __ILA_pe_act_grant__[12] ) begin
           done <= n294;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_sigm__ && __ILA_pe_act_grant__[13] ) begin
           done <= n300;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_tanh__ && __ILA_pe_act_grant__[14] ) begin
           done <= n306;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_relu__ && __ILA_pe_act_grant__[15] ) begin
           done <= n312;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_onex__ && __ILA_pe_act_grant__[16] ) begin
           done <= n318;
       end
       if ( __ILA_pe_act_decode_of_PE0_act_child_op_load_zero__ && __ILA_pe_act_grant__[5] ) begin
           done_valid <= n319;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_load__ && __ILA_pe_act_grant__[6] ) begin
           done_valid <= n320;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_store__ && __ILA_pe_act_grant__[7] ) begin
           done_valid <= n321;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_inpe__ && __ILA_pe_act_grant__[8] ) begin
           done_valid <= n322;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_outgb__ && __ILA_pe_act_grant__[9] ) begin
           done_valid <= n323;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_copy__ && __ILA_pe_act_grant__[10] ) begin
           done_valid <= n324;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_eadd__ && __ILA_pe_act_grant__[11] ) begin
           done_valid <= n325;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_emul__ && __ILA_pe_act_grant__[12] ) begin
           done_valid <= n326;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_sigm__ && __ILA_pe_act_grant__[13] ) begin
           done_valid <= n327;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_tanh__ && __ILA_pe_act_grant__[14] ) begin
           done_valid <= n328;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_relu__ && __ILA_pe_act_grant__[15] ) begin
           done_valid <= n329;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_onex__ && __ILA_pe_act_grant__[16] ) begin
           done_valid <= n330;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_done_sent__ && __ILA_pe_act_grant__[19] ) begin
           done_valid <= bv_1_0_n32;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_MNGR__ && __ILA_pe_act_grant__[0] ) begin
           pe0_act_mngr_is_valid <= n331;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_MNGR__ && __ILA_pe_act_grant__[0] ) begin
           pe0_act_mngr_is_zero_first <= n332;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_load_zero__ && __ILA_pe_act_grant__[5] ) begin
           pe0_act_mngr_is_zero_first <= n333;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_load__ && __ILA_pe_act_grant__[6] ) begin
           pe0_act_mngr_is_zero_first <= n334;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_store__ && __ILA_pe_act_grant__[7] ) begin
           pe0_act_mngr_is_zero_first <= n335;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_inpe__ && __ILA_pe_act_grant__[8] ) begin
           pe0_act_mngr_is_zero_first <= n336;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_outgb__ && __ILA_pe_act_grant__[9] ) begin
           pe0_act_mngr_is_zero_first <= n337;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_copy__ && __ILA_pe_act_grant__[10] ) begin
           pe0_act_mngr_is_zero_first <= n338;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_eadd__ && __ILA_pe_act_grant__[11] ) begin
           pe0_act_mngr_is_zero_first <= n339;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_emul__ && __ILA_pe_act_grant__[12] ) begin
           pe0_act_mngr_is_zero_first <= n340;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_sigm__ && __ILA_pe_act_grant__[13] ) begin
           pe0_act_mngr_is_zero_first <= n341;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_tanh__ && __ILA_pe_act_grant__[14] ) begin
           pe0_act_mngr_is_zero_first <= n342;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_relu__ && __ILA_pe_act_grant__[15] ) begin
           pe0_act_mngr_is_zero_first <= n343;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_onex__ && __ILA_pe_act_grant__[16] ) begin
           pe0_act_mngr_is_zero_first <= n344;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_MNGR__ && __ILA_pe_act_grant__[0] ) begin
           pe0_act_mngr_adpfloat_bias <= n345;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_MNGR__ && __ILA_pe_act_grant__[0] ) begin
           pe0_act_mngr_num_inst <= n346;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_MNGR__ && __ILA_pe_act_grant__[0] ) begin
           pe0_act_mngr_num_output <= data_in_4;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_MNGR__ && __ILA_pe_act_grant__[0] ) begin
           pe0_act_mngr_buffer_addr_base <= n348;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_MNGR__ && __ILA_pe_act_grant__[0] ) begin
           pe0_act_mngr_output_addr_base <= data_in_8;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_0_15__ && __ILA_pe_act_grant__[1] ) begin
           act_vector_0_15_Inst_0 <= data_in_0;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_0_15__ && __ILA_pe_act_grant__[1] ) begin
           act_vector_0_15_Inst_1 <= data_in_1;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_0_15__ && __ILA_pe_act_grant__[1] ) begin
           act_vector_0_15_Inst_2 <= data_in_2;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_0_15__ && __ILA_pe_act_grant__[1] ) begin
           act_vector_0_15_Inst_3 <= data_in_3;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_0_15__ && __ILA_pe_act_grant__[1] ) begin
           act_vector_0_15_Inst_4 <= data_in_4;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_0_15__ && __ILA_pe_act_grant__[1] ) begin
           act_vector_0_15_Inst_5 <= data_in_5;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_0_15__ && __ILA_pe_act_grant__[1] ) begin
           act_vector_0_15_Inst_6 <= data_in_6;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_0_15__ && __ILA_pe_act_grant__[1] ) begin
           act_vector_0_15_Inst_7 <= data_in_7;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_0_15__ && __ILA_pe_act_grant__[1] ) begin
           act_vector_0_15_Inst_8 <= data_in_8;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_0_15__ && __ILA_pe_act_grant__[1] ) begin
           act_vector_0_15_Inst_9 <= data_in_9;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_0_15__ && __ILA_pe_act_grant__[1] ) begin
           act_vector_0_15_Inst_10 <= data_in_10;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_0_15__ && __ILA_pe_act_grant__[1] ) begin
           act_vector_0_15_Inst_11 <= data_in_11;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_0_15__ && __ILA_pe_act_grant__[1] ) begin
           act_vector_0_15_Inst_12 <= data_in_12;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_0_15__ && __ILA_pe_act_grant__[1] ) begin
           act_vector_0_15_Inst_13 <= data_in_13;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_0_15__ && __ILA_pe_act_grant__[1] ) begin
           act_vector_0_15_Inst_14 <= data_in_14;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_0_15__ && __ILA_pe_act_grant__[1] ) begin
           act_vector_0_15_Inst_15 <= data_in_15;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_16_31__ && __ILA_pe_act_grant__[2] ) begin
           act_vector_16_31_Inst_0 <= data_in_0;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_16_31__ && __ILA_pe_act_grant__[2] ) begin
           act_vector_16_31_Inst_1 <= data_in_1;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_16_31__ && __ILA_pe_act_grant__[2] ) begin
           act_vector_16_31_Inst_2 <= data_in_2;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_16_31__ && __ILA_pe_act_grant__[2] ) begin
           act_vector_16_31_Inst_3 <= data_in_3;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_16_31__ && __ILA_pe_act_grant__[2] ) begin
           act_vector_16_31_Inst_4 <= data_in_4;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_16_31__ && __ILA_pe_act_grant__[2] ) begin
           act_vector_16_31_Inst_5 <= data_in_5;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_16_31__ && __ILA_pe_act_grant__[2] ) begin
           act_vector_16_31_Inst_6 <= data_in_6;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_16_31__ && __ILA_pe_act_grant__[2] ) begin
           act_vector_16_31_Inst_7 <= data_in_7;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_16_31__ && __ILA_pe_act_grant__[2] ) begin
           act_vector_16_31_Inst_8 <= data_in_8;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_16_31__ && __ILA_pe_act_grant__[2] ) begin
           act_vector_16_31_Inst_9 <= data_in_9;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_16_31__ && __ILA_pe_act_grant__[2] ) begin
           act_vector_16_31_Inst_10 <= data_in_10;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_16_31__ && __ILA_pe_act_grant__[2] ) begin
           act_vector_16_31_Inst_11 <= data_in_11;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_16_31__ && __ILA_pe_act_grant__[2] ) begin
           act_vector_16_31_Inst_12 <= data_in_12;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_16_31__ && __ILA_pe_act_grant__[2] ) begin
           act_vector_16_31_Inst_13 <= data_in_13;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_16_31__ && __ILA_pe_act_grant__[2] ) begin
           act_vector_16_31_Inst_14 <= data_in_14;
       end
       if ( __ILA_pe_act_decode_of_PE0_CONFIG_ACT_VECTOR_16_31__ && __ILA_pe_act_grant__[2] ) begin
           act_vector_16_31_Inst_15 <= data_in_15;
       end
       if ( __ILA_pe_act_decode_of_PE0_act_child_initiate__ && __ILA_pe_act_grant__[4] ) begin
           pe0_act_is_start_reg <= bv_1_1_n0;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_load_zero__ && __ILA_pe_act_grant__[5] ) begin
           pe0_act_is_start_reg <= pe0_act_is_start_reg;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_load__ && __ILA_pe_act_grant__[6] ) begin
           pe0_act_is_start_reg <= pe0_act_is_start_reg;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_store__ && __ILA_pe_act_grant__[7] ) begin
           pe0_act_is_start_reg <= pe0_act_is_start_reg;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_inpe__ && __ILA_pe_act_grant__[8] ) begin
           pe0_act_is_start_reg <= pe0_act_is_start_reg;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_outgb__ && __ILA_pe_act_grant__[9] ) begin
           pe0_act_is_start_reg <= pe0_act_is_start_reg;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_copy__ && __ILA_pe_act_grant__[10] ) begin
           pe0_act_is_start_reg <= pe0_act_is_start_reg;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_eadd__ && __ILA_pe_act_grant__[11] ) begin
           pe0_act_is_start_reg <= pe0_act_is_start_reg;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_emul__ && __ILA_pe_act_grant__[12] ) begin
           pe0_act_is_start_reg <= pe0_act_is_start_reg;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_sigm__ && __ILA_pe_act_grant__[13] ) begin
           pe0_act_is_start_reg <= pe0_act_is_start_reg;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_tanh__ && __ILA_pe_act_grant__[14] ) begin
           pe0_act_is_start_reg <= pe0_act_is_start_reg;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_relu__ && __ILA_pe_act_grant__[15] ) begin
           pe0_act_is_start_reg <= pe0_act_is_start_reg;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_onex__ && __ILA_pe_act_grant__[16] ) begin
           pe0_act_is_start_reg <= pe0_act_is_start_reg;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_reg_store__ && __ILA_pe_act_grant__[17] ) begin
           pe0_act_is_start_reg <= pe0_act_is_start_reg;
       end
       if ( __ILA_pe_act_decode_of_PE0_act_child_initiate__ && __ILA_pe_act_grant__[4] ) begin
           pe0_act_instruction_counter <= bv_6_0_n110;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_load_zero__ && __ILA_pe_act_grant__[5] ) begin
           pe0_act_instruction_counter <= n806;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_load__ && __ILA_pe_act_grant__[6] ) begin
           pe0_act_instruction_counter <= n808;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_store__ && __ILA_pe_act_grant__[7] ) begin
           pe0_act_instruction_counter <= n810;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_inpe__ && __ILA_pe_act_grant__[8] ) begin
           pe0_act_instruction_counter <= n812;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_outgb__ && __ILA_pe_act_grant__[9] ) begin
           pe0_act_instruction_counter <= n814;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_copy__ && __ILA_pe_act_grant__[10] ) begin
           pe0_act_instruction_counter <= n816;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_eadd__ && __ILA_pe_act_grant__[11] ) begin
           pe0_act_instruction_counter <= n818;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_emul__ && __ILA_pe_act_grant__[12] ) begin
           pe0_act_instruction_counter <= n820;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_sigm__ && __ILA_pe_act_grant__[13] ) begin
           pe0_act_instruction_counter <= n822;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_tanh__ && __ILA_pe_act_grant__[14] ) begin
           pe0_act_instruction_counter <= n824;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_relu__ && __ILA_pe_act_grant__[15] ) begin
           pe0_act_instruction_counter <= n826;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_onex__ && __ILA_pe_act_grant__[16] ) begin
           pe0_act_instruction_counter <= n828;
       end
       if ( __ILA_pe_act_decode_of_PE0_act_child_initiate__ && __ILA_pe_act_grant__[4] ) begin
           pe0_act_output_counter <= bv_8_0_n354;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_load_zero__ && __ILA_pe_act_grant__[5] ) begin
           pe0_act_output_counter <= n833;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_load__ && __ILA_pe_act_grant__[6] ) begin
           pe0_act_output_counter <= n838;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_store__ && __ILA_pe_act_grant__[7] ) begin
           pe0_act_output_counter <= n843;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_inpe__ && __ILA_pe_act_grant__[8] ) begin
           pe0_act_output_counter <= n848;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_outgb__ && __ILA_pe_act_grant__[9] ) begin
           pe0_act_output_counter <= n853;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_copy__ && __ILA_pe_act_grant__[10] ) begin
           pe0_act_output_counter <= n858;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_eadd__ && __ILA_pe_act_grant__[11] ) begin
           pe0_act_output_counter <= n863;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_emul__ && __ILA_pe_act_grant__[12] ) begin
           pe0_act_output_counter <= n868;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_sigm__ && __ILA_pe_act_grant__[13] ) begin
           pe0_act_output_counter <= n873;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_tanh__ && __ILA_pe_act_grant__[14] ) begin
           pe0_act_output_counter <= n878;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_relu__ && __ILA_pe_act_grant__[15] ) begin
           pe0_act_output_counter <= n883;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_onex__ && __ILA_pe_act_grant__[16] ) begin
           pe0_act_output_counter <= n888;
       end
       if ( __ILA_pe_act_decode_of_PE0_act_child_initiate__ && __ILA_pe_act_grant__[4] ) begin
           pe0_act_state <= bv_2_1_n45;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_load_zero__ && __ILA_pe_act_grant__[5] ) begin
           pe0_act_state <= bv_2_2_n224;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_load__ && __ILA_pe_act_grant__[6] ) begin
           pe0_act_state <= bv_2_2_n224;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_store__ && __ILA_pe_act_grant__[7] ) begin
           pe0_act_state <= bv_2_2_n224;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_inpe__ && __ILA_pe_act_grant__[8] ) begin
           pe0_act_state <= bv_2_2_n224;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_outgb__ && __ILA_pe_act_grant__[9] ) begin
           pe0_act_state <= bv_2_2_n224;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_copy__ && __ILA_pe_act_grant__[10] ) begin
           pe0_act_state <= bv_2_2_n224;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_eadd__ && __ILA_pe_act_grant__[11] ) begin
           pe0_act_state <= bv_2_2_n224;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_emul__ && __ILA_pe_act_grant__[12] ) begin
           pe0_act_state <= bv_2_2_n224;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_sigm__ && __ILA_pe_act_grant__[13] ) begin
           pe0_act_state <= bv_2_2_n224;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_tanh__ && __ILA_pe_act_grant__[14] ) begin
           pe0_act_state <= bv_2_2_n224;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_relu__ && __ILA_pe_act_grant__[15] ) begin
           pe0_act_state <= bv_2_2_n224;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_onex__ && __ILA_pe_act_grant__[16] ) begin
           pe0_act_state <= bv_2_2_n224;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_reg_store__ && __ILA_pe_act_grant__[17] ) begin
           pe0_act_state <= bv_2_1_n45;
       end
       if ( __ILA_pe_act_decode_of_PE0_act_child_op_load_zero__ && __ILA_pe_act_grant__[5] ) begin
           PE0_act_reg_temp_0 <= n1029;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_load__ && __ILA_pe_act_grant__[6] ) begin
           PE0_act_reg_temp_0 <= n1040;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_inpe__ && __ILA_pe_act_grant__[8] ) begin
           PE0_act_reg_temp_0 <= PE0_core_act_vector_0;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_copy__ && __ILA_pe_act_grant__[10] ) begin
           PE0_act_reg_temp_0 <= n1062;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_eadd__ && __ILA_pe_act_grant__[11] ) begin
           PE0_act_reg_temp_0 <= n1106;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_emul__ && __ILA_pe_act_grant__[12] ) begin
           PE0_act_reg_temp_0 <= n1150;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_sigm__ && __ILA_pe_act_grant__[13] ) begin
           PE0_act_reg_temp_0 <= n1174;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_tanh__ && __ILA_pe_act_grant__[14] ) begin
           PE0_act_reg_temp_0 <= n1198;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_relu__ && __ILA_pe_act_grant__[15] ) begin
           PE0_act_reg_temp_0 <= n1222;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_onex__ && __ILA_pe_act_grant__[16] ) begin
           PE0_act_reg_temp_0 <= n1246;
       end
       if ( __ILA_pe_act_decode_of_PE0_act_child_op_load_zero__ && __ILA_pe_act_grant__[5] ) begin
           PE0_act_reg_temp_1 <= n1247;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_load__ && __ILA_pe_act_grant__[6] ) begin
           PE0_act_reg_temp_1 <= n1254;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_inpe__ && __ILA_pe_act_grant__[8] ) begin
           PE0_act_reg_temp_1 <= PE0_core_act_vector_1;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_copy__ && __ILA_pe_act_grant__[10] ) begin
           PE0_act_reg_temp_1 <= n1275;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_eadd__ && __ILA_pe_act_grant__[11] ) begin
           PE0_act_reg_temp_1 <= n1319;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_emul__ && __ILA_pe_act_grant__[12] ) begin
           PE0_act_reg_temp_1 <= n1363;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_sigm__ && __ILA_pe_act_grant__[13] ) begin
           PE0_act_reg_temp_1 <= n1387;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_tanh__ && __ILA_pe_act_grant__[14] ) begin
           PE0_act_reg_temp_1 <= n1411;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_relu__ && __ILA_pe_act_grant__[15] ) begin
           PE0_act_reg_temp_1 <= n1435;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_onex__ && __ILA_pe_act_grant__[16] ) begin
           PE0_act_reg_temp_1 <= n1459;
       end
       if ( __ILA_pe_act_decode_of_PE0_act_child_op_load_zero__ && __ILA_pe_act_grant__[5] ) begin
           PE0_act_reg_temp_2 <= n1460;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_load__ && __ILA_pe_act_grant__[6] ) begin
           PE0_act_reg_temp_2 <= n1467;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_inpe__ && __ILA_pe_act_grant__[8] ) begin
           PE0_act_reg_temp_2 <= PE0_core_act_vector_2;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_copy__ && __ILA_pe_act_grant__[10] ) begin
           PE0_act_reg_temp_2 <= n1488;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_eadd__ && __ILA_pe_act_grant__[11] ) begin
           PE0_act_reg_temp_2 <= n1532;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_emul__ && __ILA_pe_act_grant__[12] ) begin
           PE0_act_reg_temp_2 <= n1576;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_sigm__ && __ILA_pe_act_grant__[13] ) begin
           PE0_act_reg_temp_2 <= n1600;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_tanh__ && __ILA_pe_act_grant__[14] ) begin
           PE0_act_reg_temp_2 <= n1624;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_relu__ && __ILA_pe_act_grant__[15] ) begin
           PE0_act_reg_temp_2 <= n1648;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_onex__ && __ILA_pe_act_grant__[16] ) begin
           PE0_act_reg_temp_2 <= n1672;
       end
       if ( __ILA_pe_act_decode_of_PE0_act_child_op_load_zero__ && __ILA_pe_act_grant__[5] ) begin
           PE0_act_reg_temp_3 <= n1673;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_load__ && __ILA_pe_act_grant__[6] ) begin
           PE0_act_reg_temp_3 <= n1680;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_inpe__ && __ILA_pe_act_grant__[8] ) begin
           PE0_act_reg_temp_3 <= PE0_core_act_vector_3;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_copy__ && __ILA_pe_act_grant__[10] ) begin
           PE0_act_reg_temp_3 <= n1701;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_eadd__ && __ILA_pe_act_grant__[11] ) begin
           PE0_act_reg_temp_3 <= n1745;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_emul__ && __ILA_pe_act_grant__[12] ) begin
           PE0_act_reg_temp_3 <= n1789;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_sigm__ && __ILA_pe_act_grant__[13] ) begin
           PE0_act_reg_temp_3 <= n1813;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_tanh__ && __ILA_pe_act_grant__[14] ) begin
           PE0_act_reg_temp_3 <= n1837;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_relu__ && __ILA_pe_act_grant__[15] ) begin
           PE0_act_reg_temp_3 <= n1861;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_onex__ && __ILA_pe_act_grant__[16] ) begin
           PE0_act_reg_temp_3 <= n1885;
       end
       if ( __ILA_pe_act_decode_of_PE0_act_child_op_load_zero__ && __ILA_pe_act_grant__[5] ) begin
           PE0_act_reg_temp_4 <= n1886;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_load__ && __ILA_pe_act_grant__[6] ) begin
           PE0_act_reg_temp_4 <= n1893;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_inpe__ && __ILA_pe_act_grant__[8] ) begin
           PE0_act_reg_temp_4 <= PE0_core_act_vector_4;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_copy__ && __ILA_pe_act_grant__[10] ) begin
           PE0_act_reg_temp_4 <= n1914;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_eadd__ && __ILA_pe_act_grant__[11] ) begin
           PE0_act_reg_temp_4 <= n1958;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_emul__ && __ILA_pe_act_grant__[12] ) begin
           PE0_act_reg_temp_4 <= n2002;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_sigm__ && __ILA_pe_act_grant__[13] ) begin
           PE0_act_reg_temp_4 <= n2026;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_tanh__ && __ILA_pe_act_grant__[14] ) begin
           PE0_act_reg_temp_4 <= n2050;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_relu__ && __ILA_pe_act_grant__[15] ) begin
           PE0_act_reg_temp_4 <= n2074;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_onex__ && __ILA_pe_act_grant__[16] ) begin
           PE0_act_reg_temp_4 <= n2098;
       end
       if ( __ILA_pe_act_decode_of_PE0_act_child_op_load_zero__ && __ILA_pe_act_grant__[5] ) begin
           PE0_act_reg_temp_5 <= n2099;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_load__ && __ILA_pe_act_grant__[6] ) begin
           PE0_act_reg_temp_5 <= n2106;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_inpe__ && __ILA_pe_act_grant__[8] ) begin
           PE0_act_reg_temp_5 <= PE0_core_act_vector_5;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_copy__ && __ILA_pe_act_grant__[10] ) begin
           PE0_act_reg_temp_5 <= n2127;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_eadd__ && __ILA_pe_act_grant__[11] ) begin
           PE0_act_reg_temp_5 <= n2171;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_emul__ && __ILA_pe_act_grant__[12] ) begin
           PE0_act_reg_temp_5 <= n2215;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_sigm__ && __ILA_pe_act_grant__[13] ) begin
           PE0_act_reg_temp_5 <= n2239;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_tanh__ && __ILA_pe_act_grant__[14] ) begin
           PE0_act_reg_temp_5 <= n2263;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_relu__ && __ILA_pe_act_grant__[15] ) begin
           PE0_act_reg_temp_5 <= n2287;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_onex__ && __ILA_pe_act_grant__[16] ) begin
           PE0_act_reg_temp_5 <= n2311;
       end
       if ( __ILA_pe_act_decode_of_PE0_act_child_op_load_zero__ && __ILA_pe_act_grant__[5] ) begin
           PE0_act_reg_temp_6 <= n2312;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_load__ && __ILA_pe_act_grant__[6] ) begin
           PE0_act_reg_temp_6 <= n2319;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_inpe__ && __ILA_pe_act_grant__[8] ) begin
           PE0_act_reg_temp_6 <= PE0_core_act_vector_6;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_copy__ && __ILA_pe_act_grant__[10] ) begin
           PE0_act_reg_temp_6 <= n2340;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_eadd__ && __ILA_pe_act_grant__[11] ) begin
           PE0_act_reg_temp_6 <= n2384;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_emul__ && __ILA_pe_act_grant__[12] ) begin
           PE0_act_reg_temp_6 <= n2428;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_sigm__ && __ILA_pe_act_grant__[13] ) begin
           PE0_act_reg_temp_6 <= n2452;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_tanh__ && __ILA_pe_act_grant__[14] ) begin
           PE0_act_reg_temp_6 <= n2476;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_relu__ && __ILA_pe_act_grant__[15] ) begin
           PE0_act_reg_temp_6 <= n2500;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_onex__ && __ILA_pe_act_grant__[16] ) begin
           PE0_act_reg_temp_6 <= n2524;
       end
       if ( __ILA_pe_act_decode_of_PE0_act_child_op_load_zero__ && __ILA_pe_act_grant__[5] ) begin
           PE0_act_reg_temp_7 <= n2525;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_load__ && __ILA_pe_act_grant__[6] ) begin
           PE0_act_reg_temp_7 <= n2532;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_inpe__ && __ILA_pe_act_grant__[8] ) begin
           PE0_act_reg_temp_7 <= PE0_core_act_vector_7;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_copy__ && __ILA_pe_act_grant__[10] ) begin
           PE0_act_reg_temp_7 <= n2553;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_eadd__ && __ILA_pe_act_grant__[11] ) begin
           PE0_act_reg_temp_7 <= n2597;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_emul__ && __ILA_pe_act_grant__[12] ) begin
           PE0_act_reg_temp_7 <= n2641;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_sigm__ && __ILA_pe_act_grant__[13] ) begin
           PE0_act_reg_temp_7 <= n2665;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_tanh__ && __ILA_pe_act_grant__[14] ) begin
           PE0_act_reg_temp_7 <= n2689;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_relu__ && __ILA_pe_act_grant__[15] ) begin
           PE0_act_reg_temp_7 <= n2713;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_onex__ && __ILA_pe_act_grant__[16] ) begin
           PE0_act_reg_temp_7 <= n2737;
       end
       if ( __ILA_pe_act_decode_of_PE0_act_child_op_load_zero__ && __ILA_pe_act_grant__[5] ) begin
           PE0_act_reg_temp_8 <= n2738;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_load__ && __ILA_pe_act_grant__[6] ) begin
           PE0_act_reg_temp_8 <= n2745;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_inpe__ && __ILA_pe_act_grant__[8] ) begin
           PE0_act_reg_temp_8 <= PE0_core_act_vector_8;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_copy__ && __ILA_pe_act_grant__[10] ) begin
           PE0_act_reg_temp_8 <= n2766;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_eadd__ && __ILA_pe_act_grant__[11] ) begin
           PE0_act_reg_temp_8 <= n2810;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_emul__ && __ILA_pe_act_grant__[12] ) begin
           PE0_act_reg_temp_8 <= n2854;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_sigm__ && __ILA_pe_act_grant__[13] ) begin
           PE0_act_reg_temp_8 <= n2878;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_tanh__ && __ILA_pe_act_grant__[14] ) begin
           PE0_act_reg_temp_8 <= n2902;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_relu__ && __ILA_pe_act_grant__[15] ) begin
           PE0_act_reg_temp_8 <= n2926;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_onex__ && __ILA_pe_act_grant__[16] ) begin
           PE0_act_reg_temp_8 <= n2950;
       end
       if ( __ILA_pe_act_decode_of_PE0_act_child_op_load_zero__ && __ILA_pe_act_grant__[5] ) begin
           PE0_act_reg_temp_9 <= n2951;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_load__ && __ILA_pe_act_grant__[6] ) begin
           PE0_act_reg_temp_9 <= n2958;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_inpe__ && __ILA_pe_act_grant__[8] ) begin
           PE0_act_reg_temp_9 <= PE0_core_act_vector_9;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_copy__ && __ILA_pe_act_grant__[10] ) begin
           PE0_act_reg_temp_9 <= n2979;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_eadd__ && __ILA_pe_act_grant__[11] ) begin
           PE0_act_reg_temp_9 <= n3023;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_emul__ && __ILA_pe_act_grant__[12] ) begin
           PE0_act_reg_temp_9 <= n3067;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_sigm__ && __ILA_pe_act_grant__[13] ) begin
           PE0_act_reg_temp_9 <= n3091;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_tanh__ && __ILA_pe_act_grant__[14] ) begin
           PE0_act_reg_temp_9 <= n3115;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_relu__ && __ILA_pe_act_grant__[15] ) begin
           PE0_act_reg_temp_9 <= n3139;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_onex__ && __ILA_pe_act_grant__[16] ) begin
           PE0_act_reg_temp_9 <= n3163;
       end
       if ( __ILA_pe_act_decode_of_PE0_act_child_op_load_zero__ && __ILA_pe_act_grant__[5] ) begin
           PE0_act_reg_temp_10 <= n3164;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_load__ && __ILA_pe_act_grant__[6] ) begin
           PE0_act_reg_temp_10 <= n3171;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_inpe__ && __ILA_pe_act_grant__[8] ) begin
           PE0_act_reg_temp_10 <= PE0_core_act_vector_10;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_copy__ && __ILA_pe_act_grant__[10] ) begin
           PE0_act_reg_temp_10 <= n3192;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_eadd__ && __ILA_pe_act_grant__[11] ) begin
           PE0_act_reg_temp_10 <= n3236;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_emul__ && __ILA_pe_act_grant__[12] ) begin
           PE0_act_reg_temp_10 <= n3280;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_sigm__ && __ILA_pe_act_grant__[13] ) begin
           PE0_act_reg_temp_10 <= n3304;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_tanh__ && __ILA_pe_act_grant__[14] ) begin
           PE0_act_reg_temp_10 <= n3328;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_relu__ && __ILA_pe_act_grant__[15] ) begin
           PE0_act_reg_temp_10 <= n3352;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_onex__ && __ILA_pe_act_grant__[16] ) begin
           PE0_act_reg_temp_10 <= n3376;
       end
       if ( __ILA_pe_act_decode_of_PE0_act_child_op_load_zero__ && __ILA_pe_act_grant__[5] ) begin
           PE0_act_reg_temp_11 <= n3377;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_load__ && __ILA_pe_act_grant__[6] ) begin
           PE0_act_reg_temp_11 <= n3384;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_inpe__ && __ILA_pe_act_grant__[8] ) begin
           PE0_act_reg_temp_11 <= PE0_core_act_vector_11;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_copy__ && __ILA_pe_act_grant__[10] ) begin
           PE0_act_reg_temp_11 <= n3405;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_eadd__ && __ILA_pe_act_grant__[11] ) begin
           PE0_act_reg_temp_11 <= n3449;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_emul__ && __ILA_pe_act_grant__[12] ) begin
           PE0_act_reg_temp_11 <= n3493;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_sigm__ && __ILA_pe_act_grant__[13] ) begin
           PE0_act_reg_temp_11 <= n3517;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_tanh__ && __ILA_pe_act_grant__[14] ) begin
           PE0_act_reg_temp_11 <= n3541;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_relu__ && __ILA_pe_act_grant__[15] ) begin
           PE0_act_reg_temp_11 <= n3565;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_onex__ && __ILA_pe_act_grant__[16] ) begin
           PE0_act_reg_temp_11 <= n3589;
       end
       if ( __ILA_pe_act_decode_of_PE0_act_child_op_load_zero__ && __ILA_pe_act_grant__[5] ) begin
           PE0_act_reg_temp_12 <= n3590;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_load__ && __ILA_pe_act_grant__[6] ) begin
           PE0_act_reg_temp_12 <= n3597;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_inpe__ && __ILA_pe_act_grant__[8] ) begin
           PE0_act_reg_temp_12 <= PE0_core_act_vector_12;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_copy__ && __ILA_pe_act_grant__[10] ) begin
           PE0_act_reg_temp_12 <= n3618;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_eadd__ && __ILA_pe_act_grant__[11] ) begin
           PE0_act_reg_temp_12 <= n3662;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_emul__ && __ILA_pe_act_grant__[12] ) begin
           PE0_act_reg_temp_12 <= n3706;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_sigm__ && __ILA_pe_act_grant__[13] ) begin
           PE0_act_reg_temp_12 <= n3730;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_tanh__ && __ILA_pe_act_grant__[14] ) begin
           PE0_act_reg_temp_12 <= n3754;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_relu__ && __ILA_pe_act_grant__[15] ) begin
           PE0_act_reg_temp_12 <= n3778;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_onex__ && __ILA_pe_act_grant__[16] ) begin
           PE0_act_reg_temp_12 <= n3802;
       end
       if ( __ILA_pe_act_decode_of_PE0_act_child_op_load_zero__ && __ILA_pe_act_grant__[5] ) begin
           PE0_act_reg_temp_13 <= n3803;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_load__ && __ILA_pe_act_grant__[6] ) begin
           PE0_act_reg_temp_13 <= n3810;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_inpe__ && __ILA_pe_act_grant__[8] ) begin
           PE0_act_reg_temp_13 <= PE0_core_act_vector_13;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_copy__ && __ILA_pe_act_grant__[10] ) begin
           PE0_act_reg_temp_13 <= n3831;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_eadd__ && __ILA_pe_act_grant__[11] ) begin
           PE0_act_reg_temp_13 <= n3875;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_emul__ && __ILA_pe_act_grant__[12] ) begin
           PE0_act_reg_temp_13 <= n3919;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_sigm__ && __ILA_pe_act_grant__[13] ) begin
           PE0_act_reg_temp_13 <= n3943;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_tanh__ && __ILA_pe_act_grant__[14] ) begin
           PE0_act_reg_temp_13 <= n3967;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_relu__ && __ILA_pe_act_grant__[15] ) begin
           PE0_act_reg_temp_13 <= n3991;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_onex__ && __ILA_pe_act_grant__[16] ) begin
           PE0_act_reg_temp_13 <= n4015;
       end
       if ( __ILA_pe_act_decode_of_PE0_act_child_op_load_zero__ && __ILA_pe_act_grant__[5] ) begin
           PE0_act_reg_temp_14 <= n4016;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_load__ && __ILA_pe_act_grant__[6] ) begin
           PE0_act_reg_temp_14 <= n4023;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_inpe__ && __ILA_pe_act_grant__[8] ) begin
           PE0_act_reg_temp_14 <= PE0_core_act_vector_14;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_copy__ && __ILA_pe_act_grant__[10] ) begin
           PE0_act_reg_temp_14 <= n4044;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_eadd__ && __ILA_pe_act_grant__[11] ) begin
           PE0_act_reg_temp_14 <= n4088;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_emul__ && __ILA_pe_act_grant__[12] ) begin
           PE0_act_reg_temp_14 <= n4132;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_sigm__ && __ILA_pe_act_grant__[13] ) begin
           PE0_act_reg_temp_14 <= n4156;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_tanh__ && __ILA_pe_act_grant__[14] ) begin
           PE0_act_reg_temp_14 <= n4180;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_relu__ && __ILA_pe_act_grant__[15] ) begin
           PE0_act_reg_temp_14 <= n4204;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_onex__ && __ILA_pe_act_grant__[16] ) begin
           PE0_act_reg_temp_14 <= n4228;
       end
       if ( __ILA_pe_act_decode_of_PE0_act_child_op_load_zero__ && __ILA_pe_act_grant__[5] ) begin
           PE0_act_reg_temp_15 <= n4229;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_load__ && __ILA_pe_act_grant__[6] ) begin
           PE0_act_reg_temp_15 <= n4236;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_inpe__ && __ILA_pe_act_grant__[8] ) begin
           PE0_act_reg_temp_15 <= PE0_core_act_vector_15;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_copy__ && __ILA_pe_act_grant__[10] ) begin
           PE0_act_reg_temp_15 <= n4257;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_eadd__ && __ILA_pe_act_grant__[11] ) begin
           PE0_act_reg_temp_15 <= n4301;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_emul__ && __ILA_pe_act_grant__[12] ) begin
           PE0_act_reg_temp_15 <= n4345;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_sigm__ && __ILA_pe_act_grant__[13] ) begin
           PE0_act_reg_temp_15 <= n4369;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_tanh__ && __ILA_pe_act_grant__[14] ) begin
           PE0_act_reg_temp_15 <= n4393;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_relu__ && __ILA_pe_act_grant__[15] ) begin
           PE0_act_reg_temp_15 <= n4417;
       end else if ( __ILA_pe_act_decode_of_PE0_act_child_op_onex__ && __ILA_pe_act_grant__[16] ) begin
           PE0_act_reg_temp_15 <= n4441;
       end
   end
end
endmodule
