
//------> ./ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   huaixil@sat8
//  Generated date: Fri Apr  8 23:11:24 2022
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
    (
  this_val, this_rdy, this_msg, data_data_rsc_z, data_addr_rsc_z, data_wstrb_rsc_z,
      data_rw_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  reg this_rdy;
  input [168:0] this_msg;
  output [127:0] data_data_rsc_z;
  output [23:0] data_addr_rsc_z;
  output [15:0] data_wstrb_rsc_z;
  output data_rw_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  wire [127:0] nl_data_data_rsci_d;
  assign nl_data_data_rsci_d = this_msg[127:0];
  wire [23:0] nl_data_addr_rsci_d;
  assign nl_data_addr_rsci_d = this_msg[151:128];
  wire [15:0] nl_data_wstrb_rsci_d;
  assign nl_data_wstrb_rsci_d = this_msg[167:152];
  wire [0:0] nl_data_rw_rsci_d;
  assign nl_data_rw_rsci_d = this_msg[168];
  ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd1),
  .width(32'sd128)) data_data_rsci (
      .d(nl_data_data_rsci_d[127:0]),
      .z(data_data_rsc_z)
    );
  ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd2),
  .width(32'sd24)) data_addr_rsci (
      .d(nl_data_addr_rsci_d[23:0]),
      .z(data_addr_rsc_z)
    );
  ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd3),
  .width(32'sd16)) data_wstrb_rsci (
      .d(nl_data_wstrb_rsci_d[15:0]),
      .z(data_wstrb_rsc_z)
    );
  ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd4),
  .width(32'sd1)) data_rw_rsci (
      .d(nl_data_rw_rsci_d[0:0]),
      .z(data_rw_rsc_z)
    );
  ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd6),
  .width(32'sd1)) return_rsci (
      .d(this_val),
      .z(return_rsc_z)
    );
  ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd114),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk ) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk ) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module ActUnit_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
    (
  this_val, this_rdy, this_msg, data_data_rsc_z, data_addr_rsc_z, data_wstrb_rsc_z,
      data_rw_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  input [168:0] this_msg;
  output [127:0] data_data_rsc_z;
  output [23:0] data_addr_rsc_z;
  output [15:0] data_wstrb_rsc_z;
  output data_rw_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .data_data_rsc_z(data_data_rsc_z),
      .data_addr_rsc_z(data_addr_rsc_z),
      .data_wstrb_rsc_z(data_wstrb_rsc_z),
      .data_rw_rsc_z(data_rw_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   huaixil@sat8
//  Generated date: Fri Apr  8 23:11:12 2022
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_ActVectorType_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_ActVectorType_Connections_SYN_PORT_PopNB_core
    (
  this_val, this_rdy, this_msg, data_data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  reg this_rdy;
  input [319:0] this_msg;
  output [319:0] data_data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  wire [319:0] nl_data_data_rsci_d;
  assign nl_data_data_rsci_d = this_msg;
  ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd12),
  .width(32'sd320)) data_data_rsci (
      .d(nl_data_data_rsci_d[319:0]),
      .z(data_data_rsc_z)
    );
  ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd14),
  .width(32'sd1)) return_rsci (
      .d(this_val),
      .z(return_rsc_z)
    );
  ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd113),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk ) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk ) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_spec_ActVectorType_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module ActUnit_Connections_InBlocking_spec_ActVectorType_Connections_SYN_PORT_PopNB (
  this_val, this_rdy, this_msg, data_data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  input [319:0] this_msg;
  output [319:0] data_data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_ActVectorType_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_spec_ActVectorType_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .data_data_rsc_z(data_data_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   huaixil@sat8
//  Generated date: Fri Apr  8 23:10:47 2022
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
    (
  this_val, this_rdy, this_msg, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_val;
  reg this_val;
  input this_rdy;
  output [127:0] this_msg;
  reg [127:0] this_msg;
  input [127:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [127:0] m_data_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_3_cse;
  wire this_val_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire [0:0] nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd48),
  .width(32'sd128)) m_data_rsci (
      .dat(m_data_rsc_dat),
      .idat(m_data_rsci_idat)
    );
  ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd112),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1
      #(.rscid(32'sd117)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld[0:0])
    );
  assign or_3_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_val_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk ) begin
    if ( ~ ccs_MIO_arst ) begin
      this_val <= 1'b0;
    end
    else if ( or_3_cse | this_val_mx0c1 ) begin
      this_val <= ~ this_val_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk ) begin
    if ( ~ ccs_MIO_arst ) begin
      this_msg <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      this_msg <= m_data_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk ) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_3_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module ActUnit_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
    (
  this_val, this_rdy, this_msg, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_val;
  input this_rdy;
  output [127:0] this_msg;
  input [127:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .m_data_rsc_dat(m_data_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   huaixil@sat8
//  Generated date: Fri Apr  8 23:10:45 2022
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
    (
  this_val, this_rdy, this_msg, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  reg this_rdy;
  input this_msg;
  output data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  wire [0:0] nl_data_rsci_d;
  assign nl_data_rsci_d = this_msg;
  ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd49),
  .width(32'sd1)) data_rsci (
      .d(nl_data_rsci_d[0:0]),
      .z(data_rsc_z)
    );
  ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd51),
  .width(32'sd1)) return_rsci (
      .d(this_val),
      .z(return_rsc_z)
    );
  ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd111),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk ) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk ) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_bool_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module ActUnit_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB (
  this_val, this_rdy, this_msg, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  input this_msg;
  output data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core_inst (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .data_rsc_z(data_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   huaixil@sat8
//  Generated date: Fri Apr  8 23:10:42 2022
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_StreamType_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_StreamType_Connections_SYN_PORT_Push_core
    (
  this_val, this_rdy, this_msg, m_data_data_rsc_dat, m_logical_addr_rsc_dat, ccs_ccore_start_rsc_dat,
      ccs_ccore_done_sync_vld, ccs_MIO_clk, ccs_MIO_arst
);
  output this_val;
  reg this_val;
  input this_rdy;
  output [137:0] this_msg;
  input [127:0] m_data_data_rsc_dat;
  input [7:0] m_logical_addr_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [127:0] m_data_data_rsci_idat;
  wire [7:0] m_logical_addr_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  reg [7:0] m_logical_addr_buf_lpi_1_dfm;
  reg [127:0] m_data_data_buf_lpi_1_dfm;
  wire and_dcpl;
  wire or_dcpl_2;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_3_cse;
  wire this_val_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire [0:0] nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd52),
  .width(32'sd128)) m_data_data_rsci (
      .dat(m_data_data_rsc_dat),
      .idat(m_data_data_rsci_idat)
    );
  ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd54),
  .width(32'sd8)) m_logical_addr_rsci (
      .dat(m_logical_addr_rsc_dat),
      .idat(m_logical_addr_rsci_idat)
    );
  ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd110),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1
      #(.rscid(32'sd116)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld[0:0])
    );
  assign this_msg = {m_logical_addr_buf_lpi_1_dfm , 2'b00 , m_data_data_buf_lpi_1_dfm};
  assign or_3_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign or_dcpl_2 = and_dcpl | (~ ccs_ccore_start_rsci_idat);
  assign this_val_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk ) begin
    if ( ~ ccs_MIO_arst ) begin
      this_val <= 1'b0;
    end
    else if ( or_3_cse | this_val_mx0c1 ) begin
      this_val <= ~ this_val_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk ) begin
    if ( ~ ccs_MIO_arst ) begin
      m_logical_addr_buf_lpi_1_dfm <= 8'b00000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_logical_addr_buf_lpi_1_dfm <= m_logical_addr_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk ) begin
    if ( ~ ccs_MIO_arst ) begin
      m_data_data_buf_lpi_1_dfm <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_data_data_buf_lpi_1_dfm <= m_data_data_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk ) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_3_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_spec_StreamType_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module ActUnit_Connections_OutBlocking_spec_StreamType_Connections_SYN_PORT_Push (
  this_val, this_rdy, this_msg, m_data_data_rsc_dat, m_logical_addr_rsc_dat, ccs_ccore_start_rsc_dat,
      ccs_ccore_done_sync_vld, ccs_MIO_clk, ccs_MIO_arst
);
  output this_val;
  input this_rdy;
  output [137:0] this_msg;
  input [127:0] m_data_data_rsc_dat;
  input [7:0] m_logical_addr_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_StreamType_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_spec_StreamType_Connections_SYN_PORT_Push_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .m_data_data_rsc_dat(m_data_data_rsc_dat),
      .m_logical_addr_rsc_dat(m_logical_addr_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./ActUnit_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ActUnit_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./ActUnit_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ActUnit_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./ActUnit_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   huaixil@sat8
//  Generated date: Fri Apr  8 23:10:35 2022
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_bool_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module ActUnit_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_bool_Connections_SYN_PORT_Push_core
    (
  this_val, this_rdy, this_msg, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_val;
  reg this_val;
  input this_rdy;
  output this_msg;
  reg this_msg;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_3_cse;
  wire this_val_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire [0:0] nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  ActUnit_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd109),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  ActUnit_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1
      #(.rscid(32'sd115)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld[0:0])
    );
  assign or_3_cse = ccs_ccore_start_rsci_idat | (io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & (~ this_rdy));
  assign this_val_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk ) begin
    if ( ~ ccs_MIO_arst ) begin
      this_val <= 1'b0;
    end
    else if ( or_3_cse | this_val_mx0c1 ) begin
      this_val <= ~ this_val_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk ) begin
    if ( ~ ccs_MIO_arst ) begin
      this_msg <= 1'b0;
    end
    else if ( (~((~ io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1) | this_rdy)) | ccs_ccore_start_rsci_idat
        ) begin
      this_msg <= 1'b1;
    end
  end
  always @(posedge ccs_MIO_clk ) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_3_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_bool_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module ActUnit_Connections_OutBlocking_bool_Connections_SYN_PORT_Push (
  this_val, this_rdy, this_msg, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_val;
  input this_rdy;
  output this_msg;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  ActUnit_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_bool_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_bool_Connections_SYN_PORT_Push_core_inst (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./ActUnit_EAdd.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   huaixil@sat8
//  Generated date: Fri Apr  8 23:11:10 2022
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    EAdd
// ------------------------------------------------------------------


module ActUnit_EAdd (
  in_1_data, in_2_data, out_data
);
  input [319:0] in_1_data;
  input [319:0] in_2_data;
  output [319:0] out_data;


  wire[19:0] for_acc_17_nl;
  wire[20:0] nl_for_acc_17_nl;
  wire[19:0] for_acc_16_nl;
  wire[20:0] nl_for_acc_16_nl;
  wire[19:0] for_acc_15_nl;
  wire[20:0] nl_for_acc_15_nl;
  wire[19:0] for_acc_14_nl;
  wire[20:0] nl_for_acc_14_nl;
  wire[19:0] for_acc_13_nl;
  wire[20:0] nl_for_acc_13_nl;
  wire[19:0] for_acc_12_nl;
  wire[20:0] nl_for_acc_12_nl;
  wire[19:0] for_acc_11_nl;
  wire[20:0] nl_for_acc_11_nl;
  wire[19:0] for_acc_10_nl;
  wire[20:0] nl_for_acc_10_nl;
  wire[19:0] for_acc_9_nl;
  wire[20:0] nl_for_acc_9_nl;
  wire[19:0] for_acc_8_nl;
  wire[20:0] nl_for_acc_8_nl;
  wire[19:0] for_acc_7_nl;
  wire[20:0] nl_for_acc_7_nl;
  wire[19:0] for_acc_6_nl;
  wire[20:0] nl_for_acc_6_nl;
  wire[19:0] for_acc_5_nl;
  wire[20:0] nl_for_acc_5_nl;
  wire[19:0] for_acc_4_nl;
  wire[20:0] nl_for_acc_4_nl;
  wire[19:0] for_acc_3_nl;
  wire[20:0] nl_for_acc_3_nl;
  wire[19:0] for_acc_1_nl;
  wire[20:0] nl_for_acc_1_nl;

  // Interconnect Declarations for Component Instantiations
  assign nl_for_acc_17_nl = (in_1_data[319:300]) + (in_2_data[319:300]);
  assign for_acc_17_nl = nl_for_acc_17_nl[19:0];
  assign nl_for_acc_16_nl = (in_1_data[299:280]) + (in_2_data[299:280]);
  assign for_acc_16_nl = nl_for_acc_16_nl[19:0];
  assign nl_for_acc_15_nl = (in_1_data[279:260]) + (in_2_data[279:260]);
  assign for_acc_15_nl = nl_for_acc_15_nl[19:0];
  assign nl_for_acc_14_nl = (in_1_data[259:240]) + (in_2_data[259:240]);
  assign for_acc_14_nl = nl_for_acc_14_nl[19:0];
  assign nl_for_acc_13_nl = (in_1_data[239:220]) + (in_2_data[239:220]);
  assign for_acc_13_nl = nl_for_acc_13_nl[19:0];
  assign nl_for_acc_12_nl = (in_1_data[219:200]) + (in_2_data[219:200]);
  assign for_acc_12_nl = nl_for_acc_12_nl[19:0];
  assign nl_for_acc_11_nl = (in_1_data[199:180]) + (in_2_data[199:180]);
  assign for_acc_11_nl = nl_for_acc_11_nl[19:0];
  assign nl_for_acc_10_nl = (in_1_data[179:160]) + (in_2_data[179:160]);
  assign for_acc_10_nl = nl_for_acc_10_nl[19:0];
  assign nl_for_acc_9_nl = (in_1_data[159:140]) + (in_2_data[159:140]);
  assign for_acc_9_nl = nl_for_acc_9_nl[19:0];
  assign nl_for_acc_8_nl = (in_1_data[139:120]) + (in_2_data[139:120]);
  assign for_acc_8_nl = nl_for_acc_8_nl[19:0];
  assign nl_for_acc_7_nl = (in_1_data[119:100]) + (in_2_data[119:100]);
  assign for_acc_7_nl = nl_for_acc_7_nl[19:0];
  assign nl_for_acc_6_nl = (in_1_data[99:80]) + (in_2_data[99:80]);
  assign for_acc_6_nl = nl_for_acc_6_nl[19:0];
  assign nl_for_acc_5_nl = (in_1_data[79:60]) + (in_2_data[79:60]);
  assign for_acc_5_nl = nl_for_acc_5_nl[19:0];
  assign nl_for_acc_4_nl = (in_1_data[59:40]) + (in_2_data[59:40]);
  assign for_acc_4_nl = nl_for_acc_4_nl[19:0];
  assign nl_for_acc_3_nl = (in_1_data[39:20]) + (in_2_data[39:20]);
  assign for_acc_3_nl = nl_for_acc_3_nl[19:0];
  assign nl_for_acc_1_nl = (in_1_data[19:0]) + (in_2_data[19:0]);
  assign for_acc_1_nl = nl_for_acc_1_nl[19:0];
  assign out_data = {for_acc_17_nl , for_acc_16_nl , for_acc_15_nl , for_acc_14_nl
      , for_acc_13_nl , for_acc_12_nl , for_acc_11_nl , for_acc_10_nl , for_acc_9_nl
      , for_acc_8_nl , for_acc_7_nl , for_acc_6_nl , for_acc_5_nl , for_acc_4_nl
      , for_acc_3_nl , for_acc_1_nl};
endmodule




//------> ./ActUnit_EMul.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   huaixil@sat8
//  Generated date: Fri Apr  8 23:11:07 2022
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    EMul
// ------------------------------------------------------------------


module ActUnit_EMul (
  in_1_data, in_2_data, out_data
);
  input [319:0] in_1_data;
  input [319:0] in_2_data;
  output [319:0] out_data;


  wire[33:0] for_mul_15_nl;
  wire signed [39:0] nl_for_mul_15_nl;
  wire[33:0] for_mul_14_nl;
  wire signed [39:0] nl_for_mul_14_nl;
  wire[33:0] for_mul_13_nl;
  wire signed [39:0] nl_for_mul_13_nl;
  wire[33:0] for_mul_12_nl;
  wire signed [39:0] nl_for_mul_12_nl;
  wire[33:0] for_mul_11_nl;
  wire signed [39:0] nl_for_mul_11_nl;
  wire[33:0] for_mul_10_nl;
  wire signed [39:0] nl_for_mul_10_nl;
  wire[33:0] for_mul_9_nl;
  wire signed [39:0] nl_for_mul_9_nl;
  wire[33:0] for_mul_8_nl;
  wire signed [39:0] nl_for_mul_8_nl;
  wire[33:0] for_mul_7_nl;
  wire signed [39:0] nl_for_mul_7_nl;
  wire[33:0] for_mul_6_nl;
  wire signed [39:0] nl_for_mul_6_nl;
  wire[33:0] for_mul_5_nl;
  wire signed [39:0] nl_for_mul_5_nl;
  wire[33:0] for_mul_4_nl;
  wire signed [39:0] nl_for_mul_4_nl;
  wire[33:0] for_mul_3_nl;
  wire signed [39:0] nl_for_mul_3_nl;
  wire[33:0] for_mul_2_nl;
  wire signed [39:0] nl_for_mul_2_nl;
  wire[33:0] for_mul_1_nl;
  wire signed [39:0] nl_for_mul_1_nl;
  wire[33:0] for_mul_nl;
  wire signed [39:0] nl_for_mul_nl;

  // Interconnect Declarations for Component Instantiations
  assign nl_for_mul_15_nl = $signed((in_1_data[319:300])) * $signed((in_2_data[319:300]));
  assign for_mul_15_nl = nl_for_mul_15_nl[33:0];
  assign nl_for_mul_14_nl = $signed((in_1_data[299:280])) * $signed((in_2_data[299:280]));
  assign for_mul_14_nl = nl_for_mul_14_nl[33:0];
  assign nl_for_mul_13_nl = $signed((in_1_data[279:260])) * $signed((in_2_data[279:260]));
  assign for_mul_13_nl = nl_for_mul_13_nl[33:0];
  assign nl_for_mul_12_nl = $signed((in_1_data[259:240])) * $signed((in_2_data[259:240]));
  assign for_mul_12_nl = nl_for_mul_12_nl[33:0];
  assign nl_for_mul_11_nl = $signed((in_1_data[239:220])) * $signed((in_2_data[239:220]));
  assign for_mul_11_nl = nl_for_mul_11_nl[33:0];
  assign nl_for_mul_10_nl = $signed((in_1_data[219:200])) * $signed((in_2_data[219:200]));
  assign for_mul_10_nl = nl_for_mul_10_nl[33:0];
  assign nl_for_mul_9_nl = $signed((in_1_data[199:180])) * $signed((in_2_data[199:180]));
  assign for_mul_9_nl = nl_for_mul_9_nl[33:0];
  assign nl_for_mul_8_nl = $signed((in_1_data[179:160])) * $signed((in_2_data[179:160]));
  assign for_mul_8_nl = nl_for_mul_8_nl[33:0];
  assign nl_for_mul_7_nl = $signed((in_1_data[159:140])) * $signed((in_2_data[159:140]));
  assign for_mul_7_nl = nl_for_mul_7_nl[33:0];
  assign nl_for_mul_6_nl = $signed((in_1_data[139:120])) * $signed((in_2_data[139:120]));
  assign for_mul_6_nl = nl_for_mul_6_nl[33:0];
  assign nl_for_mul_5_nl = $signed((in_1_data[119:100])) * $signed((in_2_data[119:100]));
  assign for_mul_5_nl = nl_for_mul_5_nl[33:0];
  assign nl_for_mul_4_nl = $signed((in_1_data[99:80])) * $signed((in_2_data[99:80]));
  assign for_mul_4_nl = nl_for_mul_4_nl[33:0];
  assign nl_for_mul_3_nl = $signed((in_1_data[79:60])) * $signed((in_2_data[79:60]));
  assign for_mul_3_nl = nl_for_mul_3_nl[33:0];
  assign nl_for_mul_2_nl = $signed((in_1_data[59:40])) * $signed((in_2_data[59:40]));
  assign for_mul_2_nl = nl_for_mul_2_nl[33:0];
  assign nl_for_mul_1_nl = $signed((in_1_data[39:20])) * $signed((in_2_data[39:20]));
  assign for_mul_1_nl = nl_for_mul_1_nl[33:0];
  assign nl_for_mul_nl = $signed((in_1_data[19:0])) * $signed((in_2_data[19:0]));
  assign for_mul_nl = nl_for_mul_nl[33:0];
  assign out_data = {(readslicef_34_20_14(for_mul_15_nl)) , (readslicef_34_20_14(for_mul_14_nl))
      , (readslicef_34_20_14(for_mul_13_nl)) , (readslicef_34_20_14(for_mul_12_nl))
      , (readslicef_34_20_14(for_mul_11_nl)) , (readslicef_34_20_14(for_mul_10_nl))
      , (readslicef_34_20_14(for_mul_9_nl)) , (readslicef_34_20_14(for_mul_8_nl))
      , (readslicef_34_20_14(for_mul_7_nl)) , (readslicef_34_20_14(for_mul_6_nl))
      , (readslicef_34_20_14(for_mul_5_nl)) , (readslicef_34_20_14(for_mul_4_nl))
      , (readslicef_34_20_14(for_mul_3_nl)) , (readslicef_34_20_14(for_mul_2_nl))
      , (readslicef_34_20_14(for_mul_1_nl)) , (readslicef_34_20_14(for_mul_nl))};

  function automatic [19:0] readslicef_34_20_14;
    input [33:0] vector;
    reg [33:0] tmp;
  begin
    tmp = vector >> 14;
    readslicef_34_20_14 = tmp[19:0];
  end
  endfunction

endmodule




//------> ./ActUnit_Sigmoid.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   huaixil@sat8
//  Generated date: Fri Apr  8 23:11:04 2022
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Sigmoid
// ------------------------------------------------------------------


module ActUnit_Sigmoid (
  in_data, out_data
);
  input [319:0] in_data;
  output [319:0] out_data;


  // Interconnect Declarations
  wire and_dcpl;
  wire and_dcpl_1;
  wire and_dcpl_2;
  wire and_dcpl_3;
  wire and_dcpl_4;
  wire and_dcpl_5;
  wire and_dcpl_6;
  wire and_dcpl_7;
  wire and_dcpl_8;
  wire and_dcpl_9;
  wire and_dcpl_10;
  wire and_dcpl_11;
  wire and_dcpl_12;
  wire and_dcpl_13;
  wire and_dcpl_14;
  wire and_dcpl_15;
  wire and_dcpl_16;
  wire and_dcpl_17;
  wire and_dcpl_18;
  wire and_dcpl_19;
  wire and_dcpl_20;
  wire and_dcpl_21;
  wire and_dcpl_22;
  wire and_dcpl_23;
  wire and_dcpl_24;
  wire and_dcpl_25;
  wire and_dcpl_26;
  wire and_dcpl_27;
  wire and_dcpl_28;
  wire and_dcpl_29;
  wire and_dcpl_30;
  wire and_dcpl_31;
  wire [9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_16_mx0w1;
  wire [10:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_16_mx0w1;
  wire [9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_31_mx0w1;
  wire [10:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_31_mx0w1;
  wire [9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_30_mx0w1;
  wire [10:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_30_mx0w1;
  wire [9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_29_mx0w1;
  wire [10:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_29_mx0w1;
  wire [9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_28_mx0w1;
  wire [10:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_28_mx0w1;
  wire [9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_27_mx0w1;
  wire [10:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_27_mx0w1;
  wire [9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_26_mx0w1;
  wire [10:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_26_mx0w1;
  wire [9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_25_mx0w1;
  wire [10:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_25_mx0w1;
  wire [9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_24_mx0w1;
  wire [10:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_24_mx0w1;
  wire [9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_23_mx0w1;
  wire [10:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_23_mx0w1;
  wire [9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_22_mx0w1;
  wire [10:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_22_mx0w1;
  wire [9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_21_mx0w1;
  wire [10:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_21_mx0w1;
  wire [9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_20_mx0w1;
  wire [10:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_20_mx0w1;
  wire [9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_19_mx0w1;
  wire [10:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_19_mx0w1;
  wire [9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_18_mx0w1;
  wire [10:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_18_mx0w1;
  wire [9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_17_mx0w1;
  wire [10:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_17_mx0w1;
  wire [17:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_16;
  wire [17:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_17;
  wire [17:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_18;
  wire [17:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_19;
  wire [17:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_20;
  wire [17:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_21;
  wire [17:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_22;
  wire [17:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_23;
  wire [17:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_24;
  wire [17:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_25;
  wire [17:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_26;
  wire [17:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_27;
  wire [17:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_28;
  wire [17:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_29;
  wire [17:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_30;
  wire [17:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_31;
  wire [19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_1_mx0;
  wire [19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_2_mx0;
  wire [19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_3_mx0;
  wire [19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_4_mx0;
  wire [19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_5_mx0;
  wire [19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_6_mx0;
  wire [19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_7_mx0;
  wire [19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_8_mx0;
  wire [19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_9_mx0;
  wire [19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_10_mx0;
  wire [19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_11_mx0;
  wire [19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_12_mx0;
  wire [19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_13_mx0;
  wire [19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_14_mx0;
  wire [19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_15_mx0;
  wire [19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_mx0;
  wire [13:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_itm_19_6_1;
  wire [13:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_1_itm_19_6_1;
  wire [13:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_2_itm_19_6_1;
  wire [13:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_3_itm_19_6_1;
  wire [13:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_4_itm_19_6_1;
  wire [13:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_5_itm_19_6_1;
  wire [13:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_6_itm_19_6_1;
  wire [13:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_7_itm_19_6_1;
  wire [13:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_8_itm_19_6_1;
  wire [13:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_9_itm_19_6_1;
  wire [13:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_10_itm_19_6_1;
  wire [13:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_11_itm_19_6_1;
  wire [13:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_12_itm_19_6_1;
  wire [13:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_13_itm_19_6_1;
  wire [13:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_14_itm_19_6_1;
  wire [13:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_15_itm_19_6_1;
  wire [12:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_15_itm_25_13;
  wire [12:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_14_itm_25_13;
  wire [12:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_13_itm_25_13;
  wire [12:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_12_itm_25_13;
  wire [12:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_11_itm_25_13;
  wire [12:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_10_itm_25_13;
  wire [12:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_9_itm_25_13;
  wire [12:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_8_itm_25_13;
  wire [12:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_7_itm_25_13;
  wire [12:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_6_itm_25_13;
  wire [12:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_5_itm_25_13;
  wire [12:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_4_itm_25_13;
  wire [12:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_3_itm_25_13;
  wire [12:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_2_itm_25_13;
  wire [12:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_1_itm_25_13;
  wire [12:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_itm_25_13;
  wire ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_15_itm_5_1;
  wire ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_14_itm_5_1;
  wire ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_13_itm_5_1;
  wire ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_12_itm_5_1;
  wire ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_11_itm_5_1;
  wire ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_10_itm_5_1;
  wire ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_9_itm_5_1;
  wire ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_8_itm_5_1;
  wire ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_7_itm_5_1;
  wire ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_6_itm_5_1;
  wire ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_5_itm_5_1;
  wire ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_4_itm_5_1;
  wire ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_3_itm_5_1;
  wire ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_2_itm_5_1;
  wire ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_1_itm_5_1;
  wire ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_itm_5_1;

  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_48_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_15_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_47_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_16_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_49_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_14_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_46_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_17_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_50_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_13_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_45_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_18_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_51_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_12_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_44_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_19_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_52_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_11_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_43_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_20_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_53_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_10_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_42_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_21_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_54_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_9_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_41_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_22_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_55_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_8_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_40_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_23_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_56_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_7_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_39_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_24_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_57_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_6_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_38_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_25_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_58_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_5_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_37_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_26_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_59_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_4_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_36_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_27_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_60_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_3_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_35_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_28_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_61_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_2_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_34_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_29_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_62_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_1_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_33_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_30_nl;
  wire[9:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_63_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_31_nl;
  wire[3:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_32_nl;
  wire[19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_nl;
  wire[20:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_nl;
  wire[8:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_1_nl;
  wire[19:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_nl;
  wire[20:0] nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_30_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_16_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_31_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_nl;
  wire[19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_1_nl;
  wire[20:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_1_nl;
  wire[8:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_3_nl;
  wire[19:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_1_nl;
  wire[20:0] nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_1_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_28_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_17_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_29_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_1_nl;
  wire[19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_2_nl;
  wire[20:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_2_nl;
  wire[8:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_5_nl;
  wire[19:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_2_nl;
  wire[20:0] nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_2_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_26_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_18_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_27_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_2_nl;
  wire[19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_3_nl;
  wire[20:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_3_nl;
  wire[8:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_7_nl;
  wire[19:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_3_nl;
  wire[20:0] nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_3_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_24_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_19_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_25_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_3_nl;
  wire[19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_4_nl;
  wire[20:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_4_nl;
  wire[8:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_9_nl;
  wire[19:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_4_nl;
  wire[20:0] nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_4_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_22_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_20_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_23_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_4_nl;
  wire[19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_5_nl;
  wire[20:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_5_nl;
  wire[8:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_11_nl;
  wire[19:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_5_nl;
  wire[20:0] nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_5_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_20_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_21_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_21_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_5_nl;
  wire[19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_6_nl;
  wire[20:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_6_nl;
  wire[8:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_13_nl;
  wire[19:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_6_nl;
  wire[20:0] nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_6_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_18_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_22_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_19_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_6_nl;
  wire[19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_7_nl;
  wire[20:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_7_nl;
  wire[8:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_15_nl;
  wire[19:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_7_nl;
  wire[20:0] nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_7_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_16_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_23_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_17_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_7_nl;
  wire[19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_8_nl;
  wire[20:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_8_nl;
  wire[8:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_17_nl;
  wire[19:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_8_nl;
  wire[20:0] nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_8_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_14_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_24_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_15_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_8_nl;
  wire[19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_9_nl;
  wire[20:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_9_nl;
  wire[8:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_19_nl;
  wire[19:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_9_nl;
  wire[20:0] nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_9_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_12_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_25_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_13_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_9_nl;
  wire[19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_10_nl;
  wire[20:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_10_nl;
  wire[8:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_21_nl;
  wire[19:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_10_nl;
  wire[20:0] nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_10_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_10_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_26_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_11_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_10_nl;
  wire[19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_11_nl;
  wire[20:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_11_nl;
  wire[8:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_23_nl;
  wire[19:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_11_nl;
  wire[20:0] nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_11_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_8_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_27_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_9_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_11_nl;
  wire[19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_12_nl;
  wire[20:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_12_nl;
  wire[8:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_25_nl;
  wire[19:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_12_nl;
  wire[20:0] nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_12_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_6_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_28_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_7_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_12_nl;
  wire[19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_13_nl;
  wire[20:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_13_nl;
  wire[8:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_27_nl;
  wire[19:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_13_nl;
  wire[20:0] nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_13_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_4_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_29_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_5_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_13_nl;
  wire[19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_14_nl;
  wire[20:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_14_nl;
  wire[8:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_29_nl;
  wire[19:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_14_nl;
  wire[20:0] nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_14_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_2_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_30_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_3_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_14_nl;
  wire[19:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_15_nl;
  wire[20:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_15_nl;
  wire[8:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_31_nl;
  wire[19:0] operator_20_0_false_AC_TRN_AC_WRAP_acc_15_nl;
  wire[20:0] nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_15_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_31_nl;
  wire[9:0] operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_1_nl;
  wire[0:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_15_nl;
  wire[7:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_30_nl;
  wire[25:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_15_nl;
  wire[29:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_15_nl;
  wire[7:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_28_nl;
  wire[25:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_14_nl;
  wire[29:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_14_nl;
  wire[7:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_26_nl;
  wire[25:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_13_nl;
  wire[29:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_13_nl;
  wire[7:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_24_nl;
  wire[25:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_12_nl;
  wire[29:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_12_nl;
  wire[7:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_22_nl;
  wire[25:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_11_nl;
  wire[29:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_11_nl;
  wire[7:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_20_nl;
  wire[25:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_10_nl;
  wire[29:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_10_nl;
  wire[7:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_18_nl;
  wire[25:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_9_nl;
  wire[29:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_9_nl;
  wire[7:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_16_nl;
  wire[25:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_8_nl;
  wire[29:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_8_nl;
  wire[7:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_14_nl;
  wire[25:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_7_nl;
  wire[29:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_7_nl;
  wire[7:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_12_nl;
  wire[25:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_6_nl;
  wire[29:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_6_nl;
  wire[7:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_10_nl;
  wire[25:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_5_nl;
  wire[29:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_5_nl;
  wire[7:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_8_nl;
  wire[25:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_4_nl;
  wire[29:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_4_nl;
  wire[7:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_6_nl;
  wire[25:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_3_nl;
  wire[29:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_3_nl;
  wire[7:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_4_nl;
  wire[25:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_2_nl;
  wire[29:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_2_nl;
  wire[7:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_2_nl;
  wire[25:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_1_nl;
  wire[29:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_1_nl;
  wire[7:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_nl;
  wire[25:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_nl;
  wire[29:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_nl;
  wire[5:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_15_nl;
  wire[6:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_15_nl;
  wire[5:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_14_nl;
  wire[6:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_14_nl;
  wire[5:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_13_nl;
  wire[6:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_13_nl;
  wire[5:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_12_nl;
  wire[6:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_12_nl;
  wire[5:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_11_nl;
  wire[6:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_11_nl;
  wire[5:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_10_nl;
  wire[6:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_10_nl;
  wire[5:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_9_nl;
  wire[6:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_9_nl;
  wire[5:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_8_nl;
  wire[6:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_8_nl;
  wire[5:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_7_nl;
  wire[6:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_7_nl;
  wire[5:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_6_nl;
  wire[6:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_6_nl;
  wire[5:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_5_nl;
  wire[6:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_5_nl;
  wire[5:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_4_nl;
  wire[6:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_4_nl;
  wire[5:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_3_nl;
  wire[6:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_3_nl;
  wire[5:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_2_nl;
  wire[6:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_2_nl;
  wire[5:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_1_nl;
  wire[6:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_1_nl;
  wire[5:0] ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_nl;
  wire[6:0] nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_nl;

  // Interconnect Declarations for Component Instantiations
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_48_nl
      = MUX_v_10_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_15_itm_19_6_1[13:4]),
      ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_16_mx0w1,
      and_dcpl_31);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_nl
      = MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_48_nl,
      10'b1111111111, and_dcpl_30);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_47_nl
      = MUX_v_4_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_15_itm_19_6_1[3:0]),
      (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_16[9:6]),
      and_dcpl_31);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_15_nl
      = MUX_v_4_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_47_nl,
      4'b1111, and_dcpl_30);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_49_nl
      = MUX_v_10_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_14_itm_19_6_1[13:4]),
      ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_31_mx0w1,
      and_dcpl_29);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_16_nl
      = MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_49_nl,
      10'b1111111111, and_dcpl_28);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_46_nl
      = MUX_v_4_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_14_itm_19_6_1[3:0]),
      (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_17[9:6]),
      and_dcpl_29);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_14_nl
      = MUX_v_4_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_46_nl,
      4'b1111, and_dcpl_28);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_50_nl
      = MUX_v_10_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_13_itm_19_6_1[13:4]),
      ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_30_mx0w1,
      and_dcpl_27);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_17_nl
      = MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_50_nl,
      10'b1111111111, and_dcpl_26);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_45_nl
      = MUX_v_4_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_13_itm_19_6_1[3:0]),
      (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_18[9:6]),
      and_dcpl_27);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_13_nl
      = MUX_v_4_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_45_nl,
      4'b1111, and_dcpl_26);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_51_nl
      = MUX_v_10_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_12_itm_19_6_1[13:4]),
      ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_29_mx0w1,
      and_dcpl_25);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_18_nl
      = MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_51_nl,
      10'b1111111111, and_dcpl_24);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_44_nl
      = MUX_v_4_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_12_itm_19_6_1[3:0]),
      (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_19[9:6]),
      and_dcpl_25);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_12_nl
      = MUX_v_4_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_44_nl,
      4'b1111, and_dcpl_24);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_52_nl
      = MUX_v_10_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_11_itm_19_6_1[13:4]),
      ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_28_mx0w1,
      and_dcpl_23);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_19_nl
      = MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_52_nl,
      10'b1111111111, and_dcpl_22);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_43_nl
      = MUX_v_4_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_11_itm_19_6_1[3:0]),
      (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_20[9:6]),
      and_dcpl_23);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_11_nl
      = MUX_v_4_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_43_nl,
      4'b1111, and_dcpl_22);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_53_nl
      = MUX_v_10_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_10_itm_19_6_1[13:4]),
      ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_27_mx0w1,
      and_dcpl_21);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_20_nl
      = MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_53_nl,
      10'b1111111111, and_dcpl_20);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_42_nl
      = MUX_v_4_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_10_itm_19_6_1[3:0]),
      (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_21[9:6]),
      and_dcpl_21);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_10_nl
      = MUX_v_4_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_42_nl,
      4'b1111, and_dcpl_20);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_54_nl
      = MUX_v_10_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_9_itm_19_6_1[13:4]),
      ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_26_mx0w1,
      and_dcpl_19);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_21_nl
      = MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_54_nl,
      10'b1111111111, and_dcpl_18);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_41_nl
      = MUX_v_4_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_9_itm_19_6_1[3:0]), (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_22[9:6]),
      and_dcpl_19);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_9_nl
      = MUX_v_4_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_41_nl,
      4'b1111, and_dcpl_18);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_55_nl
      = MUX_v_10_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_8_itm_19_6_1[13:4]),
      ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_25_mx0w1,
      and_dcpl_17);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_22_nl
      = MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_55_nl,
      10'b1111111111, and_dcpl_16);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_40_nl
      = MUX_v_4_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_8_itm_19_6_1[3:0]), (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_23[9:6]),
      and_dcpl_17);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_8_nl
      = MUX_v_4_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_40_nl,
      4'b1111, and_dcpl_16);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_56_nl
      = MUX_v_10_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_7_itm_19_6_1[13:4]),
      ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_24_mx0w1,
      and_dcpl_15);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_23_nl
      = MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_56_nl,
      10'b1111111111, and_dcpl_14);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_39_nl
      = MUX_v_4_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_7_itm_19_6_1[3:0]), (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_24[9:6]),
      and_dcpl_15);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_7_nl
      = MUX_v_4_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_39_nl,
      4'b1111, and_dcpl_14);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_57_nl
      = MUX_v_10_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_6_itm_19_6_1[13:4]),
      ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_23_mx0w1,
      and_dcpl_13);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_24_nl
      = MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_57_nl,
      10'b1111111111, and_dcpl_12);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_38_nl
      = MUX_v_4_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_6_itm_19_6_1[3:0]), (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_25[9:6]),
      and_dcpl_13);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_6_nl
      = MUX_v_4_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_38_nl,
      4'b1111, and_dcpl_12);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_58_nl
      = MUX_v_10_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_5_itm_19_6_1[13:4]),
      ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_22_mx0w1,
      and_dcpl_11);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_25_nl
      = MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_58_nl,
      10'b1111111111, and_dcpl_10);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_37_nl
      = MUX_v_4_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_5_itm_19_6_1[3:0]), (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_26[9:6]),
      and_dcpl_11);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_5_nl
      = MUX_v_4_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_37_nl,
      4'b1111, and_dcpl_10);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_59_nl
      = MUX_v_10_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_4_itm_19_6_1[13:4]),
      ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_21_mx0w1,
      and_dcpl_9);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_26_nl
      = MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_59_nl,
      10'b1111111111, and_dcpl_8);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_36_nl
      = MUX_v_4_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_4_itm_19_6_1[3:0]), (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_27[9:6]),
      and_dcpl_9);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_4_nl
      = MUX_v_4_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_36_nl,
      4'b1111, and_dcpl_8);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_60_nl
      = MUX_v_10_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_3_itm_19_6_1[13:4]),
      ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_20_mx0w1,
      and_dcpl_7);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_27_nl
      = MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_60_nl,
      10'b1111111111, and_dcpl_6);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_35_nl
      = MUX_v_4_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_3_itm_19_6_1[3:0]), (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_28[9:6]),
      and_dcpl_7);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_3_nl
      = MUX_v_4_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_35_nl,
      4'b1111, and_dcpl_6);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_61_nl
      = MUX_v_10_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_2_itm_19_6_1[13:4]),
      ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_19_mx0w1,
      and_dcpl_5);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_28_nl
      = MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_61_nl,
      10'b1111111111, and_dcpl_4);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_34_nl
      = MUX_v_4_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_2_itm_19_6_1[3:0]), (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_29[9:6]),
      and_dcpl_5);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_2_nl
      = MUX_v_4_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_34_nl,
      4'b1111, and_dcpl_4);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_62_nl
      = MUX_v_10_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_1_itm_19_6_1[13:4]),
      ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_18_mx0w1,
      and_dcpl_3);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_29_nl
      = MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_62_nl,
      10'b1111111111, and_dcpl_2);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_33_nl
      = MUX_v_4_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_1_itm_19_6_1[3:0]), (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_30[9:6]),
      and_dcpl_3);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_1_nl
      = MUX_v_4_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_33_nl,
      4'b1111, and_dcpl_2);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_63_nl
      = MUX_v_10_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_itm_19_6_1[13:4]), ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_17_mx0w1,
      and_dcpl_1);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_30_nl
      = MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_63_nl,
      10'b1111111111, and_dcpl);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_32_nl
      = MUX_v_4_2_2((operator_20_0_false_AC_TRN_AC_WRAP_acc_itm_19_6_1[3:0]), (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_31[9:6]),
      and_dcpl_1);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_31_nl
      = MUX_v_4_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_32_nl,
      4'b1111, and_dcpl);
  assign out_data = {6'b000000 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_nl
      , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_15_nl
      , 6'b000000 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_16_nl
      , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_14_nl
      , 6'b000000 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_17_nl
      , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_13_nl
      , 6'b000000 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_18_nl
      , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_12_nl
      , 6'b000000 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_19_nl
      , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_11_nl
      , 6'b000000 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_20_nl
      , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_10_nl
      , 6'b000000 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_21_nl
      , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_9_nl
      , 6'b000000 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_22_nl
      , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_8_nl
      , 6'b000000 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_23_nl
      , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_7_nl
      , 6'b000000 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_24_nl
      , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_6_nl
      , 6'b000000 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_25_nl
      , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_5_nl
      , 6'b000000 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_26_nl
      , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_4_nl
      , 6'b000000 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_27_nl
      , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_3_nl
      , 6'b000000 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_28_nl
      , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_2_nl
      , 6'b000000 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_29_nl
      , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_1_nl
      , 6'b000000 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_30_nl
      , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_or_31_nl};
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_nl
      = conv_u2u_19_20(~ (in_data[18:0])) + 20'b00000000000000000001;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_nl[19:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_1_mx0
      = MUX_v_20_2_2(({1'b0 , (in_data[18:0])}), ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_nl,
      in_data[19]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_1_nl
      = MUX_v_9_8_2(9'b000000001, 9'b010011100, 9'b100011110, 9'b101111010, 9'b110110100,
      9'b111010110, 9'b111101001, 9'b111110100, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_itm_25_13[12:10]);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_17_mx0w1
      = conv_u2u_8_10(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_31[17:10])
      + ({1'b1 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_1_nl});
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_17_mx0w1
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_17_mx0w1[9:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_16_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_30_nl
      = ~(MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_17_mx0w1,
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_16_nl));
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_31_nl
      = ~(MUX_v_10_2_2((ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_31[9:0]),
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_nl));
  assign nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_nl = ({operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_30_nl
      , operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_31_nl})
      + 20'b00000000000000000001;
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_nl = nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_nl[19:0];
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_itm_19_6_1 = readslicef_20_14_6(operator_20_0_false_AC_TRN_AC_WRAP_acc_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_1_nl
      = conv_u2u_19_20(~ (in_data[38:20])) + 20'b00000000000000000001;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_1_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_1_nl[19:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_2_mx0
      = MUX_v_20_2_2(({1'b0 , (in_data[38:20])}), ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_1_nl,
      in_data[39]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_3_nl
      = MUX_v_9_8_2(9'b000000001, 9'b010011100, 9'b100011110, 9'b101111010, 9'b110110100,
      9'b111010110, 9'b111101001, 9'b111110100, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_1_itm_25_13[12:10]);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_18_mx0w1
      = conv_u2u_8_10(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_30[17:10])
      + ({1'b1 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_3_nl});
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_18_mx0w1
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_18_mx0w1[9:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_17_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_1_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_28_nl
      = ~(MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_18_mx0w1,
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_17_nl));
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_1_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_1_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_29_nl
      = ~(MUX_v_10_2_2((ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_30[9:0]),
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_1_nl));
  assign nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_1_nl = ({operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_28_nl
      , operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_29_nl})
      + 20'b00000000000000000001;
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_1_nl = nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_1_nl[19:0];
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_1_itm_19_6_1 = readslicef_20_14_6(operator_20_0_false_AC_TRN_AC_WRAP_acc_1_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_2_nl
      = conv_u2u_19_20(~ (in_data[58:40])) + 20'b00000000000000000001;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_2_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_2_nl[19:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_3_mx0
      = MUX_v_20_2_2(({1'b0 , (in_data[58:40])}), ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_2_nl,
      in_data[59]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_5_nl
      = MUX_v_9_8_2(9'b000000001, 9'b010011100, 9'b100011110, 9'b101111010, 9'b110110100,
      9'b111010110, 9'b111101001, 9'b111110100, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_2_itm_25_13[12:10]);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_19_mx0w1
      = conv_u2u_8_10(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_29[17:10])
      + ({1'b1 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_5_nl});
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_19_mx0w1
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_19_mx0w1[9:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_18_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_2_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_26_nl
      = ~(MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_19_mx0w1,
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_18_nl));
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_2_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_2_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_27_nl
      = ~(MUX_v_10_2_2((ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_29[9:0]),
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_2_nl));
  assign nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_2_nl = ({operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_26_nl
      , operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_27_nl})
      + 20'b00000000000000000001;
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_2_nl = nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_2_nl[19:0];
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_2_itm_19_6_1 = readslicef_20_14_6(operator_20_0_false_AC_TRN_AC_WRAP_acc_2_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_3_nl
      = conv_u2u_19_20(~ (in_data[78:60])) + 20'b00000000000000000001;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_3_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_3_nl[19:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_4_mx0
      = MUX_v_20_2_2(({1'b0 , (in_data[78:60])}), ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_3_nl,
      in_data[79]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_7_nl
      = MUX_v_9_8_2(9'b000000001, 9'b010011100, 9'b100011110, 9'b101111010, 9'b110110100,
      9'b111010110, 9'b111101001, 9'b111110100, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_3_itm_25_13[12:10]);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_20_mx0w1
      = conv_u2u_8_10(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_28[17:10])
      + ({1'b1 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_7_nl});
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_20_mx0w1
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_20_mx0w1[9:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_19_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_3_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_24_nl
      = ~(MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_20_mx0w1,
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_19_nl));
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_3_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_3_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_25_nl
      = ~(MUX_v_10_2_2((ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_28[9:0]),
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_3_nl));
  assign nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_3_nl = ({operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_24_nl
      , operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_25_nl})
      + 20'b00000000000000000001;
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_3_nl = nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_3_nl[19:0];
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_3_itm_19_6_1 = readslicef_20_14_6(operator_20_0_false_AC_TRN_AC_WRAP_acc_3_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_4_nl
      = conv_u2u_19_20(~ (in_data[98:80])) + 20'b00000000000000000001;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_4_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_4_nl[19:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_5_mx0
      = MUX_v_20_2_2(({1'b0 , (in_data[98:80])}), ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_4_nl,
      in_data[99]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_9_nl
      = MUX_v_9_8_2(9'b000000001, 9'b010011100, 9'b100011110, 9'b101111010, 9'b110110100,
      9'b111010110, 9'b111101001, 9'b111110100, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_4_itm_25_13[12:10]);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_21_mx0w1
      = conv_u2u_8_10(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_27[17:10])
      + ({1'b1 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_9_nl});
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_21_mx0w1
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_21_mx0w1[9:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_20_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_4_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_22_nl
      = ~(MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_21_mx0w1,
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_20_nl));
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_4_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_4_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_23_nl
      = ~(MUX_v_10_2_2((ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_27[9:0]),
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_4_nl));
  assign nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_4_nl = ({operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_22_nl
      , operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_23_nl})
      + 20'b00000000000000000001;
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_4_nl = nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_4_nl[19:0];
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_4_itm_19_6_1 = readslicef_20_14_6(operator_20_0_false_AC_TRN_AC_WRAP_acc_4_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_5_nl
      = conv_u2u_19_20(~ (in_data[118:100])) + 20'b00000000000000000001;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_5_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_5_nl[19:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_6_mx0
      = MUX_v_20_2_2(({1'b0 , (in_data[118:100])}), ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_5_nl,
      in_data[119]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_11_nl
      = MUX_v_9_8_2(9'b000000001, 9'b010011100, 9'b100011110, 9'b101111010, 9'b110110100,
      9'b111010110, 9'b111101001, 9'b111110100, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_5_itm_25_13[12:10]);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_22_mx0w1
      = conv_u2u_8_10(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_26[17:10])
      + ({1'b1 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_11_nl});
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_22_mx0w1
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_22_mx0w1[9:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_21_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_5_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_20_nl
      = ~(MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_22_mx0w1,
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_21_nl));
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_5_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_5_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_21_nl
      = ~(MUX_v_10_2_2((ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_26[9:0]),
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_5_nl));
  assign nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_5_nl = ({operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_20_nl
      , operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_21_nl})
      + 20'b00000000000000000001;
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_5_nl = nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_5_nl[19:0];
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_5_itm_19_6_1 = readslicef_20_14_6(operator_20_0_false_AC_TRN_AC_WRAP_acc_5_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_6_nl
      = conv_u2u_19_20(~ (in_data[138:120])) + 20'b00000000000000000001;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_6_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_6_nl[19:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_7_mx0
      = MUX_v_20_2_2(({1'b0 , (in_data[138:120])}), ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_6_nl,
      in_data[139]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_13_nl
      = MUX_v_9_8_2(9'b000000001, 9'b010011100, 9'b100011110, 9'b101111010, 9'b110110100,
      9'b111010110, 9'b111101001, 9'b111110100, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_6_itm_25_13[12:10]);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_23_mx0w1
      = conv_u2u_8_10(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_25[17:10])
      + ({1'b1 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_13_nl});
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_23_mx0w1
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_23_mx0w1[9:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_22_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_6_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_18_nl
      = ~(MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_23_mx0w1,
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_22_nl));
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_6_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_6_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_19_nl
      = ~(MUX_v_10_2_2((ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_25[9:0]),
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_6_nl));
  assign nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_6_nl = ({operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_18_nl
      , operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_19_nl})
      + 20'b00000000000000000001;
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_6_nl = nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_6_nl[19:0];
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_6_itm_19_6_1 = readslicef_20_14_6(operator_20_0_false_AC_TRN_AC_WRAP_acc_6_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_7_nl
      = conv_u2u_19_20(~ (in_data[158:140])) + 20'b00000000000000000001;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_7_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_7_nl[19:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_8_mx0
      = MUX_v_20_2_2(({1'b0 , (in_data[158:140])}), ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_7_nl,
      in_data[159]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_15_nl
      = MUX_v_9_8_2(9'b000000001, 9'b010011100, 9'b100011110, 9'b101111010, 9'b110110100,
      9'b111010110, 9'b111101001, 9'b111110100, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_7_itm_25_13[12:10]);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_24_mx0w1
      = conv_u2u_8_10(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_24[17:10])
      + ({1'b1 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_15_nl});
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_24_mx0w1
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_24_mx0w1[9:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_23_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_7_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_16_nl
      = ~(MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_24_mx0w1,
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_23_nl));
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_7_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_7_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_17_nl
      = ~(MUX_v_10_2_2((ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_24[9:0]),
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_7_nl));
  assign nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_7_nl = ({operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_16_nl
      , operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_17_nl})
      + 20'b00000000000000000001;
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_7_nl = nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_7_nl[19:0];
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_7_itm_19_6_1 = readslicef_20_14_6(operator_20_0_false_AC_TRN_AC_WRAP_acc_7_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_8_nl
      = conv_u2u_19_20(~ (in_data[178:160])) + 20'b00000000000000000001;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_8_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_8_nl[19:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_9_mx0
      = MUX_v_20_2_2(({1'b0 , (in_data[178:160])}), ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_8_nl,
      in_data[179]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_17_nl
      = MUX_v_9_8_2(9'b000000001, 9'b010011100, 9'b100011110, 9'b101111010, 9'b110110100,
      9'b111010110, 9'b111101001, 9'b111110100, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_8_itm_25_13[12:10]);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_25_mx0w1
      = conv_u2u_8_10(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_23[17:10])
      + ({1'b1 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_17_nl});
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_25_mx0w1
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_25_mx0w1[9:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_24_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_8_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_14_nl
      = ~(MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_25_mx0w1,
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_24_nl));
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_8_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_8_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_15_nl
      = ~(MUX_v_10_2_2((ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_23[9:0]),
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_8_nl));
  assign nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_8_nl = ({operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_14_nl
      , operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_15_nl})
      + 20'b00000000000000000001;
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_8_nl = nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_8_nl[19:0];
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_8_itm_19_6_1 = readslicef_20_14_6(operator_20_0_false_AC_TRN_AC_WRAP_acc_8_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_9_nl
      = conv_u2u_19_20(~ (in_data[198:180])) + 20'b00000000000000000001;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_9_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_9_nl[19:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_10_mx0
      = MUX_v_20_2_2(({1'b0 , (in_data[198:180])}), ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_9_nl,
      in_data[199]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_19_nl
      = MUX_v_9_8_2(9'b000000001, 9'b010011100, 9'b100011110, 9'b101111010, 9'b110110100,
      9'b111010110, 9'b111101001, 9'b111110100, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_9_itm_25_13[12:10]);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_26_mx0w1
      = conv_u2u_8_10(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_22[17:10])
      + ({1'b1 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_19_nl});
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_26_mx0w1
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_26_mx0w1[9:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_25_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_9_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_12_nl
      = ~(MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_26_mx0w1,
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_25_nl));
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_9_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_9_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_13_nl
      = ~(MUX_v_10_2_2((ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_22[9:0]),
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_9_nl));
  assign nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_9_nl = ({operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_12_nl
      , operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_13_nl})
      + 20'b00000000000000000001;
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_9_nl = nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_9_nl[19:0];
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_9_itm_19_6_1 = readslicef_20_14_6(operator_20_0_false_AC_TRN_AC_WRAP_acc_9_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_10_nl
      = conv_u2u_19_20(~ (in_data[218:200])) + 20'b00000000000000000001;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_10_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_10_nl[19:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_11_mx0
      = MUX_v_20_2_2(({1'b0 , (in_data[218:200])}), ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_10_nl,
      in_data[219]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_21_nl
      = MUX_v_9_8_2(9'b000000001, 9'b010011100, 9'b100011110, 9'b101111010, 9'b110110100,
      9'b111010110, 9'b111101001, 9'b111110100, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_10_itm_25_13[12:10]);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_27_mx0w1
      = conv_u2u_8_10(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_21[17:10])
      + ({1'b1 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_21_nl});
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_27_mx0w1
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_27_mx0w1[9:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_26_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_10_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_10_nl
      = ~(MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_27_mx0w1,
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_26_nl));
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_10_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_10_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_11_nl
      = ~(MUX_v_10_2_2((ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_21[9:0]),
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_10_nl));
  assign nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_10_nl = ({operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_10_nl
      , operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_11_nl})
      + 20'b00000000000000000001;
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_10_nl = nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_10_nl[19:0];
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_10_itm_19_6_1 = readslicef_20_14_6(operator_20_0_false_AC_TRN_AC_WRAP_acc_10_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_11_nl
      = conv_u2u_19_20(~ (in_data[238:220])) + 20'b00000000000000000001;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_11_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_11_nl[19:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_12_mx0
      = MUX_v_20_2_2(({1'b0 , (in_data[238:220])}), ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_11_nl,
      in_data[239]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_23_nl
      = MUX_v_9_8_2(9'b000000001, 9'b010011100, 9'b100011110, 9'b101111010, 9'b110110100,
      9'b111010110, 9'b111101001, 9'b111110100, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_11_itm_25_13[12:10]);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_28_mx0w1
      = conv_u2u_8_10(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_20[17:10])
      + ({1'b1 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_23_nl});
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_28_mx0w1
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_28_mx0w1[9:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_27_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_11_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_8_nl
      = ~(MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_28_mx0w1,
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_27_nl));
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_11_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_11_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_9_nl
      = ~(MUX_v_10_2_2((ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_20[9:0]),
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_11_nl));
  assign nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_11_nl = ({operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_8_nl
      , operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_9_nl})
      + 20'b00000000000000000001;
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_11_nl = nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_11_nl[19:0];
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_11_itm_19_6_1 = readslicef_20_14_6(operator_20_0_false_AC_TRN_AC_WRAP_acc_11_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_12_nl
      = conv_u2u_19_20(~ (in_data[258:240])) + 20'b00000000000000000001;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_12_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_12_nl[19:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_13_mx0
      = MUX_v_20_2_2(({1'b0 , (in_data[258:240])}), ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_12_nl,
      in_data[259]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_25_nl
      = MUX_v_9_8_2(9'b000000001, 9'b010011100, 9'b100011110, 9'b101111010, 9'b110110100,
      9'b111010110, 9'b111101001, 9'b111110100, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_12_itm_25_13[12:10]);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_29_mx0w1
      = conv_u2u_8_10(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_19[17:10])
      + ({1'b1 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_25_nl});
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_29_mx0w1
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_29_mx0w1[9:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_28_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_12_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_6_nl
      = ~(MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_29_mx0w1,
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_28_nl));
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_12_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_12_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_7_nl
      = ~(MUX_v_10_2_2((ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_19[9:0]),
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_12_nl));
  assign nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_12_nl = ({operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_6_nl
      , operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_7_nl})
      + 20'b00000000000000000001;
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_12_nl = nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_12_nl[19:0];
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_12_itm_19_6_1 = readslicef_20_14_6(operator_20_0_false_AC_TRN_AC_WRAP_acc_12_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_13_nl
      = conv_u2u_19_20(~ (in_data[278:260])) + 20'b00000000000000000001;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_13_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_13_nl[19:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_14_mx0
      = MUX_v_20_2_2(({1'b0 , (in_data[278:260])}), ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_13_nl,
      in_data[279]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_27_nl
      = MUX_v_9_8_2(9'b000000001, 9'b010011100, 9'b100011110, 9'b101111010, 9'b110110100,
      9'b111010110, 9'b111101001, 9'b111110100, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_13_itm_25_13[12:10]);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_30_mx0w1
      = conv_u2u_8_10(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_18[17:10])
      + ({1'b1 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_27_nl});
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_30_mx0w1
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_30_mx0w1[9:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_29_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_13_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_4_nl
      = ~(MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_30_mx0w1,
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_29_nl));
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_13_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_13_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_5_nl
      = ~(MUX_v_10_2_2((ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_18[9:0]),
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_13_nl));
  assign nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_13_nl = ({operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_4_nl
      , operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_5_nl})
      + 20'b00000000000000000001;
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_13_nl = nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_13_nl[19:0];
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_13_itm_19_6_1 = readslicef_20_14_6(operator_20_0_false_AC_TRN_AC_WRAP_acc_13_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_14_nl
      = conv_u2u_19_20(~ (in_data[298:280])) + 20'b00000000000000000001;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_14_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_14_nl[19:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_15_mx0
      = MUX_v_20_2_2(({1'b0 , (in_data[298:280])}), ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_14_nl,
      in_data[299]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_29_nl
      = MUX_v_9_8_2(9'b000000001, 9'b010011100, 9'b100011110, 9'b101111010, 9'b110110100,
      9'b111010110, 9'b111101001, 9'b111110100, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_14_itm_25_13[12:10]);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_31_mx0w1
      = conv_u2u_8_10(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_17[17:10])
      + ({1'b1 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_29_nl});
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_31_mx0w1
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_31_mx0w1[9:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_30_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_14_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_2_nl
      = ~(MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_31_mx0w1,
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_30_nl));
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_14_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_14_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_3_nl
      = ~(MUX_v_10_2_2((ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_17[9:0]),
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_14_nl));
  assign nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_14_nl = ({operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_2_nl
      , operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_3_nl})
      + 20'b00000000000000000001;
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_14_nl = nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_14_nl[19:0];
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_14_itm_19_6_1 = readslicef_20_14_6(operator_20_0_false_AC_TRN_AC_WRAP_acc_14_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_15_nl
      = conv_u2u_19_20(~ (in_data[318:300])) + 20'b00000000000000000001;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_15_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_15_nl[19:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_mx0
      = MUX_v_20_2_2(({1'b0 , (in_data[318:300])}), ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qelse_acc_15_nl,
      in_data[319]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_31_nl
      = MUX_v_9_8_2(9'b000000001, 9'b010011100, 9'b100011110, 9'b101111010, 9'b110110100,
      9'b111010110, 9'b111101001, 9'b111110100, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_15_itm_25_13[12:10]);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_16_mx0w1
      = conv_u2u_8_10(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_16[17:10])
      + ({1'b1 , ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_31_nl});
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_16_mx0w1
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_16_mx0w1[9:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_31_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_15_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_nl
      = ~(MUX_v_10_2_2(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_19_10_16_mx0w1,
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_31_nl));
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_15_nl
      = ~ ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_15_itm_5_1;
  assign operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_1_nl
      = ~(MUX_v_10_2_2((ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_16[9:0]),
      10'b1111111111, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_not_15_nl));
  assign nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_15_nl = ({operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_nl
      , operator_20_0_false_AC_TRN_AC_WRAP_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_nor_1_nl})
      + 20'b00000000000000000001;
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_15_nl = nl_operator_20_0_false_AC_TRN_AC_WRAP_acc_15_nl[19:0];
  assign operator_20_0_false_AC_TRN_AC_WRAP_acc_15_itm_19_6_1 = readslicef_20_14_6(operator_20_0_false_AC_TRN_AC_WRAP_acc_15_nl);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_30_nl
      = MUX_v_8_8_2(8'b10011011, 8'b10000010, 8'b01011100, 8'b00111010, 8'b00100010,
      8'b00010011, 8'b00001010, 8'b00000110, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_15_itm_25_13[12:10]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_16
      = conv_u2u_18_18(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_30_nl
      * (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_15_itm_25_13[9:0]));
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_15_nl
      = ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_mx0
      * 10'b1100110011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_15_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_15_nl[25:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_15_itm_25_13
      = readslicef_26_13_13(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_15_nl);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_28_nl
      = MUX_v_8_8_2(8'b10011011, 8'b10000010, 8'b01011100, 8'b00111010, 8'b00100010,
      8'b00010011, 8'b00001010, 8'b00000110, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_14_itm_25_13[12:10]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_17
      = conv_u2u_18_18(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_28_nl
      * (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_14_itm_25_13[9:0]));
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_14_nl
      = ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_15_mx0
      * 10'b1100110011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_14_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_14_nl[25:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_14_itm_25_13
      = readslicef_26_13_13(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_14_nl);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_26_nl
      = MUX_v_8_8_2(8'b10011011, 8'b10000010, 8'b01011100, 8'b00111010, 8'b00100010,
      8'b00010011, 8'b00001010, 8'b00000110, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_13_itm_25_13[12:10]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_18
      = conv_u2u_18_18(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_26_nl
      * (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_13_itm_25_13[9:0]));
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_13_nl
      = ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_14_mx0
      * 10'b1100110011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_13_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_13_nl[25:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_13_itm_25_13
      = readslicef_26_13_13(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_13_nl);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_24_nl
      = MUX_v_8_8_2(8'b10011011, 8'b10000010, 8'b01011100, 8'b00111010, 8'b00100010,
      8'b00010011, 8'b00001010, 8'b00000110, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_12_itm_25_13[12:10]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_19
      = conv_u2u_18_18(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_24_nl
      * (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_12_itm_25_13[9:0]));
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_12_nl
      = ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_13_mx0
      * 10'b1100110011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_12_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_12_nl[25:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_12_itm_25_13
      = readslicef_26_13_13(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_12_nl);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_22_nl
      = MUX_v_8_8_2(8'b10011011, 8'b10000010, 8'b01011100, 8'b00111010, 8'b00100010,
      8'b00010011, 8'b00001010, 8'b00000110, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_11_itm_25_13[12:10]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_20
      = conv_u2u_18_18(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_22_nl
      * (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_11_itm_25_13[9:0]));
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_11_nl
      = ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_12_mx0
      * 10'b1100110011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_11_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_11_nl[25:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_11_itm_25_13
      = readslicef_26_13_13(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_11_nl);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_20_nl
      = MUX_v_8_8_2(8'b10011011, 8'b10000010, 8'b01011100, 8'b00111010, 8'b00100010,
      8'b00010011, 8'b00001010, 8'b00000110, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_10_itm_25_13[12:10]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_21
      = conv_u2u_18_18(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_20_nl
      * (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_10_itm_25_13[9:0]));
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_10_nl
      = ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_11_mx0
      * 10'b1100110011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_10_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_10_nl[25:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_10_itm_25_13
      = readslicef_26_13_13(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_10_nl);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_18_nl
      = MUX_v_8_8_2(8'b10011011, 8'b10000010, 8'b01011100, 8'b00111010, 8'b00100010,
      8'b00010011, 8'b00001010, 8'b00000110, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_9_itm_25_13[12:10]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_22
      = conv_u2u_18_18(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_18_nl
      * (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_9_itm_25_13[9:0]));
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_9_nl
      = ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_10_mx0
      * 10'b1100110011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_9_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_9_nl[25:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_9_itm_25_13
      = readslicef_26_13_13(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_9_nl);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_16_nl
      = MUX_v_8_8_2(8'b10011011, 8'b10000010, 8'b01011100, 8'b00111010, 8'b00100010,
      8'b00010011, 8'b00001010, 8'b00000110, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_8_itm_25_13[12:10]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_23
      = conv_u2u_18_18(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_16_nl
      * (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_8_itm_25_13[9:0]));
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_8_nl
      = ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_9_mx0
      * 10'b1100110011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_8_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_8_nl[25:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_8_itm_25_13
      = readslicef_26_13_13(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_8_nl);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_14_nl
      = MUX_v_8_8_2(8'b10011011, 8'b10000010, 8'b01011100, 8'b00111010, 8'b00100010,
      8'b00010011, 8'b00001010, 8'b00000110, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_7_itm_25_13[12:10]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_24
      = conv_u2u_18_18(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_14_nl
      * (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_7_itm_25_13[9:0]));
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_7_nl
      = ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_8_mx0
      * 10'b1100110011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_7_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_7_nl[25:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_7_itm_25_13
      = readslicef_26_13_13(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_7_nl);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_12_nl
      = MUX_v_8_8_2(8'b10011011, 8'b10000010, 8'b01011100, 8'b00111010, 8'b00100010,
      8'b00010011, 8'b00001010, 8'b00000110, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_6_itm_25_13[12:10]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_25
      = conv_u2u_18_18(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_12_nl
      * (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_6_itm_25_13[9:0]));
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_6_nl
      = ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_7_mx0
      * 10'b1100110011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_6_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_6_nl[25:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_6_itm_25_13
      = readslicef_26_13_13(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_6_nl);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_10_nl
      = MUX_v_8_8_2(8'b10011011, 8'b10000010, 8'b01011100, 8'b00111010, 8'b00100010,
      8'b00010011, 8'b00001010, 8'b00000110, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_5_itm_25_13[12:10]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_26
      = conv_u2u_18_18(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_10_nl
      * (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_5_itm_25_13[9:0]));
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_5_nl
      = ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_6_mx0
      * 10'b1100110011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_5_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_5_nl[25:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_5_itm_25_13
      = readslicef_26_13_13(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_5_nl);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_8_nl
      = MUX_v_8_8_2(8'b10011011, 8'b10000010, 8'b01011100, 8'b00111010, 8'b00100010,
      8'b00010011, 8'b00001010, 8'b00000110, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_4_itm_25_13[12:10]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_27
      = conv_u2u_18_18(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_8_nl
      * (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_4_itm_25_13[9:0]));
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_4_nl
      = ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_5_mx0
      * 10'b1100110011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_4_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_4_nl[25:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_4_itm_25_13
      = readslicef_26_13_13(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_4_nl);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_6_nl
      = MUX_v_8_8_2(8'b10011011, 8'b10000010, 8'b01011100, 8'b00111010, 8'b00100010,
      8'b00010011, 8'b00001010, 8'b00000110, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_3_itm_25_13[12:10]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_28
      = conv_u2u_18_18(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_6_nl
      * (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_3_itm_25_13[9:0]));
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_3_nl
      = ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_4_mx0
      * 10'b1100110011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_3_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_3_nl[25:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_3_itm_25_13
      = readslicef_26_13_13(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_3_nl);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_4_nl
      = MUX_v_8_8_2(8'b10011011, 8'b10000010, 8'b01011100, 8'b00111010, 8'b00100010,
      8'b00010011, 8'b00001010, 8'b00000110, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_2_itm_25_13[12:10]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_29
      = conv_u2u_18_18(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_4_nl
      * (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_2_itm_25_13[9:0]));
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_2_nl
      = ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_3_mx0
      * 10'b1100110011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_2_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_2_nl[25:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_2_itm_25_13
      = readslicef_26_13_13(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_2_nl);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_2_nl
      = MUX_v_8_8_2(8'b10011011, 8'b10000010, 8'b01011100, 8'b00111010, 8'b00100010,
      8'b00010011, 8'b00001010, 8'b00000110, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_1_itm_25_13[12:10]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_30
      = conv_u2u_18_18(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_2_nl
      * (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_1_itm_25_13[9:0]));
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_1_nl
      = ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_2_mx0
      * 10'b1100110011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_1_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_1_nl[25:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_1_itm_25_13
      = readslicef_26_13_13(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_1_nl);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_nl
      = MUX_v_8_8_2(8'b10011011, 8'b10000010, 8'b01011100, 8'b00111010, 8'b00100010,
      8'b00010011, 8'b00001010, 8'b00000110, ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_itm_25_13[12:10]);
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mul_psp_31
      = conv_u2u_18_18(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_output_pwl_mux_nl
      * (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_itm_25_13[9:0]));
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_nl
      = ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_1_mx0
      * 10'b1100110011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_nl[25:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_itm_25_13
      = readslicef_26_13_13(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_x_in_sc_mul_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_15_nl
      = (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_mx0[19:14])
      + 6'b111011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_15_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_15_nl[5:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_15_itm_5_1
      = readslicef_6_1_5(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_15_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_14_nl
      = (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_15_mx0[19:14])
      + 6'b111011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_14_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_14_nl[5:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_14_itm_5_1
      = readslicef_6_1_5(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_14_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_13_nl
      = (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_14_mx0[19:14])
      + 6'b111011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_13_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_13_nl[5:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_13_itm_5_1
      = readslicef_6_1_5(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_13_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_12_nl
      = (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_13_mx0[19:14])
      + 6'b111011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_12_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_12_nl[5:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_12_itm_5_1
      = readslicef_6_1_5(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_12_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_11_nl
      = (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_12_mx0[19:14])
      + 6'b111011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_11_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_11_nl[5:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_11_itm_5_1
      = readslicef_6_1_5(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_11_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_10_nl
      = (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_11_mx0[19:14])
      + 6'b111011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_10_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_10_nl[5:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_10_itm_5_1
      = readslicef_6_1_5(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_10_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_9_nl
      = (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_10_mx0[19:14])
      + 6'b111011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_9_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_9_nl[5:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_9_itm_5_1
      = readslicef_6_1_5(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_9_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_8_nl
      = (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_9_mx0[19:14])
      + 6'b111011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_8_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_8_nl[5:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_8_itm_5_1
      = readslicef_6_1_5(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_8_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_7_nl
      = (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_8_mx0[19:14])
      + 6'b111011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_7_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_7_nl[5:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_7_itm_5_1
      = readslicef_6_1_5(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_7_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_6_nl
      = (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_7_mx0[19:14])
      + 6'b111011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_6_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_6_nl[5:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_6_itm_5_1
      = readslicef_6_1_5(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_6_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_5_nl
      = (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_6_mx0[19:14])
      + 6'b111011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_5_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_5_nl[5:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_5_itm_5_1
      = readslicef_6_1_5(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_5_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_4_nl
      = (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_5_mx0[19:14])
      + 6'b111011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_4_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_4_nl[5:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_4_itm_5_1
      = readslicef_6_1_5(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_4_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_3_nl
      = (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_4_mx0[19:14])
      + 6'b111011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_3_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_3_nl[5:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_3_itm_5_1
      = readslicef_6_1_5(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_3_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_2_nl
      = (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_3_mx0[19:14])
      + 6'b111011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_2_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_2_nl[5:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_2_itm_5_1
      = readslicef_6_1_5(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_2_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_1_nl
      = (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_2_mx0[19:14])
      + 6'b111011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_1_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_1_nl[5:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_1_itm_5_1
      = readslicef_6_1_5(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_1_nl);
  assign nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_nl
      = (ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_1_qr_1_mx0[19:14])
      + 6'b111011;
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_nl
      = nl_ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_nl[5:0];
  assign ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_itm_5_1
      = readslicef_6_1_5(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_nl);
  assign and_dcpl = ~((in_data[19]) | ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_itm_5_1);
  assign and_dcpl_1 = (~ (in_data[19])) & ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_itm_5_1;
  assign and_dcpl_2 = ~((in_data[39]) | ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_1_itm_5_1);
  assign and_dcpl_3 = (~ (in_data[39])) & ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_1_itm_5_1;
  assign and_dcpl_4 = ~(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_2_itm_5_1
      | (in_data[59]));
  assign and_dcpl_5 = ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_2_itm_5_1
      & (~ (in_data[59]));
  assign and_dcpl_6 = ~(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_3_itm_5_1
      | (in_data[79]));
  assign and_dcpl_7 = ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_3_itm_5_1
      & (~ (in_data[79]));
  assign and_dcpl_8 = ~(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_4_itm_5_1
      | (in_data[99]));
  assign and_dcpl_9 = ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_4_itm_5_1
      & (~ (in_data[99]));
  assign and_dcpl_10 = ~(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_5_itm_5_1
      | (in_data[119]));
  assign and_dcpl_11 = ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_5_itm_5_1
      & (~ (in_data[119]));
  assign and_dcpl_12 = ~(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_6_itm_5_1
      | (in_data[139]));
  assign and_dcpl_13 = ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_6_itm_5_1
      & (~ (in_data[139]));
  assign and_dcpl_14 = ~(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_7_itm_5_1
      | (in_data[159]));
  assign and_dcpl_15 = ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_7_itm_5_1
      & (~ (in_data[159]));
  assign and_dcpl_16 = ~(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_8_itm_5_1
      | (in_data[179]));
  assign and_dcpl_17 = ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_8_itm_5_1
      & (~ (in_data[179]));
  assign and_dcpl_18 = ~(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_9_itm_5_1
      | (in_data[199]));
  assign and_dcpl_19 = ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_9_itm_5_1
      & (~ (in_data[199]));
  assign and_dcpl_20 = ~(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_10_itm_5_1
      | (in_data[219]));
  assign and_dcpl_21 = ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_10_itm_5_1
      & (~ (in_data[219]));
  assign and_dcpl_22 = ~(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_11_itm_5_1
      | (in_data[239]));
  assign and_dcpl_23 = ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_11_itm_5_1
      & (~ (in_data[239]));
  assign and_dcpl_24 = ~(ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_12_itm_5_1
      | (in_data[259]));
  assign and_dcpl_25 = ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_12_itm_5_1
      & (~ (in_data[259]));
  assign and_dcpl_26 = ~((in_data[279]) | ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_13_itm_5_1);
  assign and_dcpl_27 = (~ (in_data[279])) & ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_13_itm_5_1;
  assign and_dcpl_28 = ~((in_data[299]) | ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_14_itm_5_1);
  assign and_dcpl_29 = (~ (in_data[299])) & ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_14_itm_5_1;
  assign and_dcpl_30 = ~((in_data[319]) | ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_15_itm_5_1);
  assign and_dcpl_31 = (~ (in_data[319])) & ac_math_ac_sigmoid_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_AC_TRN_AC_WRAP_if_2_acc_15_itm_5_1;

  function automatic [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function automatic [19:0] MUX_v_20_2_2;
    input [19:0] input_0;
    input [19:0] input_1;
    input [0:0] sel;
    reg [19:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_20_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_8_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [2:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_8_8_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_8_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [8:0] input_2;
    input [8:0] input_3;
    input [8:0] input_4;
    input [8:0] input_5;
    input [8:0] input_6;
    input [8:0] input_7;
    input [2:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_9_8_2 = result;
  end
  endfunction


  function automatic [13:0] readslicef_20_14_6;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_20_14_6 = tmp[13:0];
  end
  endfunction


  function automatic [12:0] readslicef_26_13_13;
    input [25:0] vector;
    reg [25:0] tmp;
  begin
    tmp = vector >> 13;
    readslicef_26_13_13 = tmp[12:0];
  end
  endfunction


  function automatic [0:0] readslicef_6_1_5;
    input [5:0] vector;
    reg [5:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_6_1_5 = tmp[0:0];
  end
  endfunction


  function automatic [9:0] conv_u2u_8_10 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_10 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [17:0] conv_u2u_18_18 ;
    input [17:0]  vector ;
  begin
    conv_u2u_18_18 = vector;
  end
  endfunction


  function automatic [19:0] conv_u2u_19_20 ;
    input [18:0]  vector ;
  begin
    conv_u2u_19_20 = {1'b0, vector};
  end
  endfunction

endmodule




//------> ./ActUnit_Tanh.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   huaixil@sat8
//  Generated date: Fri Apr  8 23:10:59 2022
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Tanh
// ------------------------------------------------------------------


module ActUnit_Tanh (
  in_data, out_data
);
  input [319:0] in_data;
  output [319:0] out_data;


  // Interconnect Declarations
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_1_mx0;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_2_mx0;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_3_mx0;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_4_mx0;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_5_mx0;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_6_mx0;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_7_mx0;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_8_mx0;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_9_mx0;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_10_mx0;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_11_mx0;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_12_mx0;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_13_mx0;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_14_mx0;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_15_mx0;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_mx0;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_16;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_17;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_18;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_19;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_20;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_21;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_22;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_23;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_24;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_25;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_26;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_27;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_28;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_29;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_30;
  wire [17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_31;
  wire [10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_1_mx0w2_20_10;
  wire [11:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_1_mx0w2_20_10;
  wire [10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_2_mx0w2_20_10;
  wire [11:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_2_mx0w2_20_10;
  wire [10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_3_mx0w2_20_10;
  wire [11:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_3_mx0w2_20_10;
  wire [10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_4_mx0w2_20_10;
  wire [11:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_4_mx0w2_20_10;
  wire [10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_5_mx0w2_20_10;
  wire [11:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_5_mx0w2_20_10;
  wire [10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_6_mx0w2_20_10;
  wire [11:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_6_mx0w2_20_10;
  wire [10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_7_mx0w2_20_10;
  wire [11:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_7_mx0w2_20_10;
  wire [10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_8_mx0w2_20_10;
  wire [11:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_8_mx0w2_20_10;
  wire [10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_9_mx0w2_20_10;
  wire [11:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_9_mx0w2_20_10;
  wire [10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_10_mx0w2_20_10;
  wire [11:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_10_mx0w2_20_10;
  wire [10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_11_mx0w2_20_10;
  wire [11:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_11_mx0w2_20_10;
  wire [10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_12_mx0w2_20_10;
  wire [11:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_12_mx0w2_20_10;
  wire [10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_13_mx0w2_20_10;
  wire [11:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_13_mx0w2_20_10;
  wire [10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_14_mx0w2_20_10;
  wire [11:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_14_mx0w2_20_10;
  wire [10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_15_mx0w2_20_10;
  wire [11:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_15_mx0w2_20_10;
  wire [10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mx0w2_20_10;
  wire [11:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mx0w2_20_10;
  wire operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_15_itm_5_1;
  wire operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_14_itm_5_1;
  wire operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_13_itm_5_1;
  wire operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_12_itm_5_1;
  wire operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_11_itm_5_1;
  wire operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_10_itm_5_1;
  wire operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_9_itm_5_1;
  wire operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_8_itm_5_1;
  wire operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_7_itm_5_1;
  wire operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_6_itm_5_1;
  wire operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_5_itm_5_1;
  wire operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_4_itm_5_1;
  wire operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_3_itm_5_1;
  wire operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_2_itm_5_1;
  wire operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_1_itm_5_1;
  wire operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_itm_5_1;

  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_15_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TR000000;
  wire[15:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TR000000;
  wire[10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_32_nl;
  wire[3:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_32_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_nl;
  wire[0:0] nor_nl;
  wire[0:0] and_31_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_14_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_15_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000;
  wire[15:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_15_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000;
  wire[10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_30_nl;
  wire[3:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_7_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_38_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_1_nl;
  wire[0:0] nor_1_nl;
  wire[0:0] and_29_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_13_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_14_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000;
  wire[15:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_14_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000;
  wire[10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_28_nl;
  wire[3:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_14_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_44_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_2_nl;
  wire[0:0] nor_2_nl;
  wire[0:0] and_27_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_12_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_13_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000;
  wire[15:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_13_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000;
  wire[10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_26_nl;
  wire[3:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_21_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_50_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_3_nl;
  wire[0:0] nor_3_nl;
  wire[0:0] and_25_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_11_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_12_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000;
  wire[15:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_12_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000;
  wire[10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_24_nl;
  wire[3:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_28_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_56_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_4_nl;
  wire[0:0] nor_4_nl;
  wire[0:0] and_23_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_10_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_11_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000;
  wire[15:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_11_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000;
  wire[10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_22_nl;
  wire[3:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_35_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_62_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_5_nl;
  wire[0:0] nor_5_nl;
  wire[0:0] and_21_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_9_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_10_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000;
  wire[15:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_10_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000;
  wire[10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_20_nl;
  wire[3:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_42_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_68_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_6_nl;
  wire[0:0] nor_6_nl;
  wire[0:0] and_19_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_8_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_9_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000;
  wire[15:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_9_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000;
  wire[10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_18_nl;
  wire[3:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_49_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_74_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_7_nl;
  wire[0:0] nor_7_nl;
  wire[0:0] and_17_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_7_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_8_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000;
  wire[15:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_8_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000;
  wire[10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_16_nl;
  wire[3:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_56_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_80_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_8_nl;
  wire[0:0] nor_8_nl;
  wire[0:0] and_15_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_6_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_7_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000;
  wire[15:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_7_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000;
  wire[10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_14_nl;
  wire[3:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_63_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_86_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_9_nl;
  wire[0:0] nor_9_nl;
  wire[0:0] and_13_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_5_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_6_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000;
  wire[15:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_6_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000;
  wire[10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_12_nl;
  wire[3:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_70_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_92_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_10_nl;
  wire[0:0] nor_10_nl;
  wire[0:0] and_11_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_4_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_5_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000;
  wire[15:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_5_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000;
  wire[10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_10_nl;
  wire[3:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_77_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_98_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_11_nl;
  wire[0:0] nor_11_nl;
  wire[0:0] and_9_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_3_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_4_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000;
  wire[15:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_4_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000;
  wire[10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_8_nl;
  wire[3:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_84_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_104_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_12_nl;
  wire[0:0] nor_12_nl;
  wire[0:0] and_7_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_2_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_3_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000;
  wire[15:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_3_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000;
  wire[10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_6_nl;
  wire[3:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_91_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_110_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_13_nl;
  wire[0:0] nor_13_nl;
  wire[0:0] and_5_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_1_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_2_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000;
  wire[15:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_2_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000;
  wire[10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_4_nl;
  wire[3:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_98_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_116_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_14_nl;
  wire[0:0] nor_14_nl;
  wire[0:0] and_3_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_nl;
  wire[14:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_1_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000;
  wire[15:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_1_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000;
  wire[10:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_nl;
  wire[3:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_105_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_122_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_15_nl;
  wire[0:0] nor_15_nl;
  wire[0:0] and_1_nl;
  wire[17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_nl;
  wire[18:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_nl;
  wire[9:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_1_nl;
  wire[17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_1_nl;
  wire[18:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_1_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_1_nl;
  wire[9:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_3_nl;
  wire[17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_2_nl;
  wire[18:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_2_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_2_nl;
  wire[9:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_5_nl;
  wire[17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_3_nl;
  wire[18:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_3_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_3_nl;
  wire[9:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_7_nl;
  wire[17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_4_nl;
  wire[18:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_4_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_4_nl;
  wire[9:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_9_nl;
  wire[17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_5_nl;
  wire[18:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_5_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_5_nl;
  wire[9:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_11_nl;
  wire[17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_6_nl;
  wire[18:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_6_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_6_nl;
  wire[9:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_13_nl;
  wire[17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_7_nl;
  wire[18:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_7_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_7_nl;
  wire[9:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_15_nl;
  wire[17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_8_nl;
  wire[18:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_8_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_8_nl;
  wire[9:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_17_nl;
  wire[17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_9_nl;
  wire[18:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_9_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_9_nl;
  wire[9:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_19_nl;
  wire[17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_10_nl;
  wire[18:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_10_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_10_nl;
  wire[9:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_21_nl;
  wire[17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_11_nl;
  wire[18:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_11_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_11_nl;
  wire[9:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_23_nl;
  wire[17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_12_nl;
  wire[18:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_12_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_12_nl;
  wire[9:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_25_nl;
  wire[17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_13_nl;
  wire[18:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_13_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_13_nl;
  wire[9:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_27_nl;
  wire[17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_14_nl;
  wire[18:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_14_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_14_nl;
  wire[9:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_29_nl;
  wire[17:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_15_nl;
  wire[18:0] nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_15_nl;
  wire[0:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_15_nl;
  wire[9:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_31_nl;
  wire[7:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_33_nl;
  wire[7:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_34_nl;
  wire[7:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_35_nl;
  wire[7:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_36_nl;
  wire[7:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_37_nl;
  wire[7:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_38_nl;
  wire[7:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_39_nl;
  wire[7:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_40_nl;
  wire[7:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_41_nl;
  wire[7:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_42_nl;
  wire[7:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_43_nl;
  wire[7:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_44_nl;
  wire[7:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_45_nl;
  wire[7:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_46_nl;
  wire[7:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_2_nl;
  wire[7:0] ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_47_nl;
  wire[5:0] operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_15_nl;
  wire[6:0] nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_15_nl;
  wire[5:0] operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_14_nl;
  wire[6:0] nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_14_nl;
  wire[5:0] operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_13_nl;
  wire[6:0] nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_13_nl;
  wire[5:0] operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_12_nl;
  wire[6:0] nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_12_nl;
  wire[5:0] operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_11_nl;
  wire[6:0] nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_11_nl;
  wire[5:0] operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_10_nl;
  wire[6:0] nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_10_nl;
  wire[5:0] operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_9_nl;
  wire[6:0] nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_9_nl;
  wire[5:0] operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_8_nl;
  wire[6:0] nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_8_nl;
  wire[5:0] operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_7_nl;
  wire[6:0] nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_7_nl;
  wire[5:0] operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_6_nl;
  wire[6:0] nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_6_nl;
  wire[5:0] operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_5_nl;
  wire[6:0] nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_5_nl;
  wire[5:0] operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_4_nl;
  wire[6:0] nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_4_nl;
  wire[5:0] operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_3_nl;
  wire[6:0] nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_3_nl;
  wire[5:0] operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_2_nl;
  wire[6:0] nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_2_nl;
  wire[5:0] operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_1_nl;
  wire[6:0] nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_1_nl;
  wire[5:0] operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_nl;
  wire[6:0] nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_nl;

  // Interconnect Declarations for Component Instantiations
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_32_nl
      = MUX_v_11_2_2(11'b01111111111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mx0w2_20_10,
      operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_15_itm_5_1);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_32_nl
      = ~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_15_itm_5_1;
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_nl
      = ~(MUX_v_4_2_2((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_16[9:6]),
      4'b1111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_32_nl));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_nl
      = (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_16[0])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_15_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_16[1])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_15_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_16[2])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_15_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_16[3])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_15_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_16[4])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_15_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_16[5])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_15_itm_5_1)));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TR000000
      = ({(~ ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_32_nl)
      , ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_nl})
      + conv_u2s_1_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TR000000
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TR000000[14:0];
  assign nor_nl = ~((in_data[319]) | operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_15_itm_5_1);
  assign and_31_nl = (~ (in_data[319])) & operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_15_itm_5_1;
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_15_nl
      = MUX1HOT_v_15_3_2(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TR000000,
      15'b011111111111111, ({ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mx0w2_20_10
      , (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_16[9:6])}),
      {(in_data[319]) , nor_nl , and_31_nl});
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_30_nl
      = MUX_v_11_2_2(11'b01111111111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_15_mx0w2_20_10,
      operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_14_itm_5_1);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_38_nl
      = ~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_14_itm_5_1;
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_7_nl
      = ~(MUX_v_4_2_2((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_17[9:6]),
      4'b1111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_38_nl));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_1_nl
      = (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_17[0])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_14_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_17[1])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_14_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_17[2])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_14_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_17[3])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_14_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_17[4])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_14_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_17[5])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_14_itm_5_1)));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_15_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000
      = ({(~ ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_30_nl)
      , ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_7_nl})
      + conv_u2s_1_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_1_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_15_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_15_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000[14:0];
  assign nor_1_nl = ~((in_data[299]) | operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_14_itm_5_1);
  assign and_29_nl = (~ (in_data[299])) & operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_14_itm_5_1;
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_14_nl
      = MUX1HOT_v_15_3_2(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_15_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000,
      15'b011111111111111, ({ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_15_mx0w2_20_10
      , (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_17[9:6])}),
      {(in_data[299]) , nor_1_nl , and_29_nl});
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_28_nl
      = MUX_v_11_2_2(11'b01111111111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_14_mx0w2_20_10,
      operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_13_itm_5_1);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_44_nl
      = ~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_13_itm_5_1;
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_14_nl
      = ~(MUX_v_4_2_2((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_18[9:6]),
      4'b1111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_44_nl));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_2_nl
      = (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_18[0])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_13_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_18[1])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_13_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_18[2])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_13_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_18[3])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_13_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_18[4])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_13_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_18[5])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_13_itm_5_1)));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_14_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000
      = ({(~ ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_28_nl)
      , ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_14_nl})
      + conv_u2s_1_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_2_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_14_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_14_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000[14:0];
  assign nor_2_nl = ~((in_data[279]) | operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_13_itm_5_1);
  assign and_27_nl = (~ (in_data[279])) & operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_13_itm_5_1;
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_13_nl
      = MUX1HOT_v_15_3_2(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_14_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000,
      15'b011111111111111, ({ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_14_mx0w2_20_10
      , (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_18[9:6])}),
      {(in_data[279]) , nor_2_nl , and_27_nl});
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_26_nl
      = MUX_v_11_2_2(11'b01111111111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_13_mx0w2_20_10,
      operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_12_itm_5_1);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_50_nl
      = ~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_12_itm_5_1;
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_21_nl
      = ~(MUX_v_4_2_2((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_19[9:6]),
      4'b1111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_50_nl));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_3_nl
      = (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_19[0])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_12_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_19[1])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_12_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_19[2])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_12_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_19[3])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_12_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_19[4])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_12_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_19[5])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_12_itm_5_1)));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_13_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000
      = ({(~ ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_26_nl)
      , ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_21_nl})
      + conv_u2s_1_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_3_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_13_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_13_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000[14:0];
  assign nor_3_nl = ~(operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_12_itm_5_1 |
      (in_data[259]));
  assign and_25_nl = operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_12_itm_5_1 &
      (~ (in_data[259]));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_12_nl
      = MUX1HOT_v_15_3_2(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_13_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000,
      15'b011111111111111, ({ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_13_mx0w2_20_10
      , (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_19[9:6])}),
      {(in_data[259]) , nor_3_nl , and_25_nl});
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_24_nl
      = MUX_v_11_2_2(11'b01111111111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_12_mx0w2_20_10,
      operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_11_itm_5_1);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_56_nl
      = ~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_11_itm_5_1;
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_28_nl
      = ~(MUX_v_4_2_2((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_20[9:6]),
      4'b1111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_56_nl));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_4_nl
      = (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_20[0])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_11_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_20[1])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_11_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_20[2])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_11_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_20[3])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_11_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_20[4])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_11_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_20[5])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_11_itm_5_1)));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_12_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000
      = ({(~ ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_24_nl)
      , ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_28_nl})
      + conv_u2s_1_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_4_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_12_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_12_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000[14:0];
  assign nor_4_nl = ~(operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_11_itm_5_1 |
      (in_data[239]));
  assign and_23_nl = operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_11_itm_5_1 &
      (~ (in_data[239]));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_11_nl
      = MUX1HOT_v_15_3_2(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_12_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000,
      15'b011111111111111, ({ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_12_mx0w2_20_10
      , (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_20[9:6])}),
      {(in_data[239]) , nor_4_nl , and_23_nl});
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_22_nl
      = MUX_v_11_2_2(11'b01111111111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_11_mx0w2_20_10,
      operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_10_itm_5_1);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_62_nl
      = ~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_10_itm_5_1;
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_35_nl
      = ~(MUX_v_4_2_2((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_21[9:6]),
      4'b1111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_62_nl));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_5_nl
      = (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_21[0])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_10_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_21[1])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_10_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_21[2])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_10_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_21[3])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_10_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_21[4])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_10_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_21[5])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_10_itm_5_1)));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_11_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000
      = ({(~ ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_22_nl)
      , ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_35_nl})
      + conv_u2s_1_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_5_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_11_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_11_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000[14:0];
  assign nor_5_nl = ~(operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_10_itm_5_1 |
      (in_data[219]));
  assign and_21_nl = operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_10_itm_5_1 &
      (~ (in_data[219]));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_10_nl
      = MUX1HOT_v_15_3_2(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_11_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000,
      15'b011111111111111, ({ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_11_mx0w2_20_10
      , (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_21[9:6])}),
      {(in_data[219]) , nor_5_nl , and_21_nl});
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_20_nl
      = MUX_v_11_2_2(11'b01111111111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_10_mx0w2_20_10,
      operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_9_itm_5_1);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_68_nl
      = ~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_9_itm_5_1;
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_42_nl
      = ~(MUX_v_4_2_2((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_22[9:6]),
      4'b1111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_68_nl));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_6_nl
      = (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_22[0])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_9_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_22[1])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_9_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_22[2])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_9_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_22[3])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_9_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_22[4])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_9_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_22[5])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_9_itm_5_1)));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_10_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000
      = ({(~ ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_20_nl)
      , ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_42_nl})
      + conv_u2s_1_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_6_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_10_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_10_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000[14:0];
  assign nor_6_nl = ~(operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_9_itm_5_1 |
      (in_data[199]));
  assign and_19_nl = operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_9_itm_5_1 & (~
      (in_data[199]));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_9_nl
      = MUX1HOT_v_15_3_2(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_10_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC000000,
      15'b011111111111111, ({ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_10_mx0w2_20_10
      , (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_22[9:6])}),
      {(in_data[199]) , nor_6_nl , and_19_nl});
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_18_nl
      = MUX_v_11_2_2(11'b01111111111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_9_mx0w2_20_10,
      operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_8_itm_5_1);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_74_nl
      = ~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_8_itm_5_1;
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_49_nl
      = ~(MUX_v_4_2_2((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_23[9:6]),
      4'b1111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_74_nl));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_7_nl
      = (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_23[0])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_8_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_23[1])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_8_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_23[2])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_8_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_23[3])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_8_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_23[4])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_8_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_23[5])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_8_itm_5_1)));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_9_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000
      = ({(~ ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_18_nl)
      , ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_49_nl})
      + conv_u2s_1_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_7_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_9_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_9_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000[14:0];
  assign nor_7_nl = ~(operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_8_itm_5_1 |
      (in_data[179]));
  assign and_17_nl = operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_8_itm_5_1 & (~
      (in_data[179]));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_8_nl
      = MUX1HOT_v_15_3_2(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_9_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000,
      15'b011111111111111, ({ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_9_mx0w2_20_10
      , (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_23[9:6])}),
      {(in_data[179]) , nor_7_nl , and_17_nl});
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_16_nl
      = MUX_v_11_2_2(11'b01111111111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_8_mx0w2_20_10,
      operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_7_itm_5_1);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_80_nl
      = ~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_7_itm_5_1;
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_56_nl
      = ~(MUX_v_4_2_2((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_24[9:6]),
      4'b1111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_80_nl));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_8_nl
      = (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_24[0])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_7_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_24[1])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_7_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_24[2])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_7_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_24[3])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_7_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_24[4])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_7_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_24[5])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_7_itm_5_1)));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_8_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000
      = ({(~ ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_16_nl)
      , ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_56_nl})
      + conv_u2s_1_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_8_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_8_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_8_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000[14:0];
  assign nor_8_nl = ~(operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_7_itm_5_1 |
      (in_data[159]));
  assign and_15_nl = operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_7_itm_5_1 & (~
      (in_data[159]));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_7_nl
      = MUX1HOT_v_15_3_2(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_8_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000,
      15'b011111111111111, ({ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_8_mx0w2_20_10
      , (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_24[9:6])}),
      {(in_data[159]) , nor_8_nl , and_15_nl});
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_14_nl
      = MUX_v_11_2_2(11'b01111111111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_7_mx0w2_20_10,
      operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_6_itm_5_1);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_86_nl
      = ~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_6_itm_5_1;
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_63_nl
      = ~(MUX_v_4_2_2((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_25[9:6]),
      4'b1111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_86_nl));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_9_nl
      = (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_25[0])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_6_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_25[1])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_6_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_25[2])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_6_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_25[3])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_6_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_25[4])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_6_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_25[5])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_6_itm_5_1)));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_7_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000
      = ({(~ ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_14_nl)
      , ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_63_nl})
      + conv_u2s_1_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_9_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_7_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_7_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000[14:0];
  assign nor_9_nl = ~(operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_6_itm_5_1 |
      (in_data[139]));
  assign and_13_nl = operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_6_itm_5_1 & (~
      (in_data[139]));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_6_nl
      = MUX1HOT_v_15_3_2(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_7_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000,
      15'b011111111111111, ({ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_7_mx0w2_20_10
      , (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_25[9:6])}),
      {(in_data[139]) , nor_9_nl , and_13_nl});
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_12_nl
      = MUX_v_11_2_2(11'b01111111111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_6_mx0w2_20_10,
      operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_5_itm_5_1);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_92_nl
      = ~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_5_itm_5_1;
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_70_nl
      = ~(MUX_v_4_2_2((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_26[9:6]),
      4'b1111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_92_nl));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_10_nl
      = (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_26[0])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_5_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_26[1])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_5_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_26[2])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_5_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_26[3])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_5_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_26[4])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_5_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_26[5])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_5_itm_5_1)));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_6_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000
      = ({(~ ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_12_nl)
      , ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_70_nl})
      + conv_u2s_1_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_10_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_6_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_6_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000[14:0];
  assign nor_10_nl = ~(operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_5_itm_5_1 |
      (in_data[119]));
  assign and_11_nl = operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_5_itm_5_1 & (~
      (in_data[119]));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_5_nl
      = MUX1HOT_v_15_3_2(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_6_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000,
      15'b011111111111111, ({ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_6_mx0w2_20_10
      , (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_26[9:6])}),
      {(in_data[119]) , nor_10_nl , and_11_nl});
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_10_nl
      = MUX_v_11_2_2(11'b01111111111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_5_mx0w2_20_10,
      operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_4_itm_5_1);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_98_nl
      = ~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_4_itm_5_1;
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_77_nl
      = ~(MUX_v_4_2_2((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_27[9:6]),
      4'b1111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_98_nl));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_11_nl
      = (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_27[0])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_4_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_27[1])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_4_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_27[2])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_4_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_27[3])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_4_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_27[4])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_4_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_27[5])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_4_itm_5_1)));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_5_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000
      = ({(~ ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_10_nl)
      , ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_77_nl})
      + conv_u2s_1_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_11_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_5_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_5_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000[14:0];
  assign nor_11_nl = ~(operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_4_itm_5_1 |
      (in_data[99]));
  assign and_9_nl = operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_4_itm_5_1 & (~
      (in_data[99]));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_4_nl
      = MUX1HOT_v_15_3_2(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_5_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000,
      15'b011111111111111, ({ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_5_mx0w2_20_10
      , (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_27[9:6])}),
      {(in_data[99]) , nor_11_nl , and_9_nl});
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_8_nl
      = MUX_v_11_2_2(11'b01111111111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_4_mx0w2_20_10,
      operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_3_itm_5_1);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_104_nl
      = ~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_3_itm_5_1;
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_84_nl
      = ~(MUX_v_4_2_2((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_28[9:6]),
      4'b1111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_104_nl));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_12_nl
      = (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_28[0])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_3_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_28[1])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_3_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_28[2])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_3_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_28[3])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_3_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_28[4])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_3_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_28[5])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_3_itm_5_1)));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_4_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000
      = ({(~ ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_8_nl)
      , ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_84_nl})
      + conv_u2s_1_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_12_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_4_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_4_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000[14:0];
  assign nor_12_nl = ~(operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_3_itm_5_1 |
      (in_data[79]));
  assign and_7_nl = operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_3_itm_5_1 & (~
      (in_data[79]));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_3_nl
      = MUX1HOT_v_15_3_2(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_4_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000,
      15'b011111111111111, ({ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_4_mx0w2_20_10
      , (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_28[9:6])}),
      {(in_data[79]) , nor_12_nl , and_7_nl});
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_6_nl
      = MUX_v_11_2_2(11'b01111111111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_3_mx0w2_20_10,
      operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_2_itm_5_1);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_110_nl
      = ~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_2_itm_5_1;
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_91_nl
      = ~(MUX_v_4_2_2((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_29[9:6]),
      4'b1111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_110_nl));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_13_nl
      = (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_29[0])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_2_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_29[1])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_2_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_29[2])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_2_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_29[3])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_2_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_29[4])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_2_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_29[5])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_2_itm_5_1)));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_3_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000
      = ({(~ ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_6_nl)
      , ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_91_nl})
      + conv_u2s_1_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_13_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_3_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_3_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000[14:0];
  assign nor_13_nl = ~(operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_2_itm_5_1 |
      (in_data[59]));
  assign and_5_nl = operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_2_itm_5_1 & (~
      (in_data[59]));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_2_nl
      = MUX1HOT_v_15_3_2(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_3_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000,
      15'b011111111111111, ({ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_3_mx0w2_20_10
      , (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_29[9:6])}),
      {(in_data[59]) , nor_13_nl , and_5_nl});
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_4_nl
      = MUX_v_11_2_2(11'b01111111111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_2_mx0w2_20_10,
      operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_1_itm_5_1);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_116_nl
      = ~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_1_itm_5_1;
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_98_nl
      = ~(MUX_v_4_2_2((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_30[9:6]),
      4'b1111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_116_nl));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_14_nl
      = (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_30[0])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_1_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_30[1])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_1_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_30[2])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_1_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_30[3])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_1_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_30[4])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_1_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_30[5])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_1_itm_5_1)));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_2_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000
      = ({(~ ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_4_nl)
      , ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_98_nl})
      + conv_u2s_1_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_14_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_2_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_2_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000[14:0];
  assign nor_14_nl = ~((in_data[39]) | operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_1_itm_5_1);
  assign and_3_nl = (~ (in_data[39])) & operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_1_itm_5_1;
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_1_nl
      = MUX1HOT_v_15_3_2(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_2_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000,
      15'b011111111111111, ({ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_2_mx0w2_20_10
      , (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_30[9:6])}),
      {(in_data[39]) , nor_14_nl , and_3_nl});
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_nl
      = MUX_v_11_2_2(11'b01111111111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_1_mx0w2_20_10,
      operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_itm_5_1);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_122_nl
      = ~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_itm_5_1;
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_105_nl
      = ~(MUX_v_4_2_2((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_31[9:6]),
      4'b1111, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_not_122_nl));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_15_nl
      = (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_31[0])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_31[1])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_31[2])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_31[3])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_31[4])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_itm_5_1))) & (~((ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_31[5])
      | (~ operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_itm_5_1)));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_1_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000
      = ({(~ ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_nl)
      , ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_nor_105_nl})
      + conv_u2s_1_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_and_15_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_1_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_1_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000[14:0];
  assign nor_15_nl = ~((in_data[19]) | operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_itm_5_1);
  assign and_1_nl = (~ (in_data[19])) & operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_itm_5_1;
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_nl
      = MUX1HOT_v_15_3_2(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_1_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_000000,
      15'b011111111111111, ({ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_1_mx0w2_20_10
      , (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_31[9:6])}),
      {(in_data[19]) , nor_15_nl , and_1_nl});
  assign out_data = signext_320_315({ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_15_nl
      , (signext_20_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_14_nl))
      , (signext_20_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_13_nl))
      , (signext_20_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_12_nl))
      , (signext_20_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_11_nl))
      , (signext_20_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_10_nl))
      , (signext_20_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_9_nl))
      , (signext_20_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_8_nl))
      , (signext_20_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_7_nl))
      , (signext_20_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_6_nl))
      , (signext_20_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_5_nl))
      , (signext_20_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_4_nl))
      , (signext_20_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_3_nl))
      , (signext_20_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_2_nl))
      , (signext_20_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_1_nl))
      , (signext_20_15(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux1h_nl))});
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_nl
      = ~((in_data[1:0]!=2'b00));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_nl
      = conv_u2u_17_18(~ (in_data[18:2])) + conv_u2u_1_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_nl
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_nl[17:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_1_mx0
      = MUX_v_18_2_2(({1'b0 , (in_data[18:2])}), ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_nl,
      in_data[19]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_1_nl
      = MUX_v_10_12_2(10'b0000000001, 10'b0011111100, 10'b0111011100, 10'b1010001101,
      10'b1100001111, 10'b1101100111, 10'b1110100000, 10'b1111000101, 10'b1111011100,
      10'b1111101010, 10'b1111110011, 10'b1111111000, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_1_mx0[13:10]);
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_1_mx0w2_20_10
      = conv_u2u_8_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_31[17:10])
      + conv_u2u_10_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_1_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_1_mx0w2_20_10
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_1_mx0w2_20_10[10:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_1_nl
      = ~((in_data[21:20]!=2'b00));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_1_nl
      = conv_u2u_17_18(~ (in_data[38:22])) + conv_u2u_1_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_1_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_1_nl
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_1_nl[17:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_2_mx0
      = MUX_v_18_2_2(({1'b0 , (in_data[38:22])}), ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_1_nl,
      in_data[39]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_3_nl
      = MUX_v_10_12_2(10'b0000000001, 10'b0011111100, 10'b0111011100, 10'b1010001101,
      10'b1100001111, 10'b1101100111, 10'b1110100000, 10'b1111000101, 10'b1111011100,
      10'b1111101010, 10'b1111110011, 10'b1111111000, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_2_mx0[13:10]);
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_2_mx0w2_20_10
      = conv_u2u_8_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_30[17:10])
      + conv_u2u_10_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_3_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_2_mx0w2_20_10
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_2_mx0w2_20_10[10:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_2_nl
      = ~((in_data[41:40]!=2'b00));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_2_nl
      = conv_u2u_17_18(~ (in_data[58:42])) + conv_u2u_1_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_2_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_2_nl
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_2_nl[17:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_3_mx0
      = MUX_v_18_2_2(({1'b0 , (in_data[58:42])}), ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_2_nl,
      in_data[59]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_5_nl
      = MUX_v_10_12_2(10'b0000000001, 10'b0011111100, 10'b0111011100, 10'b1010001101,
      10'b1100001111, 10'b1101100111, 10'b1110100000, 10'b1111000101, 10'b1111011100,
      10'b1111101010, 10'b1111110011, 10'b1111111000, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_3_mx0[13:10]);
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_3_mx0w2_20_10
      = conv_u2u_8_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_29[17:10])
      + conv_u2u_10_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_5_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_3_mx0w2_20_10
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_3_mx0w2_20_10[10:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_3_nl
      = ~((in_data[61:60]!=2'b00));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_3_nl
      = conv_u2u_17_18(~ (in_data[78:62])) + conv_u2u_1_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_3_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_3_nl
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_3_nl[17:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_4_mx0
      = MUX_v_18_2_2(({1'b0 , (in_data[78:62])}), ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_3_nl,
      in_data[79]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_7_nl
      = MUX_v_10_12_2(10'b0000000001, 10'b0011111100, 10'b0111011100, 10'b1010001101,
      10'b1100001111, 10'b1101100111, 10'b1110100000, 10'b1111000101, 10'b1111011100,
      10'b1111101010, 10'b1111110011, 10'b1111111000, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_4_mx0[13:10]);
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_4_mx0w2_20_10
      = conv_u2u_8_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_28[17:10])
      + conv_u2u_10_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_7_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_4_mx0w2_20_10
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_4_mx0w2_20_10[10:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_4_nl
      = ~((in_data[81:80]!=2'b00));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_4_nl
      = conv_u2u_17_18(~ (in_data[98:82])) + conv_u2u_1_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_4_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_4_nl
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_4_nl[17:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_5_mx0
      = MUX_v_18_2_2(({1'b0 , (in_data[98:82])}), ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_4_nl,
      in_data[99]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_9_nl
      = MUX_v_10_12_2(10'b0000000001, 10'b0011111100, 10'b0111011100, 10'b1010001101,
      10'b1100001111, 10'b1101100111, 10'b1110100000, 10'b1111000101, 10'b1111011100,
      10'b1111101010, 10'b1111110011, 10'b1111111000, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_5_mx0[13:10]);
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_5_mx0w2_20_10
      = conv_u2u_8_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_27[17:10])
      + conv_u2u_10_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_9_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_5_mx0w2_20_10
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_5_mx0w2_20_10[10:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_5_nl
      = ~((in_data[101:100]!=2'b00));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_5_nl
      = conv_u2u_17_18(~ (in_data[118:102])) + conv_u2u_1_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_5_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_5_nl
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_5_nl[17:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_6_mx0
      = MUX_v_18_2_2(({1'b0 , (in_data[118:102])}), ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_5_nl,
      in_data[119]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_11_nl
      = MUX_v_10_12_2(10'b0000000001, 10'b0011111100, 10'b0111011100, 10'b1010001101,
      10'b1100001111, 10'b1101100111, 10'b1110100000, 10'b1111000101, 10'b1111011100,
      10'b1111101010, 10'b1111110011, 10'b1111111000, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_6_mx0[13:10]);
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_6_mx0w2_20_10
      = conv_u2u_8_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_26[17:10])
      + conv_u2u_10_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_11_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_6_mx0w2_20_10
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_6_mx0w2_20_10[10:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_6_nl
      = ~((in_data[121:120]!=2'b00));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_6_nl
      = conv_u2u_17_18(~ (in_data[138:122])) + conv_u2u_1_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_6_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_6_nl
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_6_nl[17:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_7_mx0
      = MUX_v_18_2_2(({1'b0 , (in_data[138:122])}), ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_6_nl,
      in_data[139]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_13_nl
      = MUX_v_10_12_2(10'b0000000001, 10'b0011111100, 10'b0111011100, 10'b1010001101,
      10'b1100001111, 10'b1101100111, 10'b1110100000, 10'b1111000101, 10'b1111011100,
      10'b1111101010, 10'b1111110011, 10'b1111111000, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_7_mx0[13:10]);
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_7_mx0w2_20_10
      = conv_u2u_8_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_25[17:10])
      + conv_u2u_10_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_13_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_7_mx0w2_20_10
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_7_mx0w2_20_10[10:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_7_nl
      = ~((in_data[141:140]!=2'b00));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_7_nl
      = conv_u2u_17_18(~ (in_data[158:142])) + conv_u2u_1_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_7_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_7_nl
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_7_nl[17:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_8_mx0
      = MUX_v_18_2_2(({1'b0 , (in_data[158:142])}), ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_7_nl,
      in_data[159]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_15_nl
      = MUX_v_10_12_2(10'b0000000001, 10'b0011111100, 10'b0111011100, 10'b1010001101,
      10'b1100001111, 10'b1101100111, 10'b1110100000, 10'b1111000101, 10'b1111011100,
      10'b1111101010, 10'b1111110011, 10'b1111111000, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_8_mx0[13:10]);
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_8_mx0w2_20_10
      = conv_u2u_8_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_24[17:10])
      + conv_u2u_10_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_15_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_8_mx0w2_20_10
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_8_mx0w2_20_10[10:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_8_nl
      = ~((in_data[161:160]!=2'b00));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_8_nl
      = conv_u2u_17_18(~ (in_data[178:162])) + conv_u2u_1_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_8_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_8_nl
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_8_nl[17:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_9_mx0
      = MUX_v_18_2_2(({1'b0 , (in_data[178:162])}), ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_8_nl,
      in_data[179]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_17_nl
      = MUX_v_10_12_2(10'b0000000001, 10'b0011111100, 10'b0111011100, 10'b1010001101,
      10'b1100001111, 10'b1101100111, 10'b1110100000, 10'b1111000101, 10'b1111011100,
      10'b1111101010, 10'b1111110011, 10'b1111111000, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_9_mx0[13:10]);
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_9_mx0w2_20_10
      = conv_u2u_8_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_23[17:10])
      + conv_u2u_10_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_17_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_9_mx0w2_20_10
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_9_mx0w2_20_10[10:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_9_nl
      = ~((in_data[181:180]!=2'b00));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_9_nl
      = conv_u2u_17_18(~ (in_data[198:182])) + conv_u2u_1_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_9_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_9_nl
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_9_nl[17:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_10_mx0
      = MUX_v_18_2_2(({1'b0 , (in_data[198:182])}), ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_9_nl,
      in_data[199]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_19_nl
      = MUX_v_10_12_2(10'b0000000001, 10'b0011111100, 10'b0111011100, 10'b1010001101,
      10'b1100001111, 10'b1101100111, 10'b1110100000, 10'b1111000101, 10'b1111011100,
      10'b1111101010, 10'b1111110011, 10'b1111111000, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_10_mx0[13:10]);
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_10_mx0w2_20_10
      = conv_u2u_8_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_22[17:10])
      + conv_u2u_10_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_19_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_10_mx0w2_20_10
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_10_mx0w2_20_10[10:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_10_nl
      = ~((in_data[201:200]!=2'b00));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_10_nl
      = conv_u2u_17_18(~ (in_data[218:202])) + conv_u2u_1_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_10_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_10_nl
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_10_nl[17:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_11_mx0
      = MUX_v_18_2_2(({1'b0 , (in_data[218:202])}), ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_10_nl,
      in_data[219]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_21_nl
      = MUX_v_10_12_2(10'b0000000001, 10'b0011111100, 10'b0111011100, 10'b1010001101,
      10'b1100001111, 10'b1101100111, 10'b1110100000, 10'b1111000101, 10'b1111011100,
      10'b1111101010, 10'b1111110011, 10'b1111111000, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_11_mx0[13:10]);
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_11_mx0w2_20_10
      = conv_u2u_8_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_21[17:10])
      + conv_u2u_10_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_21_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_11_mx0w2_20_10
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_11_mx0w2_20_10[10:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_11_nl
      = ~((in_data[221:220]!=2'b00));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_11_nl
      = conv_u2u_17_18(~ (in_data[238:222])) + conv_u2u_1_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_11_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_11_nl
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_11_nl[17:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_12_mx0
      = MUX_v_18_2_2(({1'b0 , (in_data[238:222])}), ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_11_nl,
      in_data[239]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_23_nl
      = MUX_v_10_12_2(10'b0000000001, 10'b0011111100, 10'b0111011100, 10'b1010001101,
      10'b1100001111, 10'b1101100111, 10'b1110100000, 10'b1111000101, 10'b1111011100,
      10'b1111101010, 10'b1111110011, 10'b1111111000, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_12_mx0[13:10]);
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_12_mx0w2_20_10
      = conv_u2u_8_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_20[17:10])
      + conv_u2u_10_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_23_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_12_mx0w2_20_10
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_12_mx0w2_20_10[10:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_12_nl
      = ~((in_data[241:240]!=2'b00));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_12_nl
      = conv_u2u_17_18(~ (in_data[258:242])) + conv_u2u_1_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_12_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_12_nl
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_12_nl[17:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_13_mx0
      = MUX_v_18_2_2(({1'b0 , (in_data[258:242])}), ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_12_nl,
      in_data[259]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_25_nl
      = MUX_v_10_12_2(10'b0000000001, 10'b0011111100, 10'b0111011100, 10'b1010001101,
      10'b1100001111, 10'b1101100111, 10'b1110100000, 10'b1111000101, 10'b1111011100,
      10'b1111101010, 10'b1111110011, 10'b1111111000, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_13_mx0[13:10]);
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_13_mx0w2_20_10
      = conv_u2u_8_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_19[17:10])
      + conv_u2u_10_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_25_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_13_mx0w2_20_10
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_13_mx0w2_20_10[10:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_13_nl
      = ~((in_data[261:260]!=2'b00));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_13_nl
      = conv_u2u_17_18(~ (in_data[278:262])) + conv_u2u_1_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_13_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_13_nl
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_13_nl[17:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_14_mx0
      = MUX_v_18_2_2(({1'b0 , (in_data[278:262])}), ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_13_nl,
      in_data[279]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_27_nl
      = MUX_v_10_12_2(10'b0000000001, 10'b0011111100, 10'b0111011100, 10'b1010001101,
      10'b1100001111, 10'b1101100111, 10'b1110100000, 10'b1111000101, 10'b1111011100,
      10'b1111101010, 10'b1111110011, 10'b1111111000, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_14_mx0[13:10]);
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_14_mx0w2_20_10
      = conv_u2u_8_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_18[17:10])
      + conv_u2u_10_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_27_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_14_mx0w2_20_10
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_14_mx0w2_20_10[10:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_14_nl
      = ~((in_data[281:280]!=2'b00));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_14_nl
      = conv_u2u_17_18(~ (in_data[298:282])) + conv_u2u_1_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_14_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_14_nl
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_14_nl[17:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_15_mx0
      = MUX_v_18_2_2(({1'b0 , (in_data[298:282])}), ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_14_nl,
      in_data[299]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_29_nl
      = MUX_v_10_12_2(10'b0000000001, 10'b0011111100, 10'b0111011100, 10'b1010001101,
      10'b1100001111, 10'b1101100111, 10'b1110100000, 10'b1111000101, 10'b1111011100,
      10'b1111101010, 10'b1111110011, 10'b1111111000, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_15_mx0[13:10]);
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_15_mx0w2_20_10
      = conv_u2u_8_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_17[17:10])
      + conv_u2u_10_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_29_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_15_mx0w2_20_10
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_15_mx0w2_20_10[10:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_15_nl
      = ~((in_data[301:300]!=2'b00));
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_15_nl
      = conv_u2u_17_18(~ (in_data[318:302])) + conv_u2u_1_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_nor_15_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_15_nl
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_15_nl[17:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_mx0
      = MUX_v_18_2_2(({1'b0 , (in_data[318:302])}), ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qelse_acc_15_nl,
      in_data[319]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_31_nl
      = MUX_v_10_12_2(10'b0000000001, 10'b0011111100, 10'b0111011100, 10'b1010001101,
      10'b1100001111, 10'b1101100111, 10'b1110100000, 10'b1111000101, 10'b1111011100,
      10'b1111101010, 10'b1111110011, 10'b1111111000, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_mx0[13:10]);
  assign nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mx0w2_20_10
      = conv_u2u_8_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_16[17:10])
      + conv_u2u_10_11(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_31_nl);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mx0w2_20_10
      = nl_ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mx0w2_20_10[10:0];
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_33_nl
      = MUX_v_8_12_2(8'b11111011, 8'b11100000, 8'b10110001, 8'b10000001, 8'b01011000,
      8'b00111001, 8'b00100101, 8'b00010111, 8'b00001110, 8'b00001001, 8'b00000101,
      8'b00000011, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_mx0[13:10]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_16
      = conv_u2u_18_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_33_nl
      * (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_mx0[9:0]));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_34_nl
      = MUX_v_8_12_2(8'b11111011, 8'b11100000, 8'b10110001, 8'b10000001, 8'b01011000,
      8'b00111001, 8'b00100101, 8'b00010111, 8'b00001110, 8'b00001001, 8'b00000101,
      8'b00000011, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_15_mx0[13:10]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_17
      = conv_u2u_18_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_34_nl
      * (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_15_mx0[9:0]));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_35_nl
      = MUX_v_8_12_2(8'b11111011, 8'b11100000, 8'b10110001, 8'b10000001, 8'b01011000,
      8'b00111001, 8'b00100101, 8'b00010111, 8'b00001110, 8'b00001001, 8'b00000101,
      8'b00000011, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_14_mx0[13:10]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_18
      = conv_u2u_18_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_35_nl
      * (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_14_mx0[9:0]));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_36_nl
      = MUX_v_8_12_2(8'b11111011, 8'b11100000, 8'b10110001, 8'b10000001, 8'b01011000,
      8'b00111001, 8'b00100101, 8'b00010111, 8'b00001110, 8'b00001001, 8'b00000101,
      8'b00000011, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_13_mx0[13:10]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_19
      = conv_u2u_18_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_36_nl
      * (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_13_mx0[9:0]));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_37_nl
      = MUX_v_8_12_2(8'b11111011, 8'b11100000, 8'b10110001, 8'b10000001, 8'b01011000,
      8'b00111001, 8'b00100101, 8'b00010111, 8'b00001110, 8'b00001001, 8'b00000101,
      8'b00000011, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_12_mx0[13:10]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_20
      = conv_u2u_18_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_37_nl
      * (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_12_mx0[9:0]));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_38_nl
      = MUX_v_8_12_2(8'b11111011, 8'b11100000, 8'b10110001, 8'b10000001, 8'b01011000,
      8'b00111001, 8'b00100101, 8'b00010111, 8'b00001110, 8'b00001001, 8'b00000101,
      8'b00000011, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_11_mx0[13:10]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_21
      = conv_u2u_18_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_38_nl
      * (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_11_mx0[9:0]));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_39_nl
      = MUX_v_8_12_2(8'b11111011, 8'b11100000, 8'b10110001, 8'b10000001, 8'b01011000,
      8'b00111001, 8'b00100101, 8'b00010111, 8'b00001110, 8'b00001001, 8'b00000101,
      8'b00000011, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_10_mx0[13:10]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_22
      = conv_u2u_18_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_39_nl
      * (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_10_mx0[9:0]));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_40_nl
      = MUX_v_8_12_2(8'b11111011, 8'b11100000, 8'b10110001, 8'b10000001, 8'b01011000,
      8'b00111001, 8'b00100101, 8'b00010111, 8'b00001110, 8'b00001001, 8'b00000101,
      8'b00000011, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_9_mx0[13:10]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_23
      = conv_u2u_18_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_40_nl
      * (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_9_mx0[9:0]));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_41_nl
      = MUX_v_8_12_2(8'b11111011, 8'b11100000, 8'b10110001, 8'b10000001, 8'b01011000,
      8'b00111001, 8'b00100101, 8'b00010111, 8'b00001110, 8'b00001001, 8'b00000101,
      8'b00000011, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_8_mx0[13:10]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_24
      = conv_u2u_18_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_41_nl
      * (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_8_mx0[9:0]));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_42_nl
      = MUX_v_8_12_2(8'b11111011, 8'b11100000, 8'b10110001, 8'b10000001, 8'b01011000,
      8'b00111001, 8'b00100101, 8'b00010111, 8'b00001110, 8'b00001001, 8'b00000101,
      8'b00000011, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_7_mx0[13:10]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_25
      = conv_u2u_18_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_42_nl
      * (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_7_mx0[9:0]));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_43_nl
      = MUX_v_8_12_2(8'b11111011, 8'b11100000, 8'b10110001, 8'b10000001, 8'b01011000,
      8'b00111001, 8'b00100101, 8'b00010111, 8'b00001110, 8'b00001001, 8'b00000101,
      8'b00000011, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_6_mx0[13:10]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_26
      = conv_u2u_18_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_43_nl
      * (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_6_mx0[9:0]));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_44_nl
      = MUX_v_8_12_2(8'b11111011, 8'b11100000, 8'b10110001, 8'b10000001, 8'b01011000,
      8'b00111001, 8'b00100101, 8'b00010111, 8'b00001110, 8'b00001001, 8'b00000101,
      8'b00000011, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_5_mx0[13:10]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_27
      = conv_u2u_18_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_44_nl
      * (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_5_mx0[9:0]));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_45_nl
      = MUX_v_8_12_2(8'b11111011, 8'b11100000, 8'b10110001, 8'b10000001, 8'b01011000,
      8'b00111001, 8'b00100101, 8'b00010111, 8'b00001110, 8'b00001001, 8'b00000101,
      8'b00000011, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_4_mx0[13:10]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_28
      = conv_u2u_18_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_45_nl
      * (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_4_mx0[9:0]));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_46_nl
      = MUX_v_8_12_2(8'b11111011, 8'b11100000, 8'b10110001, 8'b10000001, 8'b01011000,
      8'b00111001, 8'b00100101, 8'b00010111, 8'b00001110, 8'b00001001, 8'b00000101,
      8'b00000011, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_3_mx0[13:10]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_29
      = conv_u2u_18_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_46_nl
      * (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_3_mx0[9:0]));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_2_nl
      = MUX_v_8_12_2(8'b11111011, 8'b11100000, 8'b10110001, 8'b10000001, 8'b01011000,
      8'b00111001, 8'b00100101, 8'b00010111, 8'b00001110, 8'b00001001, 8'b00000101,
      8'b00000011, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_2_mx0[13:10]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_30
      = conv_u2u_18_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_2_nl
      * (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_2_mx0[9:0]));
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_47_nl
      = MUX_v_8_12_2(8'b11111011, 8'b11100000, 8'b10110001, 8'b10000001, 8'b01011000,
      8'b00111001, 8'b00100101, 8'b00010111, 8'b00001110, 8'b00001001, 8'b00000101,
      8'b00000011, ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_1_mx0[13:10]);
  assign ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mul_sdt_31
      = conv_u2u_18_18(ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_output_pwl_mux_47_nl
      * (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_1_mx0[9:0]));
  assign nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_15_nl = (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_mx0[17:12])
      + 6'b111101;
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_15_nl = nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_15_nl[5:0];
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_15_itm_5_1 = readslicef_6_1_5(operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_15_nl);
  assign nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_14_nl = (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_15_mx0[17:12])
      + 6'b111101;
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_14_nl = nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_14_nl[5:0];
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_14_itm_5_1 = readslicef_6_1_5(operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_14_nl);
  assign nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_13_nl = (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_14_mx0[17:12])
      + 6'b111101;
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_13_nl = nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_13_nl[5:0];
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_13_itm_5_1 = readslicef_6_1_5(operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_13_nl);
  assign nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_12_nl = (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_13_mx0[17:12])
      + 6'b111101;
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_12_nl = nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_12_nl[5:0];
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_12_itm_5_1 = readslicef_6_1_5(operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_12_nl);
  assign nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_11_nl = (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_12_mx0[17:12])
      + 6'b111101;
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_11_nl = nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_11_nl[5:0];
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_11_itm_5_1 = readslicef_6_1_5(operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_11_nl);
  assign nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_10_nl = (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_11_mx0[17:12])
      + 6'b111101;
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_10_nl = nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_10_nl[5:0];
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_10_itm_5_1 = readslicef_6_1_5(operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_10_nl);
  assign nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_9_nl = (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_10_mx0[17:12])
      + 6'b111101;
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_9_nl = nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_9_nl[5:0];
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_9_itm_5_1 = readslicef_6_1_5(operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_9_nl);
  assign nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_8_nl = (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_9_mx0[17:12])
      + 6'b111101;
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_8_nl = nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_8_nl[5:0];
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_8_itm_5_1 = readslicef_6_1_5(operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_8_nl);
  assign nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_7_nl = (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_8_mx0[17:12])
      + 6'b111101;
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_7_nl = nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_7_nl[5:0];
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_7_itm_5_1 = readslicef_6_1_5(operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_7_nl);
  assign nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_6_nl = (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_7_mx0[17:12])
      + 6'b111101;
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_6_nl = nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_6_nl[5:0];
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_6_itm_5_1 = readslicef_6_1_5(operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_6_nl);
  assign nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_5_nl = (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_6_mx0[17:12])
      + 6'b111101;
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_5_nl = nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_5_nl[5:0];
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_5_itm_5_1 = readslicef_6_1_5(operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_5_nl);
  assign nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_4_nl = (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_5_mx0[17:12])
      + 6'b111101;
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_4_nl = nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_4_nl[5:0];
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_4_itm_5_1 = readslicef_6_1_5(operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_4_nl);
  assign nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_3_nl = (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_4_mx0[17:12])
      + 6'b111101;
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_3_nl = nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_3_nl[5:0];
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_3_itm_5_1 = readslicef_6_1_5(operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_3_nl);
  assign nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_2_nl = (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_3_mx0[17:12])
      + 6'b111101;
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_2_nl = nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_2_nl[5:0];
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_2_itm_5_1 = readslicef_6_1_5(operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_2_nl);
  assign nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_1_nl = (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_2_mx0[17:12])
      + 6'b111101;
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_1_nl = nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_1_nl[5:0];
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_1_itm_5_1 = readslicef_6_1_5(operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_1_nl);
  assign nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_nl = (ac_math_ac_tanh_pwl_AC_TRN_20_6_true_AC_TRN_AC_WRAP_20_6_false_AC_TRN_AC_WRAP_if_1_qr_19_2_1_mx0[17:12])
      + 6'b111101;
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_nl = nl_operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_nl[5:0];
  assign operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_itm_5_1 = readslicef_6_1_5(operator_20_6_false_AC_TRN_AC_WRAP_2_false_acc_nl);

  function automatic [14:0] MUX1HOT_v_15_3_2;
    input [14:0] input_2;
    input [14:0] input_1;
    input [14:0] input_0;
    input [2:0] sel;
    reg [14:0] result;
  begin
    result = input_0 & {15{sel[0]}};
    result = result | ( input_1 & {15{sel[1]}});
    result = result | ( input_2 & {15{sel[2]}});
    MUX1HOT_v_15_3_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_12_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [9:0] input_2;
    input [9:0] input_3;
    input [9:0] input_4;
    input [9:0] input_5;
    input [9:0] input_6;
    input [9:0] input_7;
    input [9:0] input_8;
    input [9:0] input_9;
    input [9:0] input_10;
    input [9:0] input_11;
    input [3:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      default : begin
        result = input_11;
      end
    endcase
    MUX_v_10_12_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [0:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [17:0] MUX_v_18_2_2;
    input [17:0] input_0;
    input [17:0] input_1;
    input [0:0] sel;
    reg [17:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_18_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_12_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [7:0] input_8;
    input [7:0] input_9;
    input [7:0] input_10;
    input [7:0] input_11;
    input [3:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      default : begin
        result = input_11;
      end
    endcase
    MUX_v_8_12_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_6_1_5;
    input [5:0] vector;
    reg [5:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_6_1_5 = tmp[0:0];
  end
  endfunction


  function automatic [19:0] signext_20_15;
    input [14:0] vector;
  begin
    signext_20_15= {{5{vector[14]}}, vector};
  end
  endfunction


  function automatic [319:0] signext_320_315;
    input [314:0] vector;
  begin
    signext_320_315= {{5{vector[314]}}, vector};
  end
  endfunction


  function automatic [14:0] conv_u2s_1_15 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_15 = {{14{1'b0}}, vector};
  end
  endfunction


  function automatic [17:0] conv_u2u_1_18 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_18 = {{17{1'b0}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_8_11 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_11 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction


  function automatic [17:0] conv_u2u_17_18 ;
    input [16:0]  vector ;
  begin
    conv_u2u_17_18 = {1'b0, vector};
  end
  endfunction


  function automatic [17:0] conv_u2u_18_18 ;
    input [17:0]  vector ;
  begin
    conv_u2u_18_18 = vector;
  end
  endfunction

endmodule




//------> ./ActUnit_Relu.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   huaixil@sat8
//  Generated date: Fri Apr  8 23:10:52 2022
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Relu
// ------------------------------------------------------------------


module ActUnit_Relu (
  in_data, out_data
);
  input [319:0] in_data;
  output [319:0] out_data;


  wire[18:0] for_if_for_if_and_nl;
  wire[0:0] for_if_not_nl;
  wire[18:0] for_if_for_if_and_1_nl;
  wire[0:0] for_if_not_1_nl;
  wire[18:0] for_if_for_if_and_2_nl;
  wire[0:0] for_if_not_2_nl;
  wire[18:0] for_if_for_if_and_3_nl;
  wire[0:0] for_if_not_3_nl;
  wire[18:0] for_if_for_if_and_4_nl;
  wire[0:0] for_if_not_4_nl;
  wire[18:0] for_if_for_if_and_5_nl;
  wire[0:0] for_if_not_5_nl;
  wire[18:0] for_if_for_if_and_6_nl;
  wire[0:0] for_if_not_6_nl;
  wire[18:0] for_if_for_if_and_7_nl;
  wire[0:0] for_if_not_7_nl;
  wire[18:0] for_if_for_if_and_8_nl;
  wire[0:0] for_if_not_8_nl;
  wire[18:0] for_if_for_if_and_9_nl;
  wire[0:0] for_if_not_9_nl;
  wire[18:0] for_if_for_if_and_10_nl;
  wire[0:0] for_if_not_10_nl;
  wire[18:0] for_if_for_if_and_11_nl;
  wire[0:0] for_if_not_11_nl;
  wire[18:0] for_if_for_if_and_12_nl;
  wire[0:0] for_if_not_12_nl;
  wire[18:0] for_if_for_if_and_13_nl;
  wire[0:0] for_if_not_13_nl;
  wire[18:0] for_if_for_if_and_14_nl;
  wire[0:0] for_if_not_14_nl;
  wire[18:0] for_if_for_if_and_15_nl;
  wire[0:0] for_if_not_15_nl;

  // Interconnect Declarations for Component Instantiations
  assign for_if_not_nl = ~ (in_data[319]);
  assign for_if_for_if_and_nl = MUX_v_19_2_2(19'b0000000000000000000, (in_data[318:300]),
      for_if_not_nl);
  assign for_if_not_1_nl = ~ (in_data[299]);
  assign for_if_for_if_and_1_nl = MUX_v_19_2_2(19'b0000000000000000000, (in_data[298:280]),
      for_if_not_1_nl);
  assign for_if_not_2_nl = ~ (in_data[279]);
  assign for_if_for_if_and_2_nl = MUX_v_19_2_2(19'b0000000000000000000, (in_data[278:260]),
      for_if_not_2_nl);
  assign for_if_not_3_nl = ~ (in_data[259]);
  assign for_if_for_if_and_3_nl = MUX_v_19_2_2(19'b0000000000000000000, (in_data[258:240]),
      for_if_not_3_nl);
  assign for_if_not_4_nl = ~ (in_data[239]);
  assign for_if_for_if_and_4_nl = MUX_v_19_2_2(19'b0000000000000000000, (in_data[238:220]),
      for_if_not_4_nl);
  assign for_if_not_5_nl = ~ (in_data[219]);
  assign for_if_for_if_and_5_nl = MUX_v_19_2_2(19'b0000000000000000000, (in_data[218:200]),
      for_if_not_5_nl);
  assign for_if_not_6_nl = ~ (in_data[199]);
  assign for_if_for_if_and_6_nl = MUX_v_19_2_2(19'b0000000000000000000, (in_data[198:180]),
      for_if_not_6_nl);
  assign for_if_not_7_nl = ~ (in_data[179]);
  assign for_if_for_if_and_7_nl = MUX_v_19_2_2(19'b0000000000000000000, (in_data[178:160]),
      for_if_not_7_nl);
  assign for_if_not_8_nl = ~ (in_data[159]);
  assign for_if_for_if_and_8_nl = MUX_v_19_2_2(19'b0000000000000000000, (in_data[158:140]),
      for_if_not_8_nl);
  assign for_if_not_9_nl = ~ (in_data[139]);
  assign for_if_for_if_and_9_nl = MUX_v_19_2_2(19'b0000000000000000000, (in_data[138:120]),
      for_if_not_9_nl);
  assign for_if_not_10_nl = ~ (in_data[119]);
  assign for_if_for_if_and_10_nl = MUX_v_19_2_2(19'b0000000000000000000, (in_data[118:100]),
      for_if_not_10_nl);
  assign for_if_not_11_nl = ~ (in_data[99]);
  assign for_if_for_if_and_11_nl = MUX_v_19_2_2(19'b0000000000000000000, (in_data[98:80]),
      for_if_not_11_nl);
  assign for_if_not_12_nl = ~ (in_data[79]);
  assign for_if_for_if_and_12_nl = MUX_v_19_2_2(19'b0000000000000000000, (in_data[78:60]),
      for_if_not_12_nl);
  assign for_if_not_13_nl = ~ (in_data[59]);
  assign for_if_for_if_and_13_nl = MUX_v_19_2_2(19'b0000000000000000000, (in_data[58:40]),
      for_if_not_13_nl);
  assign for_if_not_14_nl = ~ (in_data[39]);
  assign for_if_for_if_and_14_nl = MUX_v_19_2_2(19'b0000000000000000000, (in_data[38:20]),
      for_if_not_14_nl);
  assign for_if_not_15_nl = ~ (in_data[19]);
  assign for_if_for_if_and_15_nl = MUX_v_19_2_2(19'b0000000000000000000, (in_data[18:0]),
      for_if_not_15_nl);
  assign out_data = {1'b0 , for_if_for_if_and_nl , 1'b0 , for_if_for_if_and_1_nl
      , 1'b0 , for_if_for_if_and_2_nl , 1'b0 , for_if_for_if_and_3_nl , 1'b0 , for_if_for_if_and_4_nl
      , 1'b0 , for_if_for_if_and_5_nl , 1'b0 , for_if_for_if_and_6_nl , 1'b0 , for_if_for_if_and_7_nl
      , 1'b0 , for_if_for_if_and_8_nl , 1'b0 , for_if_for_if_and_9_nl , 1'b0 , for_if_for_if_and_10_nl
      , 1'b0 , for_if_for_if_and_11_nl , 1'b0 , for_if_for_if_and_12_nl , 1'b0 ,
      for_if_for_if_and_13_nl , 1'b0 , for_if_for_if_and_14_nl , 1'b0 , for_if_for_if_and_15_nl};

  function automatic [18:0] MUX_v_19_2_2;
    input [18:0] input_0;
    input [18:0] input_1;
    input [0:0] sel;
    reg [18:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_19_2_2 = result;
  end
  endfunction

endmodule




//------> ./ActUnit_OneX.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   huaixil@sat8
//  Generated date: Fri Apr  8 23:10:50 2022
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    OneX
// ------------------------------------------------------------------


module ActUnit_OneX (
  in_data, out_data
);
  input [319:0] in_data;
  output [319:0] out_data;


  wire[19:0] operator_20_true_acc_15_nl;
  wire[20:0] nl_operator_20_true_acc_15_nl;
  wire[19:0] operator_20_true_acc_14_nl;
  wire[20:0] nl_operator_20_true_acc_14_nl;
  wire[19:0] operator_20_true_acc_13_nl;
  wire[20:0] nl_operator_20_true_acc_13_nl;
  wire[19:0] operator_20_true_acc_12_nl;
  wire[20:0] nl_operator_20_true_acc_12_nl;
  wire[19:0] operator_20_true_acc_11_nl;
  wire[20:0] nl_operator_20_true_acc_11_nl;
  wire[19:0] operator_20_true_acc_10_nl;
  wire[20:0] nl_operator_20_true_acc_10_nl;
  wire[19:0] operator_20_true_acc_9_nl;
  wire[20:0] nl_operator_20_true_acc_9_nl;
  wire[19:0] operator_20_true_acc_8_nl;
  wire[20:0] nl_operator_20_true_acc_8_nl;
  wire[19:0] operator_20_true_acc_7_nl;
  wire[20:0] nl_operator_20_true_acc_7_nl;
  wire[19:0] operator_20_true_acc_6_nl;
  wire[20:0] nl_operator_20_true_acc_6_nl;
  wire[19:0] operator_20_true_acc_5_nl;
  wire[20:0] nl_operator_20_true_acc_5_nl;
  wire[19:0] operator_20_true_acc_4_nl;
  wire[20:0] nl_operator_20_true_acc_4_nl;
  wire[19:0] operator_20_true_acc_3_nl;
  wire[20:0] nl_operator_20_true_acc_3_nl;
  wire[19:0] operator_20_true_acc_2_nl;
  wire[20:0] nl_operator_20_true_acc_2_nl;
  wire[19:0] operator_20_true_acc_1_nl;
  wire[20:0] nl_operator_20_true_acc_1_nl;
  wire[19:0] operator_20_true_acc_nl;
  wire[20:0] nl_operator_20_true_acc_nl;

  // Interconnect Declarations for Component Instantiations
  assign nl_operator_20_true_acc_15_nl = (~ (in_data[319:300])) + 20'b00000100000000000001;
  assign operator_20_true_acc_15_nl = nl_operator_20_true_acc_15_nl[19:0];
  assign nl_operator_20_true_acc_14_nl = (~ (in_data[299:280])) + 20'b00000100000000000001;
  assign operator_20_true_acc_14_nl = nl_operator_20_true_acc_14_nl[19:0];
  assign nl_operator_20_true_acc_13_nl = (~ (in_data[279:260])) + 20'b00000100000000000001;
  assign operator_20_true_acc_13_nl = nl_operator_20_true_acc_13_nl[19:0];
  assign nl_operator_20_true_acc_12_nl = (~ (in_data[259:240])) + 20'b00000100000000000001;
  assign operator_20_true_acc_12_nl = nl_operator_20_true_acc_12_nl[19:0];
  assign nl_operator_20_true_acc_11_nl = (~ (in_data[239:220])) + 20'b00000100000000000001;
  assign operator_20_true_acc_11_nl = nl_operator_20_true_acc_11_nl[19:0];
  assign nl_operator_20_true_acc_10_nl = (~ (in_data[219:200])) + 20'b00000100000000000001;
  assign operator_20_true_acc_10_nl = nl_operator_20_true_acc_10_nl[19:0];
  assign nl_operator_20_true_acc_9_nl = (~ (in_data[199:180])) + 20'b00000100000000000001;
  assign operator_20_true_acc_9_nl = nl_operator_20_true_acc_9_nl[19:0];
  assign nl_operator_20_true_acc_8_nl = (~ (in_data[179:160])) + 20'b00000100000000000001;
  assign operator_20_true_acc_8_nl = nl_operator_20_true_acc_8_nl[19:0];
  assign nl_operator_20_true_acc_7_nl = (~ (in_data[159:140])) + 20'b00000100000000000001;
  assign operator_20_true_acc_7_nl = nl_operator_20_true_acc_7_nl[19:0];
  assign nl_operator_20_true_acc_6_nl = (~ (in_data[139:120])) + 20'b00000100000000000001;
  assign operator_20_true_acc_6_nl = nl_operator_20_true_acc_6_nl[19:0];
  assign nl_operator_20_true_acc_5_nl = (~ (in_data[119:100])) + 20'b00000100000000000001;
  assign operator_20_true_acc_5_nl = nl_operator_20_true_acc_5_nl[19:0];
  assign nl_operator_20_true_acc_4_nl = (~ (in_data[99:80])) + 20'b00000100000000000001;
  assign operator_20_true_acc_4_nl = nl_operator_20_true_acc_4_nl[19:0];
  assign nl_operator_20_true_acc_3_nl = (~ (in_data[79:60])) + 20'b00000100000000000001;
  assign operator_20_true_acc_3_nl = nl_operator_20_true_acc_3_nl[19:0];
  assign nl_operator_20_true_acc_2_nl = (~ (in_data[59:40])) + 20'b00000100000000000001;
  assign operator_20_true_acc_2_nl = nl_operator_20_true_acc_2_nl[19:0];
  assign nl_operator_20_true_acc_1_nl = (~ (in_data[39:20])) + 20'b00000100000000000001;
  assign operator_20_true_acc_1_nl = nl_operator_20_true_acc_1_nl[19:0];
  assign nl_operator_20_true_acc_nl = (~ (in_data[19:0])) + 20'b00000100000000000001;
  assign operator_20_true_acc_nl = nl_operator_20_true_acc_nl[19:0];
  assign out_data = {operator_20_true_acc_15_nl , operator_20_true_acc_14_nl , operator_20_true_acc_13_nl
      , operator_20_true_acc_12_nl , operator_20_true_acc_11_nl , operator_20_true_acc_10_nl
      , operator_20_true_acc_9_nl , operator_20_true_acc_8_nl , operator_20_true_acc_7_nl
      , operator_20_true_acc_6_nl , operator_20_true_acc_5_nl , operator_20_true_acc_4_nl
      , operator_20_true_acc_3_nl , operator_20_true_acc_2_nl , operator_20_true_acc_1_nl
      , operator_20_true_acc_nl};
endmodule




//------> ./ActUnit_Adpfloat2Fixed_mgc_shift_l_beh_v5.v 
module ActUnit_Adpfloat2Fixed_mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./ActUnit_Adpfloat2Fixed.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   huaixil@sat8
//  Generated date: Fri Apr  8 23:10:39 2022
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Adpfloat2Fixed
// ------------------------------------------------------------------


module ActUnit_Adpfloat2Fixed (
  in_data, out_data, adpfloat_bias
);
  input [127:0] in_data;
  output [319:0] out_data;
  input [2:0] adpfloat_bias;


  // Interconnect Declarations
  wire [18:0] input_adpfloat_to_fixed_20U_14U_lshift_psp_31;
  wire [18:0] input_adpfloat_to_fixed_20U_14U_lshift_psp_30;
  wire [18:0] input_adpfloat_to_fixed_20U_14U_lshift_psp_29;
  wire [18:0] input_adpfloat_to_fixed_20U_14U_lshift_psp_28;
  wire [18:0] input_adpfloat_to_fixed_20U_14U_lshift_psp_27;
  wire [18:0] input_adpfloat_to_fixed_20U_14U_lshift_psp_26;
  wire [18:0] input_adpfloat_to_fixed_20U_14U_lshift_psp_25;
  wire [18:0] input_adpfloat_to_fixed_20U_14U_lshift_psp_24;
  wire [18:0] input_adpfloat_to_fixed_20U_14U_lshift_psp_23;
  wire [18:0] input_adpfloat_to_fixed_20U_14U_lshift_psp_22;
  wire [18:0] input_adpfloat_to_fixed_20U_14U_lshift_psp_21;
  wire [18:0] input_adpfloat_to_fixed_20U_14U_lshift_psp_20;
  wire [18:0] input_adpfloat_to_fixed_20U_14U_lshift_psp_19;
  wire [18:0] input_adpfloat_to_fixed_20U_14U_lshift_psp_18;
  wire [18:0] input_adpfloat_to_fixed_20U_14U_lshift_psp_17;
  wire [18:0] input_adpfloat_to_fixed_20U_14U_lshift_psp_16;
  wire or_15_tmp;
  wire or_14_tmp;
  wire or_13_tmp;
  wire or_12_tmp;
  wire or_11_tmp;
  wire or_10_tmp;
  wire or_9_tmp;
  wire or_8_tmp;
  wire or_7_tmp;
  wire or_6_tmp;
  wire or_5_tmp;
  wire or_4_tmp;
  wire or_3_tmp;
  wire or_2_tmp;
  wire or_1_tmp;
  wire or_tmp;
  wire input_adpfloat_to_fixed_20U_14U_if_and_ssc;
  wire input_adpfloat_to_fixed_20U_14U_if_and_1_ssc;
  wire input_adpfloat_to_fixed_20U_14U_if_and_2_ssc;
  wire input_adpfloat_to_fixed_20U_14U_if_and_3_ssc;
  wire input_adpfloat_to_fixed_20U_14U_if_and_4_ssc;
  wire input_adpfloat_to_fixed_20U_14U_if_and_5_ssc;
  wire input_adpfloat_to_fixed_20U_14U_if_and_6_ssc;
  wire input_adpfloat_to_fixed_20U_14U_if_and_7_ssc;
  wire input_adpfloat_to_fixed_20U_14U_if_and_8_ssc;
  wire input_adpfloat_to_fixed_20U_14U_if_and_9_ssc;
  wire input_adpfloat_to_fixed_20U_14U_if_and_10_ssc;
  wire input_adpfloat_to_fixed_20U_14U_if_and_11_ssc;
  wire input_adpfloat_to_fixed_20U_14U_if_and_12_ssc;
  wire input_adpfloat_to_fixed_20U_14U_if_and_13_ssc;
  wire input_adpfloat_to_fixed_20U_14U_if_and_14_ssc;
  wire input_adpfloat_to_fixed_20U_14U_if_and_15_ssc;

  wire[19:0] input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_mux_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_1_acc_15_nl;
  wire[19:0] nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_15_nl;
  wire[19:0] input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_1_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_mux_16_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_1_acc_14_nl;
  wire[19:0] nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_14_nl;
  wire[19:0] input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_2_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_mux_17_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_1_acc_13_nl;
  wire[19:0] nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_13_nl;
  wire[19:0] input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_3_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_mux_18_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_1_acc_12_nl;
  wire[19:0] nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_12_nl;
  wire[19:0] input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_4_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_mux_19_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_1_acc_11_nl;
  wire[19:0] nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_11_nl;
  wire[19:0] input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_5_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_mux_20_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_1_acc_10_nl;
  wire[19:0] nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_10_nl;
  wire[19:0] input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_6_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_mux_21_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_1_acc_9_nl;
  wire[19:0] nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_9_nl;
  wire[19:0] input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_7_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_mux_22_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_1_acc_8_nl;
  wire[19:0] nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_8_nl;
  wire[19:0] input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_8_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_mux_23_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_1_acc_7_nl;
  wire[19:0] nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_7_nl;
  wire[19:0] input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_9_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_mux_24_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_1_acc_6_nl;
  wire[19:0] nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_6_nl;
  wire[19:0] input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_10_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_mux_25_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_1_acc_5_nl;
  wire[19:0] nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_5_nl;
  wire[19:0] input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_11_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_mux_26_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_1_acc_4_nl;
  wire[19:0] nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_4_nl;
  wire[19:0] input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_12_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_mux_27_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_1_acc_3_nl;
  wire[19:0] nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_3_nl;
  wire[19:0] input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_13_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_mux_28_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_1_acc_2_nl;
  wire[19:0] nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_2_nl;
  wire[19:0] input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_14_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_mux_29_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_1_acc_1_nl;
  wire[19:0] nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_1_nl;
  wire[19:0] input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_15_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_mux_30_nl;
  wire[18:0] input_adpfloat_to_fixed_20U_14U_if_1_acc_nl;
  wire[19:0] nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_nl;

  // Interconnect Declarations for Component Instantiations
  wire [4:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_rg_a;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_rg_a = {1'b1 , (in_data[3:0])};
  wire [3:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_rg_s;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_rg_s = conv_u2u_3_4(in_data[6:4])
      + conv_u2u_3_4(adpfloat_bias);
  wire [4:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_1_rg_a;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_1_rg_a = {1'b1 , (in_data[11:8])};
  wire [3:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_1_rg_s;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_1_rg_s = conv_u2u_3_4(in_data[14:12])
      + conv_u2u_3_4(adpfloat_bias);
  wire [4:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_2_rg_a;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_2_rg_a = {1'b1 , (in_data[19:16])};
  wire [3:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_2_rg_s;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_2_rg_s = conv_u2u_3_4(in_data[22:20])
      + conv_u2u_3_4(adpfloat_bias);
  wire [4:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_3_rg_a;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_3_rg_a = {1'b1 , (in_data[27:24])};
  wire [3:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_3_rg_s;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_3_rg_s = conv_u2u_3_4(in_data[30:28])
      + conv_u2u_3_4(adpfloat_bias);
  wire [4:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_4_rg_a;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_4_rg_a = {1'b1 , (in_data[35:32])};
  wire [3:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_4_rg_s;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_4_rg_s = conv_u2u_3_4(in_data[38:36])
      + conv_u2u_3_4(adpfloat_bias);
  wire [4:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_5_rg_a;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_5_rg_a = {1'b1 , (in_data[43:40])};
  wire [3:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_5_rg_s;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_5_rg_s = conv_u2u_3_4(in_data[46:44])
      + conv_u2u_3_4(adpfloat_bias);
  wire [4:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_6_rg_a;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_6_rg_a = {1'b1 , (in_data[51:48])};
  wire [3:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_6_rg_s;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_6_rg_s = conv_u2u_3_4(in_data[54:52])
      + conv_u2u_3_4(adpfloat_bias);
  wire [4:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_7_rg_a;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_7_rg_a = {1'b1 , (in_data[59:56])};
  wire [3:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_7_rg_s;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_7_rg_s = conv_u2u_3_4(in_data[62:60])
      + conv_u2u_3_4(adpfloat_bias);
  wire [4:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_8_rg_a;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_8_rg_a = {1'b1 , (in_data[67:64])};
  wire [3:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_8_rg_s;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_8_rg_s = conv_u2u_3_4(in_data[70:68])
      + conv_u2u_3_4(adpfloat_bias);
  wire [4:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_9_rg_a;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_9_rg_a = {1'b1 , (in_data[75:72])};
  wire [3:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_9_rg_s;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_9_rg_s = conv_u2u_3_4(in_data[78:76])
      + conv_u2u_3_4(adpfloat_bias);
  wire [4:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_10_rg_a;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_10_rg_a = {1'b1 , (in_data[83:80])};
  wire [3:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_10_rg_s;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_10_rg_s = conv_u2u_3_4(in_data[86:84])
      + conv_u2u_3_4(adpfloat_bias);
  wire [4:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_11_rg_a;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_11_rg_a = {1'b1 , (in_data[91:88])};
  wire [3:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_11_rg_s;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_11_rg_s = conv_u2u_3_4(in_data[94:92])
      + conv_u2u_3_4(adpfloat_bias);
  wire [4:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_12_rg_a;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_12_rg_a = {1'b1 , (in_data[99:96])};
  wire [3:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_12_rg_s;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_12_rg_s = conv_u2u_3_4(in_data[102:100])
      + conv_u2u_3_4(adpfloat_bias);
  wire [4:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_13_rg_a;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_13_rg_a = {1'b1 , (in_data[107:104])};
  wire [3:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_13_rg_s;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_13_rg_s = conv_u2u_3_4(in_data[110:108])
      + conv_u2u_3_4(adpfloat_bias);
  wire [4:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_14_rg_a;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_14_rg_a = {1'b1 , (in_data[115:112])};
  wire [3:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_14_rg_s;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_14_rg_s = conv_u2u_3_4(in_data[118:116])
      + conv_u2u_3_4(adpfloat_bias);
  wire [4:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_15_rg_a;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_15_rg_a = {1'b1 , (in_data[123:120])};
  wire [3:0] nl_input_adpfloat_to_fixed_20U_14U_lshift_15_rg_s;
  assign nl_input_adpfloat_to_fixed_20U_14U_lshift_15_rg_s = conv_u2u_3_4(in_data[126:124])
      + conv_u2u_3_4(adpfloat_bias);
  ActUnit_Adpfloat2Fixed_mgc_shift_l_v5 #(.width_a(32'sd5),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd19)) input_adpfloat_to_fixed_20U_14U_lshift_rg (
      .a(nl_input_adpfloat_to_fixed_20U_14U_lshift_rg_a[4:0]),
      .s(nl_input_adpfloat_to_fixed_20U_14U_lshift_rg_s[3:0]),
      .z(input_adpfloat_to_fixed_20U_14U_lshift_psp_16)
    );
  ActUnit_Adpfloat2Fixed_mgc_shift_l_v5 #(.width_a(32'sd5),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd19)) input_adpfloat_to_fixed_20U_14U_lshift_1_rg (
      .a(nl_input_adpfloat_to_fixed_20U_14U_lshift_1_rg_a[4:0]),
      .s(nl_input_adpfloat_to_fixed_20U_14U_lshift_1_rg_s[3:0]),
      .z(input_adpfloat_to_fixed_20U_14U_lshift_psp_17)
    );
  ActUnit_Adpfloat2Fixed_mgc_shift_l_v5 #(.width_a(32'sd5),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd19)) input_adpfloat_to_fixed_20U_14U_lshift_2_rg (
      .a(nl_input_adpfloat_to_fixed_20U_14U_lshift_2_rg_a[4:0]),
      .s(nl_input_adpfloat_to_fixed_20U_14U_lshift_2_rg_s[3:0]),
      .z(input_adpfloat_to_fixed_20U_14U_lshift_psp_18)
    );
  ActUnit_Adpfloat2Fixed_mgc_shift_l_v5 #(.width_a(32'sd5),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd19)) input_adpfloat_to_fixed_20U_14U_lshift_3_rg (
      .a(nl_input_adpfloat_to_fixed_20U_14U_lshift_3_rg_a[4:0]),
      .s(nl_input_adpfloat_to_fixed_20U_14U_lshift_3_rg_s[3:0]),
      .z(input_adpfloat_to_fixed_20U_14U_lshift_psp_19)
    );
  ActUnit_Adpfloat2Fixed_mgc_shift_l_v5 #(.width_a(32'sd5),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd19)) input_adpfloat_to_fixed_20U_14U_lshift_4_rg (
      .a(nl_input_adpfloat_to_fixed_20U_14U_lshift_4_rg_a[4:0]),
      .s(nl_input_adpfloat_to_fixed_20U_14U_lshift_4_rg_s[3:0]),
      .z(input_adpfloat_to_fixed_20U_14U_lshift_psp_20)
    );
  ActUnit_Adpfloat2Fixed_mgc_shift_l_v5 #(.width_a(32'sd5),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd19)) input_adpfloat_to_fixed_20U_14U_lshift_5_rg (
      .a(nl_input_adpfloat_to_fixed_20U_14U_lshift_5_rg_a[4:0]),
      .s(nl_input_adpfloat_to_fixed_20U_14U_lshift_5_rg_s[3:0]),
      .z(input_adpfloat_to_fixed_20U_14U_lshift_psp_21)
    );
  ActUnit_Adpfloat2Fixed_mgc_shift_l_v5 #(.width_a(32'sd5),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd19)) input_adpfloat_to_fixed_20U_14U_lshift_6_rg (
      .a(nl_input_adpfloat_to_fixed_20U_14U_lshift_6_rg_a[4:0]),
      .s(nl_input_adpfloat_to_fixed_20U_14U_lshift_6_rg_s[3:0]),
      .z(input_adpfloat_to_fixed_20U_14U_lshift_psp_22)
    );
  ActUnit_Adpfloat2Fixed_mgc_shift_l_v5 #(.width_a(32'sd5),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd19)) input_adpfloat_to_fixed_20U_14U_lshift_7_rg (
      .a(nl_input_adpfloat_to_fixed_20U_14U_lshift_7_rg_a[4:0]),
      .s(nl_input_adpfloat_to_fixed_20U_14U_lshift_7_rg_s[3:0]),
      .z(input_adpfloat_to_fixed_20U_14U_lshift_psp_23)
    );
  ActUnit_Adpfloat2Fixed_mgc_shift_l_v5 #(.width_a(32'sd5),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd19)) input_adpfloat_to_fixed_20U_14U_lshift_8_rg (
      .a(nl_input_adpfloat_to_fixed_20U_14U_lshift_8_rg_a[4:0]),
      .s(nl_input_adpfloat_to_fixed_20U_14U_lshift_8_rg_s[3:0]),
      .z(input_adpfloat_to_fixed_20U_14U_lshift_psp_24)
    );
  ActUnit_Adpfloat2Fixed_mgc_shift_l_v5 #(.width_a(32'sd5),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd19)) input_adpfloat_to_fixed_20U_14U_lshift_9_rg (
      .a(nl_input_adpfloat_to_fixed_20U_14U_lshift_9_rg_a[4:0]),
      .s(nl_input_adpfloat_to_fixed_20U_14U_lshift_9_rg_s[3:0]),
      .z(input_adpfloat_to_fixed_20U_14U_lshift_psp_25)
    );
  ActUnit_Adpfloat2Fixed_mgc_shift_l_v5 #(.width_a(32'sd5),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd19)) input_adpfloat_to_fixed_20U_14U_lshift_10_rg (
      .a(nl_input_adpfloat_to_fixed_20U_14U_lshift_10_rg_a[4:0]),
      .s(nl_input_adpfloat_to_fixed_20U_14U_lshift_10_rg_s[3:0]),
      .z(input_adpfloat_to_fixed_20U_14U_lshift_psp_26)
    );
  ActUnit_Adpfloat2Fixed_mgc_shift_l_v5 #(.width_a(32'sd5),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd19)) input_adpfloat_to_fixed_20U_14U_lshift_11_rg (
      .a(nl_input_adpfloat_to_fixed_20U_14U_lshift_11_rg_a[4:0]),
      .s(nl_input_adpfloat_to_fixed_20U_14U_lshift_11_rg_s[3:0]),
      .z(input_adpfloat_to_fixed_20U_14U_lshift_psp_27)
    );
  ActUnit_Adpfloat2Fixed_mgc_shift_l_v5 #(.width_a(32'sd5),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd19)) input_adpfloat_to_fixed_20U_14U_lshift_12_rg (
      .a(nl_input_adpfloat_to_fixed_20U_14U_lshift_12_rg_a[4:0]),
      .s(nl_input_adpfloat_to_fixed_20U_14U_lshift_12_rg_s[3:0]),
      .z(input_adpfloat_to_fixed_20U_14U_lshift_psp_28)
    );
  ActUnit_Adpfloat2Fixed_mgc_shift_l_v5 #(.width_a(32'sd5),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd19)) input_adpfloat_to_fixed_20U_14U_lshift_13_rg (
      .a(nl_input_adpfloat_to_fixed_20U_14U_lshift_13_rg_a[4:0]),
      .s(nl_input_adpfloat_to_fixed_20U_14U_lshift_13_rg_s[3:0]),
      .z(input_adpfloat_to_fixed_20U_14U_lshift_psp_29)
    );
  ActUnit_Adpfloat2Fixed_mgc_shift_l_v5 #(.width_a(32'sd5),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd19)) input_adpfloat_to_fixed_20U_14U_lshift_14_rg (
      .a(nl_input_adpfloat_to_fixed_20U_14U_lshift_14_rg_a[4:0]),
      .s(nl_input_adpfloat_to_fixed_20U_14U_lshift_14_rg_s[3:0]),
      .z(input_adpfloat_to_fixed_20U_14U_lshift_psp_30)
    );
  ActUnit_Adpfloat2Fixed_mgc_shift_l_v5 #(.width_a(32'sd5),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd19)) input_adpfloat_to_fixed_20U_14U_lshift_15_rg (
      .a(nl_input_adpfloat_to_fixed_20U_14U_lshift_15_rg_a[4:0]),
      .s(nl_input_adpfloat_to_fixed_20U_14U_lshift_15_rg_s[3:0]),
      .z(input_adpfloat_to_fixed_20U_14U_lshift_psp_31)
    );
  assign or_15_tmp = (in_data[126:120]!=7'b0000000);
  assign or_14_tmp = (in_data[118:112]!=7'b0000000);
  assign or_13_tmp = (in_data[110:104]!=7'b0000000);
  assign or_12_tmp = (in_data[102:96]!=7'b0000000);
  assign or_11_tmp = (in_data[94:88]!=7'b0000000);
  assign or_10_tmp = (in_data[86:80]!=7'b0000000);
  assign or_9_tmp = (in_data[78:72]!=7'b0000000);
  assign or_8_tmp = (in_data[70:64]!=7'b0000000);
  assign or_7_tmp = (in_data[62:56]!=7'b0000000);
  assign or_6_tmp = (in_data[54:48]!=7'b0000000);
  assign or_5_tmp = (in_data[46:40]!=7'b0000000);
  assign or_4_tmp = (in_data[38:32]!=7'b0000000);
  assign or_3_tmp = (in_data[30:24]!=7'b0000000);
  assign or_2_tmp = (in_data[22:16]!=7'b0000000);
  assign or_1_tmp = (in_data[14:8]!=7'b0000000);
  assign or_tmp = (in_data[6:0]!=7'b0000000);
  assign input_adpfloat_to_fixed_20U_14U_if_and_ssc = (in_data[127]) & or_15_tmp;
  assign input_adpfloat_to_fixed_20U_14U_if_and_1_ssc = (in_data[119]) & or_14_tmp;
  assign input_adpfloat_to_fixed_20U_14U_if_and_2_ssc = (in_data[111]) & or_13_tmp;
  assign input_adpfloat_to_fixed_20U_14U_if_and_3_ssc = (in_data[103]) & or_12_tmp;
  assign input_adpfloat_to_fixed_20U_14U_if_and_4_ssc = (in_data[95]) & or_11_tmp;
  assign input_adpfloat_to_fixed_20U_14U_if_and_5_ssc = (in_data[87]) & or_10_tmp;
  assign input_adpfloat_to_fixed_20U_14U_if_and_6_ssc = (in_data[79]) & or_9_tmp;
  assign input_adpfloat_to_fixed_20U_14U_if_and_7_ssc = (in_data[71]) & or_8_tmp;
  assign input_adpfloat_to_fixed_20U_14U_if_and_8_ssc = (in_data[63]) & or_7_tmp;
  assign input_adpfloat_to_fixed_20U_14U_if_and_9_ssc = (in_data[55]) & or_6_tmp;
  assign input_adpfloat_to_fixed_20U_14U_if_and_10_ssc = (in_data[47]) & or_5_tmp;
  assign input_adpfloat_to_fixed_20U_14U_if_and_11_ssc = (in_data[39]) & or_4_tmp;
  assign input_adpfloat_to_fixed_20U_14U_if_and_12_ssc = (in_data[31]) & or_3_tmp;
  assign input_adpfloat_to_fixed_20U_14U_if_and_13_ssc = (in_data[23]) & or_2_tmp;
  assign input_adpfloat_to_fixed_20U_14U_if_and_14_ssc = (in_data[15]) & or_1_tmp;
  assign input_adpfloat_to_fixed_20U_14U_if_and_15_ssc = (in_data[7]) & or_tmp;
  assign nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_15_nl = (~ input_adpfloat_to_fixed_20U_14U_lshift_psp_31)
      + 19'b0000000000000000001;
  assign input_adpfloat_to_fixed_20U_14U_if_1_acc_15_nl = nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_15_nl[18:0];
  assign input_adpfloat_to_fixed_20U_14U_if_mux_nl = MUX_v_19_2_2(input_adpfloat_to_fixed_20U_14U_lshift_psp_31,
      input_adpfloat_to_fixed_20U_14U_if_1_acc_15_nl, input_adpfloat_to_fixed_20U_14U_if_and_ssc);
  assign input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_nl
      = MUX_v_20_2_2(20'b00000000000000000000, ({input_adpfloat_to_fixed_20U_14U_if_and_ssc
      , input_adpfloat_to_fixed_20U_14U_if_mux_nl}), or_15_tmp);
  assign nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_14_nl = (~ input_adpfloat_to_fixed_20U_14U_lshift_psp_30)
      + 19'b0000000000000000001;
  assign input_adpfloat_to_fixed_20U_14U_if_1_acc_14_nl = nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_14_nl[18:0];
  assign input_adpfloat_to_fixed_20U_14U_if_mux_16_nl = MUX_v_19_2_2(input_adpfloat_to_fixed_20U_14U_lshift_psp_30,
      input_adpfloat_to_fixed_20U_14U_if_1_acc_14_nl, input_adpfloat_to_fixed_20U_14U_if_and_1_ssc);
  assign input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_1_nl
      = MUX_v_20_2_2(20'b00000000000000000000, ({input_adpfloat_to_fixed_20U_14U_if_and_1_ssc
      , input_adpfloat_to_fixed_20U_14U_if_mux_16_nl}), or_14_tmp);
  assign nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_13_nl = (~ input_adpfloat_to_fixed_20U_14U_lshift_psp_29)
      + 19'b0000000000000000001;
  assign input_adpfloat_to_fixed_20U_14U_if_1_acc_13_nl = nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_13_nl[18:0];
  assign input_adpfloat_to_fixed_20U_14U_if_mux_17_nl = MUX_v_19_2_2(input_adpfloat_to_fixed_20U_14U_lshift_psp_29,
      input_adpfloat_to_fixed_20U_14U_if_1_acc_13_nl, input_adpfloat_to_fixed_20U_14U_if_and_2_ssc);
  assign input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_2_nl
      = MUX_v_20_2_2(20'b00000000000000000000, ({input_adpfloat_to_fixed_20U_14U_if_and_2_ssc
      , input_adpfloat_to_fixed_20U_14U_if_mux_17_nl}), or_13_tmp);
  assign nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_12_nl = (~ input_adpfloat_to_fixed_20U_14U_lshift_psp_28)
      + 19'b0000000000000000001;
  assign input_adpfloat_to_fixed_20U_14U_if_1_acc_12_nl = nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_12_nl[18:0];
  assign input_adpfloat_to_fixed_20U_14U_if_mux_18_nl = MUX_v_19_2_2(input_adpfloat_to_fixed_20U_14U_lshift_psp_28,
      input_adpfloat_to_fixed_20U_14U_if_1_acc_12_nl, input_adpfloat_to_fixed_20U_14U_if_and_3_ssc);
  assign input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_3_nl
      = MUX_v_20_2_2(20'b00000000000000000000, ({input_adpfloat_to_fixed_20U_14U_if_and_3_ssc
      , input_adpfloat_to_fixed_20U_14U_if_mux_18_nl}), or_12_tmp);
  assign nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_11_nl = (~ input_adpfloat_to_fixed_20U_14U_lshift_psp_27)
      + 19'b0000000000000000001;
  assign input_adpfloat_to_fixed_20U_14U_if_1_acc_11_nl = nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_11_nl[18:0];
  assign input_adpfloat_to_fixed_20U_14U_if_mux_19_nl = MUX_v_19_2_2(input_adpfloat_to_fixed_20U_14U_lshift_psp_27,
      input_adpfloat_to_fixed_20U_14U_if_1_acc_11_nl, input_adpfloat_to_fixed_20U_14U_if_and_4_ssc);
  assign input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_4_nl
      = MUX_v_20_2_2(20'b00000000000000000000, ({input_adpfloat_to_fixed_20U_14U_if_and_4_ssc
      , input_adpfloat_to_fixed_20U_14U_if_mux_19_nl}), or_11_tmp);
  assign nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_10_nl = (~ input_adpfloat_to_fixed_20U_14U_lshift_psp_26)
      + 19'b0000000000000000001;
  assign input_adpfloat_to_fixed_20U_14U_if_1_acc_10_nl = nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_10_nl[18:0];
  assign input_adpfloat_to_fixed_20U_14U_if_mux_20_nl = MUX_v_19_2_2(input_adpfloat_to_fixed_20U_14U_lshift_psp_26,
      input_adpfloat_to_fixed_20U_14U_if_1_acc_10_nl, input_adpfloat_to_fixed_20U_14U_if_and_5_ssc);
  assign input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_5_nl
      = MUX_v_20_2_2(20'b00000000000000000000, ({input_adpfloat_to_fixed_20U_14U_if_and_5_ssc
      , input_adpfloat_to_fixed_20U_14U_if_mux_20_nl}), or_10_tmp);
  assign nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_9_nl = (~ input_adpfloat_to_fixed_20U_14U_lshift_psp_25)
      + 19'b0000000000000000001;
  assign input_adpfloat_to_fixed_20U_14U_if_1_acc_9_nl = nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_9_nl[18:0];
  assign input_adpfloat_to_fixed_20U_14U_if_mux_21_nl = MUX_v_19_2_2(input_adpfloat_to_fixed_20U_14U_lshift_psp_25,
      input_adpfloat_to_fixed_20U_14U_if_1_acc_9_nl, input_adpfloat_to_fixed_20U_14U_if_and_6_ssc);
  assign input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_6_nl
      = MUX_v_20_2_2(20'b00000000000000000000, ({input_adpfloat_to_fixed_20U_14U_if_and_6_ssc
      , input_adpfloat_to_fixed_20U_14U_if_mux_21_nl}), or_9_tmp);
  assign nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_8_nl = (~ input_adpfloat_to_fixed_20U_14U_lshift_psp_24)
      + 19'b0000000000000000001;
  assign input_adpfloat_to_fixed_20U_14U_if_1_acc_8_nl = nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_8_nl[18:0];
  assign input_adpfloat_to_fixed_20U_14U_if_mux_22_nl = MUX_v_19_2_2(input_adpfloat_to_fixed_20U_14U_lshift_psp_24,
      input_adpfloat_to_fixed_20U_14U_if_1_acc_8_nl, input_adpfloat_to_fixed_20U_14U_if_and_7_ssc);
  assign input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_7_nl
      = MUX_v_20_2_2(20'b00000000000000000000, ({input_adpfloat_to_fixed_20U_14U_if_and_7_ssc
      , input_adpfloat_to_fixed_20U_14U_if_mux_22_nl}), or_8_tmp);
  assign nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_7_nl = (~ input_adpfloat_to_fixed_20U_14U_lshift_psp_23)
      + 19'b0000000000000000001;
  assign input_adpfloat_to_fixed_20U_14U_if_1_acc_7_nl = nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_7_nl[18:0];
  assign input_adpfloat_to_fixed_20U_14U_if_mux_23_nl = MUX_v_19_2_2(input_adpfloat_to_fixed_20U_14U_lshift_psp_23,
      input_adpfloat_to_fixed_20U_14U_if_1_acc_7_nl, input_adpfloat_to_fixed_20U_14U_if_and_8_ssc);
  assign input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_8_nl
      = MUX_v_20_2_2(20'b00000000000000000000, ({input_adpfloat_to_fixed_20U_14U_if_and_8_ssc
      , input_adpfloat_to_fixed_20U_14U_if_mux_23_nl}), or_7_tmp);
  assign nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_6_nl = (~ input_adpfloat_to_fixed_20U_14U_lshift_psp_22)
      + 19'b0000000000000000001;
  assign input_adpfloat_to_fixed_20U_14U_if_1_acc_6_nl = nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_6_nl[18:0];
  assign input_adpfloat_to_fixed_20U_14U_if_mux_24_nl = MUX_v_19_2_2(input_adpfloat_to_fixed_20U_14U_lshift_psp_22,
      input_adpfloat_to_fixed_20U_14U_if_1_acc_6_nl, input_adpfloat_to_fixed_20U_14U_if_and_9_ssc);
  assign input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_9_nl
      = MUX_v_20_2_2(20'b00000000000000000000, ({input_adpfloat_to_fixed_20U_14U_if_and_9_ssc
      , input_adpfloat_to_fixed_20U_14U_if_mux_24_nl}), or_6_tmp);
  assign nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_5_nl = (~ input_adpfloat_to_fixed_20U_14U_lshift_psp_21)
      + 19'b0000000000000000001;
  assign input_adpfloat_to_fixed_20U_14U_if_1_acc_5_nl = nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_5_nl[18:0];
  assign input_adpfloat_to_fixed_20U_14U_if_mux_25_nl = MUX_v_19_2_2(input_adpfloat_to_fixed_20U_14U_lshift_psp_21,
      input_adpfloat_to_fixed_20U_14U_if_1_acc_5_nl, input_adpfloat_to_fixed_20U_14U_if_and_10_ssc);
  assign input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_10_nl
      = MUX_v_20_2_2(20'b00000000000000000000, ({input_adpfloat_to_fixed_20U_14U_if_and_10_ssc
      , input_adpfloat_to_fixed_20U_14U_if_mux_25_nl}), or_5_tmp);
  assign nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_4_nl = (~ input_adpfloat_to_fixed_20U_14U_lshift_psp_20)
      + 19'b0000000000000000001;
  assign input_adpfloat_to_fixed_20U_14U_if_1_acc_4_nl = nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_4_nl[18:0];
  assign input_adpfloat_to_fixed_20U_14U_if_mux_26_nl = MUX_v_19_2_2(input_adpfloat_to_fixed_20U_14U_lshift_psp_20,
      input_adpfloat_to_fixed_20U_14U_if_1_acc_4_nl, input_adpfloat_to_fixed_20U_14U_if_and_11_ssc);
  assign input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_11_nl
      = MUX_v_20_2_2(20'b00000000000000000000, ({input_adpfloat_to_fixed_20U_14U_if_and_11_ssc
      , input_adpfloat_to_fixed_20U_14U_if_mux_26_nl}), or_4_tmp);
  assign nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_3_nl = (~ input_adpfloat_to_fixed_20U_14U_lshift_psp_19)
      + 19'b0000000000000000001;
  assign input_adpfloat_to_fixed_20U_14U_if_1_acc_3_nl = nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_3_nl[18:0];
  assign input_adpfloat_to_fixed_20U_14U_if_mux_27_nl = MUX_v_19_2_2(input_adpfloat_to_fixed_20U_14U_lshift_psp_19,
      input_adpfloat_to_fixed_20U_14U_if_1_acc_3_nl, input_adpfloat_to_fixed_20U_14U_if_and_12_ssc);
  assign input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_12_nl
      = MUX_v_20_2_2(20'b00000000000000000000, ({input_adpfloat_to_fixed_20U_14U_if_and_12_ssc
      , input_adpfloat_to_fixed_20U_14U_if_mux_27_nl}), or_3_tmp);
  assign nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_2_nl = (~ input_adpfloat_to_fixed_20U_14U_lshift_psp_18)
      + 19'b0000000000000000001;
  assign input_adpfloat_to_fixed_20U_14U_if_1_acc_2_nl = nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_2_nl[18:0];
  assign input_adpfloat_to_fixed_20U_14U_if_mux_28_nl = MUX_v_19_2_2(input_adpfloat_to_fixed_20U_14U_lshift_psp_18,
      input_adpfloat_to_fixed_20U_14U_if_1_acc_2_nl, input_adpfloat_to_fixed_20U_14U_if_and_13_ssc);
  assign input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_13_nl
      = MUX_v_20_2_2(20'b00000000000000000000, ({input_adpfloat_to_fixed_20U_14U_if_and_13_ssc
      , input_adpfloat_to_fixed_20U_14U_if_mux_28_nl}), or_2_tmp);
  assign nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_1_nl = (~ input_adpfloat_to_fixed_20U_14U_lshift_psp_17)
      + 19'b0000000000000000001;
  assign input_adpfloat_to_fixed_20U_14U_if_1_acc_1_nl = nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_1_nl[18:0];
  assign input_adpfloat_to_fixed_20U_14U_if_mux_29_nl = MUX_v_19_2_2(input_adpfloat_to_fixed_20U_14U_lshift_psp_17,
      input_adpfloat_to_fixed_20U_14U_if_1_acc_1_nl, input_adpfloat_to_fixed_20U_14U_if_and_14_ssc);
  assign input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_14_nl
      = MUX_v_20_2_2(20'b00000000000000000000, ({input_adpfloat_to_fixed_20U_14U_if_and_14_ssc
      , input_adpfloat_to_fixed_20U_14U_if_mux_29_nl}), or_1_tmp);
  assign nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_nl = (~ input_adpfloat_to_fixed_20U_14U_lshift_psp_16)
      + 19'b0000000000000000001;
  assign input_adpfloat_to_fixed_20U_14U_if_1_acc_nl = nl_input_adpfloat_to_fixed_20U_14U_if_1_acc_nl[18:0];
  assign input_adpfloat_to_fixed_20U_14U_if_mux_30_nl = MUX_v_19_2_2(input_adpfloat_to_fixed_20U_14U_lshift_psp_16,
      input_adpfloat_to_fixed_20U_14U_if_1_acc_nl, input_adpfloat_to_fixed_20U_14U_if_and_15_ssc);
  assign input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_15_nl
      = MUX_v_20_2_2(20'b00000000000000000000, ({input_adpfloat_to_fixed_20U_14U_if_and_15_ssc
      , input_adpfloat_to_fixed_20U_14U_if_mux_30_nl}), or_tmp);
  assign out_data = {input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_nl
      , input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_1_nl
      , input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_2_nl
      , input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_3_nl
      , input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_4_nl
      , input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_5_nl
      , input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_6_nl
      , input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_7_nl
      , input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_8_nl
      , input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_9_nl
      , input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_10_nl
      , input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_11_nl
      , input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_12_nl
      , input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_13_nl
      , input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_14_nl
      , input_adpfloat_to_fixed_20U_14U_if_input_adpfloat_to_fixed_20U_14U_if_and_15_nl};

  function automatic [18:0] MUX_v_19_2_2;
    input [18:0] input_0;
    input [18:0] input_1;
    input [0:0] sel;
    reg [18:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_19_2_2 = result;
  end
  endfunction


  function automatic [19:0] MUX_v_20_2_2;
    input [19:0] input_0;
    input [19:0] input_1;
    input [0:0] sel;
    reg [19:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_20_2_2 = result;
  end
  endfunction


  function automatic [3:0] conv_u2u_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_4 = {1'b0, vector};
  end
  endfunction

endmodule




//------> ./ActUnit_Fixed2Adpfloat_mgc_shift_l_beh_v5.v 
module ActUnit_Fixed2Adpfloat_mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./ActUnit_Fixed2Adpfloat_leading_sign_20_1_1_0.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   huaixil@sat8
//  Generated date: Fri Apr  8 23:11:14 2022
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    leading_sign_20_1_1_0
// ------------------------------------------------------------------


module ActUnit_Fixed2Adpfloat_leading_sign_20_1_1_0 (
  mantissa, all_same, rtn
);
  input [19:0] mantissa;
  output all_same;
  output [4:0] rtn;


  // Interconnect Declarations
  wire ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_2;
  wire ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_18_3_sdt_3;
  wire ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_26_2_sdt_2;
  wire ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_42_4_sdt_4;
  wire ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_54_5_sdt_5;
  wire ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_1;
  wire ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_14_2_sdt_1;
  wire ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_26_2_sdt_1;
  wire ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_34_2_sdt_1;
  wire ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_48_2_sdt_1;
  wire [18:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_xor_18_0;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire c_h_1_8;

  wire[0:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_and_nl;
  wire[0:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_and_1_nl;
  wire[1:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_or_1_nl;
  wire[0:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_and_74_nl;
  wire[0:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_and_76_nl;

  // Interconnect Declarations for Component Instantiations
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_xor_18_0
      = (mantissa[18:0]) ^ (signext_19_1(~ (mantissa[19])));
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_2
      = (ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_xor_18_0[16:15]==2'b11);
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_1
      = (ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_xor_18_0[18:17]==2'b11);
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_14_2_sdt_1
      = (ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_xor_18_0[14:13]==2'b11);
  assign c_h_1_2 = ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_1
      & ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_2;
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_18_3_sdt_3
      = (ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_xor_18_0[12:11]==2'b11)
      & ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_14_2_sdt_1;
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_26_2_sdt_2
      = (ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_xor_18_0[8:7]==2'b11);
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_26_2_sdt_1
      = (ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_xor_18_0[10:9]==2'b11);
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_34_2_sdt_1
      = (ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_xor_18_0[6:5]==2'b11);
  assign c_h_1_5 = ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_26_2_sdt_1
      & ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_18_3_sdt_3;
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_42_4_sdt_4
      = (ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_xor_18_0[4:3]==2'b11)
      & ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_34_2_sdt_1
      & c_h_1_5;
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_48_2_sdt_1
      = (ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_xor_18_0[2:1]==2'b11);
  assign c_h_1_8 = c_h_1_6 & ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_42_4_sdt_4;
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_54_5_sdt_5
      = (ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_xor_18_0[0])
      & ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_48_2_sdt_1
      & c_h_1_8;
  assign all_same = ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_54_5_sdt_5;
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_and_nl
      = c_h_1_6 & (~ ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_42_4_sdt_4);
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_and_1_nl
      = c_h_1_2 & (c_h_1_5 | (~ ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_18_3_sdt_3))
      & (~ c_h_1_8);
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_and_74_nl
      = ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_1
      & (ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_14_2_sdt_1
      | (~ ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_2))
      & (~((~(ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_26_2_sdt_1
      & (ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_34_2_sdt_1
      | (~ ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_26_2_sdt_2))))
      & c_h_1_6)) & (ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_48_2_sdt_1
      | (~ c_h_1_8));
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_and_76_nl
      = (ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_xor_18_0[18])
      & ((ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_xor_18_0[17:16]!=2'b10))
      & (~((~((ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_xor_18_0[14])
      & ((ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_xor_18_0[13:12]!=2'b10))))
      & c_h_1_2)) & (~((~((ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_xor_18_0[10])
      & ((ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_xor_18_0[9:8]!=2'b10))
      & (~((~((ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_xor_18_0[6])
      & ((ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_xor_18_0[5:4]!=2'b10))))
      & c_h_1_5)))) & c_h_1_6)) & (~((~((ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_xor_18_0[2:1]==2'b10)))
      & c_h_1_8));
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_or_1_nl
      = MUX_v_2_2_2(({ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_and_74_nl
      , ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_and_76_nl}),
      2'b11, ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_54_5_sdt_5);
  assign rtn = {c_h_1_8 , ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_and_nl
      , ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_and_1_nl
      , ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_if_all_sign_1_or_1_nl};

  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [18:0] signext_19_1;
    input [0:0] vector;
  begin
    signext_19_1= {{18{vector[0]}}, vector};
  end
  endfunction

endmodule




//------> ./ActUnit_Fixed2Adpfloat.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   huaixil@sat8
//  Generated date: Fri Apr  8 23:11:20 2022
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Fixed2Adpfloat
// ------------------------------------------------------------------


module ActUnit_Fixed2Adpfloat (
  in_data, out_data, adpfloat_bias
);
  input [319:0] in_data;
  output [127:0] out_data;
  input [2:0] adpfloat_bias;


  // Interconnect Declarations
  wire [6:0] ac_float_cctor_round_20_if_m_1_acc_15_tmp;
  wire [7:0] nl_ac_float_cctor_round_20_if_m_1_acc_15_tmp;
  wire [6:0] ac_float_cctor_round_20_if_m_1_acc_14_tmp;
  wire [7:0] nl_ac_float_cctor_round_20_if_m_1_acc_14_tmp;
  wire [6:0] ac_float_cctor_round_20_if_m_1_acc_13_tmp;
  wire [7:0] nl_ac_float_cctor_round_20_if_m_1_acc_13_tmp;
  wire [6:0] ac_float_cctor_round_20_if_m_1_acc_12_tmp;
  wire [7:0] nl_ac_float_cctor_round_20_if_m_1_acc_12_tmp;
  wire [6:0] ac_float_cctor_round_20_if_m_1_acc_11_tmp;
  wire [7:0] nl_ac_float_cctor_round_20_if_m_1_acc_11_tmp;
  wire [6:0] ac_float_cctor_round_20_if_m_1_acc_10_tmp;
  wire [7:0] nl_ac_float_cctor_round_20_if_m_1_acc_10_tmp;
  wire [6:0] ac_float_cctor_round_20_if_m_1_acc_9_tmp;
  wire [7:0] nl_ac_float_cctor_round_20_if_m_1_acc_9_tmp;
  wire [6:0] ac_float_cctor_round_20_if_m_1_acc_8_tmp;
  wire [7:0] nl_ac_float_cctor_round_20_if_m_1_acc_8_tmp;
  wire [6:0] ac_float_cctor_round_20_if_m_1_acc_7_tmp;
  wire [7:0] nl_ac_float_cctor_round_20_if_m_1_acc_7_tmp;
  wire [6:0] ac_float_cctor_round_20_if_m_1_acc_6_tmp;
  wire [7:0] nl_ac_float_cctor_round_20_if_m_1_acc_6_tmp;
  wire [6:0] ac_float_cctor_round_20_if_m_1_acc_5_tmp;
  wire [7:0] nl_ac_float_cctor_round_20_if_m_1_acc_5_tmp;
  wire [6:0] ac_float_cctor_round_20_if_m_1_acc_4_tmp;
  wire [7:0] nl_ac_float_cctor_round_20_if_m_1_acc_4_tmp;
  wire [6:0] ac_float_cctor_round_20_if_m_1_acc_3_tmp;
  wire [7:0] nl_ac_float_cctor_round_20_if_m_1_acc_3_tmp;
  wire [6:0] ac_float_cctor_round_20_if_m_1_acc_2_tmp;
  wire [7:0] nl_ac_float_cctor_round_20_if_m_1_acc_2_tmp;
  wire [6:0] ac_float_cctor_round_20_if_m_1_acc_1_tmp;
  wire [7:0] nl_ac_float_cctor_round_20_if_m_1_acc_1_tmp;
  wire [6:0] ac_float_cctor_round_20_if_m_1_acc_tmp;
  wire [7:0] nl_ac_float_cctor_round_20_if_m_1_acc_tmp;
  wire or_dcpl_96;
  wire or_dcpl_115;
  wire and_dcpl_20;
  wire and_dcpl_22;
  wire or_dcpl_116;
  wire or_dcpl_135;
  wire and_dcpl_43;
  wire and_dcpl_45;
  wire or_dcpl_136;
  wire or_dcpl_155;
  wire and_dcpl_66;
  wire and_dcpl_68;
  wire or_dcpl_156;
  wire or_dcpl_175;
  wire and_dcpl_89;
  wire and_dcpl_91;
  wire or_dcpl_176;
  wire or_dcpl_195;
  wire and_dcpl_112;
  wire and_dcpl_114;
  wire or_dcpl_196;
  wire or_dcpl_215;
  wire and_dcpl_135;
  wire and_dcpl_137;
  wire or_dcpl_216;
  wire or_dcpl_235;
  wire and_dcpl_158;
  wire and_dcpl_160;
  wire or_dcpl_236;
  wire or_dcpl_255;
  wire and_dcpl_181;
  wire and_dcpl_183;
  wire or_dcpl_256;
  wire or_dcpl_275;
  wire and_dcpl_204;
  wire and_dcpl_206;
  wire or_dcpl_276;
  wire or_dcpl_295;
  wire and_dcpl_227;
  wire and_dcpl_229;
  wire or_dcpl_296;
  wire or_dcpl_315;
  wire and_dcpl_250;
  wire and_dcpl_252;
  wire or_dcpl_316;
  wire or_dcpl_335;
  wire and_dcpl_273;
  wire and_dcpl_275;
  wire or_dcpl_336;
  wire or_dcpl_355;
  wire and_dcpl_296;
  wire and_dcpl_298;
  wire or_dcpl_356;
  wire or_dcpl_375;
  wire and_dcpl_319;
  wire and_dcpl_321;
  wire or_dcpl_376;
  wire or_dcpl_395;
  wire and_dcpl_342;
  wire and_dcpl_344;
  wire or_dcpl_396;
  wire or_dcpl_415;
  wire and_dcpl_365;
  wire and_dcpl_367;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_mx0;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_15_mx0;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_14_mx0;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_13_mx0;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_12_mx0;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_11_mx0;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_10_mx0;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_9_mx0;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_8_mx0;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_7_mx0;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_6_mx0;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_5_mx0;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_4_mx0;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_3_mx0;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_2_mx0;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_1_mx0;
  wire [19:0] operator_20_6_true_AC_TRN_AC_WRAP_lshift_15_itm;
  wire [19:0] operator_20_6_true_AC_TRN_AC_WRAP_lshift_14_itm;
  wire [19:0] operator_20_6_true_AC_TRN_AC_WRAP_lshift_13_itm;
  wire [19:0] operator_20_6_true_AC_TRN_AC_WRAP_lshift_12_itm;
  wire [19:0] operator_20_6_true_AC_TRN_AC_WRAP_lshift_11_itm;
  wire [19:0] operator_20_6_true_AC_TRN_AC_WRAP_lshift_10_itm;
  wire [19:0] operator_20_6_true_AC_TRN_AC_WRAP_lshift_9_itm;
  wire [19:0] operator_20_6_true_AC_TRN_AC_WRAP_lshift_8_itm;
  wire [19:0] operator_20_6_true_AC_TRN_AC_WRAP_lshift_7_itm;
  wire [19:0] operator_20_6_true_AC_TRN_AC_WRAP_lshift_6_itm;
  wire [19:0] operator_20_6_true_AC_TRN_AC_WRAP_lshift_5_itm;
  wire [19:0] operator_20_6_true_AC_TRN_AC_WRAP_lshift_4_itm;
  wire [19:0] operator_20_6_true_AC_TRN_AC_WRAP_lshift_3_itm;
  wire [19:0] operator_20_6_true_AC_TRN_AC_WRAP_lshift_2_itm;
  wire [19:0] operator_20_6_true_AC_TRN_AC_WRAP_lshift_1_itm;
  wire [19:0] operator_20_6_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_16;
  wire [6:0] nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_16;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_17;
  wire [6:0] nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_17;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_18;
  wire [6:0] nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_18;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_19;
  wire [6:0] nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_19;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_20;
  wire [6:0] nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_20;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_21;
  wire [6:0] nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_21;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_22;
  wire [6:0] nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_22;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_23;
  wire [6:0] nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_23;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_24;
  wire [6:0] nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_24;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_25;
  wire [6:0] nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_25;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_26;
  wire [6:0] nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_26;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_27;
  wire [6:0] nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_27;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_28;
  wire [6:0] nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_28;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_29;
  wire [6:0] nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_29;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_30;
  wire [6:0] nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_30;
  wire [5:0] out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_31;
  wire [6:0] nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_31;
  wire [4:0] operator_24_true_operator_24_true_conc_mx0w1_5_1;
  wire [5:0] nl_operator_24_true_operator_24_true_conc_mx0w1_5_1;
  wire [4:0] operator_24_true_operator_24_true_conc_3_mx0w1_5_1;
  wire [5:0] nl_operator_24_true_operator_24_true_conc_3_mx0w1_5_1;
  wire [4:0] operator_24_true_operator_24_true_conc_5_mx0w1_5_1;
  wire [5:0] nl_operator_24_true_operator_24_true_conc_5_mx0w1_5_1;
  wire [4:0] operator_24_true_operator_24_true_conc_7_mx0w1_5_1;
  wire [5:0] nl_operator_24_true_operator_24_true_conc_7_mx0w1_5_1;
  wire [4:0] operator_24_true_operator_24_true_conc_9_mx0w1_5_1;
  wire [5:0] nl_operator_24_true_operator_24_true_conc_9_mx0w1_5_1;
  wire [4:0] operator_24_true_operator_24_true_conc_11_mx0w1_5_1;
  wire [5:0] nl_operator_24_true_operator_24_true_conc_11_mx0w1_5_1;
  wire [4:0] operator_24_true_operator_24_true_conc_13_mx0w1_5_1;
  wire [5:0] nl_operator_24_true_operator_24_true_conc_13_mx0w1_5_1;
  wire [4:0] operator_24_true_operator_24_true_conc_15_mx0w1_5_1;
  wire [5:0] nl_operator_24_true_operator_24_true_conc_15_mx0w1_5_1;
  wire [4:0] operator_24_true_operator_24_true_conc_17_mx0w1_5_1;
  wire [5:0] nl_operator_24_true_operator_24_true_conc_17_mx0w1_5_1;
  wire [4:0] operator_24_true_operator_24_true_conc_19_mx0w1_5_1;
  wire [5:0] nl_operator_24_true_operator_24_true_conc_19_mx0w1_5_1;
  wire [4:0] operator_24_true_operator_24_true_conc_21_mx0w1_5_1;
  wire [5:0] nl_operator_24_true_operator_24_true_conc_21_mx0w1_5_1;
  wire [4:0] operator_24_true_operator_24_true_conc_23_mx0w1_5_1;
  wire [5:0] nl_operator_24_true_operator_24_true_conc_23_mx0w1_5_1;
  wire [4:0] operator_24_true_operator_24_true_conc_25_mx0w1_5_1;
  wire [5:0] nl_operator_24_true_operator_24_true_conc_25_mx0w1_5_1;
  wire [4:0] operator_24_true_operator_24_true_conc_27_mx0w1_5_1;
  wire [5:0] nl_operator_24_true_operator_24_true_conc_27_mx0w1_5_1;
  wire [4:0] operator_24_true_operator_24_true_conc_29_mx0w1_5_1;
  wire [5:0] nl_operator_24_true_operator_24_true_conc_29_mx0w1_5_1;
  wire [4:0] operator_24_true_operator_24_true_conc_31_mx0w1_5_1;
  wire [5:0] nl_operator_24_true_operator_24_true_conc_31_mx0w1_5_1;
  wire libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_32;
  wire [4:0] libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_48;
  wire libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_33;
  wire [4:0] libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_49;
  wire libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_34;
  wire [4:0] libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_50;
  wire libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_35;
  wire [4:0] libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_51;
  wire libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_36;
  wire [4:0] libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_52;
  wire libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_37;
  wire [4:0] libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_53;
  wire libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_38;
  wire [4:0] libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_54;
  wire libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_39;
  wire [4:0] libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_55;
  wire libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_40;
  wire [4:0] libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_56;
  wire libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_41;
  wire [4:0] libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_57;
  wire libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_42;
  wire [4:0] libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_58;
  wire libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_43;
  wire [4:0] libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_59;
  wire libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_44;
  wire [4:0] libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_60;
  wire libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_45;
  wire [4:0] libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_61;
  wire libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_46;
  wire [4:0] libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_62;
  wire libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_47;
  wire [4:0] libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_63;
  wire operator_23_true_acc_15_itm_2_1;
  wire operator_23_true_acc_14_itm_2_1;
  wire operator_23_true_acc_13_itm_2_1;
  wire operator_23_true_acc_12_itm_2_1;
  wire operator_23_true_acc_11_itm_2_1;
  wire operator_23_true_acc_10_itm_2_1;
  wire operator_23_true_acc_9_itm_2_1;
  wire operator_23_true_acc_8_itm_2_1;
  wire operator_23_true_acc_7_itm_2_1;
  wire operator_23_true_acc_6_itm_2_1;
  wire operator_23_true_acc_5_itm_2_1;
  wire operator_23_true_acc_4_itm_2_1;
  wire operator_23_true_acc_3_itm_2_1;
  wire operator_23_true_acc_2_itm_2_1;
  wire operator_23_true_acc_1_itm_2_1;
  wire operator_23_true_acc_itm_2_1;

  wire[0:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_nl;
  wire[2:0] x_max_lut_x_max_lut_or_nl;
  wire[2:0] x_max_lut_and_nl;
  wire[0:0] not_384_nl;
  wire[3:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_nl;
  wire[3:0] out_adpfloat_AdpfloatType_and_nl;
  wire[3:0] out_adpfloat_AdpfloatType_mux_nl;
  wire[3:0] out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_15_nl;
  wire[4:0] nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_15_nl;
  wire[0:0] out_adpfloat_AdpfloatType_and_1_nl;
  wire[0:0] not_385_nl;
  wire[0:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_1_nl;
  wire[2:0] x_max_lut_x_max_lut_or_1_nl;
  wire[2:0] x_max_lut_and_1_nl;
  wire[0:0] not_386_nl;
  wire[3:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_1_nl;
  wire[3:0] out_adpfloat_AdpfloatType_and_2_nl;
  wire[3:0] out_adpfloat_AdpfloatType_mux_16_nl;
  wire[3:0] out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_14_nl;
  wire[4:0] nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_14_nl;
  wire[0:0] out_adpfloat_AdpfloatType_and_3_nl;
  wire[0:0] not_387_nl;
  wire[0:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_2_nl;
  wire[2:0] x_max_lut_x_max_lut_or_2_nl;
  wire[2:0] x_max_lut_and_2_nl;
  wire[0:0] not_388_nl;
  wire[3:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_2_nl;
  wire[3:0] out_adpfloat_AdpfloatType_and_4_nl;
  wire[3:0] out_adpfloat_AdpfloatType_mux_17_nl;
  wire[3:0] out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_13_nl;
  wire[4:0] nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_13_nl;
  wire[0:0] out_adpfloat_AdpfloatType_and_5_nl;
  wire[0:0] not_389_nl;
  wire[0:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_3_nl;
  wire[2:0] x_max_lut_x_max_lut_or_3_nl;
  wire[2:0] x_max_lut_and_3_nl;
  wire[0:0] not_390_nl;
  wire[3:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_3_nl;
  wire[3:0] out_adpfloat_AdpfloatType_and_6_nl;
  wire[3:0] out_adpfloat_AdpfloatType_mux_18_nl;
  wire[3:0] out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_12_nl;
  wire[4:0] nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_12_nl;
  wire[0:0] out_adpfloat_AdpfloatType_and_7_nl;
  wire[0:0] not_391_nl;
  wire[0:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_4_nl;
  wire[2:0] x_max_lut_x_max_lut_or_4_nl;
  wire[2:0] x_max_lut_and_4_nl;
  wire[0:0] not_392_nl;
  wire[3:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_4_nl;
  wire[3:0] out_adpfloat_AdpfloatType_and_8_nl;
  wire[3:0] out_adpfloat_AdpfloatType_mux_19_nl;
  wire[3:0] out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_11_nl;
  wire[4:0] nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_11_nl;
  wire[0:0] out_adpfloat_AdpfloatType_and_9_nl;
  wire[0:0] not_393_nl;
  wire[0:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_5_nl;
  wire[2:0] x_max_lut_x_max_lut_or_5_nl;
  wire[2:0] x_max_lut_and_5_nl;
  wire[0:0] not_394_nl;
  wire[3:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_5_nl;
  wire[3:0] out_adpfloat_AdpfloatType_and_10_nl;
  wire[3:0] out_adpfloat_AdpfloatType_mux_20_nl;
  wire[3:0] out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_10_nl;
  wire[4:0] nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_10_nl;
  wire[0:0] out_adpfloat_AdpfloatType_and_11_nl;
  wire[0:0] not_395_nl;
  wire[0:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_6_nl;
  wire[2:0] x_max_lut_x_max_lut_or_6_nl;
  wire[2:0] x_max_lut_and_6_nl;
  wire[0:0] not_396_nl;
  wire[3:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_6_nl;
  wire[3:0] out_adpfloat_AdpfloatType_and_12_nl;
  wire[3:0] out_adpfloat_AdpfloatType_mux_21_nl;
  wire[3:0] out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_9_nl;
  wire[4:0] nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_9_nl;
  wire[0:0] out_adpfloat_AdpfloatType_and_13_nl;
  wire[0:0] not_397_nl;
  wire[0:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_7_nl;
  wire[2:0] x_max_lut_x_max_lut_or_7_nl;
  wire[2:0] x_max_lut_and_7_nl;
  wire[0:0] not_398_nl;
  wire[3:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_7_nl;
  wire[3:0] out_adpfloat_AdpfloatType_and_14_nl;
  wire[3:0] out_adpfloat_AdpfloatType_mux_22_nl;
  wire[3:0] out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_8_nl;
  wire[4:0] nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_8_nl;
  wire[0:0] out_adpfloat_AdpfloatType_and_15_nl;
  wire[0:0] not_399_nl;
  wire[0:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_8_nl;
  wire[2:0] x_max_lut_x_max_lut_or_8_nl;
  wire[2:0] x_max_lut_and_8_nl;
  wire[0:0] not_400_nl;
  wire[3:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_8_nl;
  wire[3:0] out_adpfloat_AdpfloatType_and_16_nl;
  wire[3:0] out_adpfloat_AdpfloatType_mux_23_nl;
  wire[3:0] out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_7_nl;
  wire[4:0] nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_7_nl;
  wire[0:0] out_adpfloat_AdpfloatType_and_17_nl;
  wire[0:0] not_401_nl;
  wire[0:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_9_nl;
  wire[2:0] x_max_lut_x_max_lut_or_9_nl;
  wire[2:0] x_max_lut_and_9_nl;
  wire[0:0] not_402_nl;
  wire[3:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_9_nl;
  wire[3:0] out_adpfloat_AdpfloatType_and_18_nl;
  wire[3:0] out_adpfloat_AdpfloatType_mux_24_nl;
  wire[3:0] out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_6_nl;
  wire[4:0] nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_6_nl;
  wire[0:0] out_adpfloat_AdpfloatType_and_19_nl;
  wire[0:0] not_403_nl;
  wire[0:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_10_nl;
  wire[2:0] x_max_lut_x_max_lut_or_10_nl;
  wire[2:0] x_max_lut_and_10_nl;
  wire[0:0] not_404_nl;
  wire[3:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_10_nl;
  wire[3:0] out_adpfloat_AdpfloatType_and_20_nl;
  wire[3:0] out_adpfloat_AdpfloatType_mux_25_nl;
  wire[3:0] out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_5_nl;
  wire[4:0] nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_5_nl;
  wire[0:0] out_adpfloat_AdpfloatType_and_21_nl;
  wire[0:0] not_405_nl;
  wire[0:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_11_nl;
  wire[2:0] x_max_lut_x_max_lut_or_11_nl;
  wire[2:0] x_max_lut_and_11_nl;
  wire[0:0] not_406_nl;
  wire[3:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_11_nl;
  wire[3:0] out_adpfloat_AdpfloatType_and_22_nl;
  wire[3:0] out_adpfloat_AdpfloatType_mux_26_nl;
  wire[3:0] out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_4_nl;
  wire[4:0] nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_4_nl;
  wire[0:0] out_adpfloat_AdpfloatType_and_23_nl;
  wire[0:0] not_407_nl;
  wire[0:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_12_nl;
  wire[2:0] x_max_lut_x_max_lut_or_12_nl;
  wire[2:0] x_max_lut_and_12_nl;
  wire[0:0] not_408_nl;
  wire[3:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_12_nl;
  wire[3:0] out_adpfloat_AdpfloatType_and_24_nl;
  wire[3:0] out_adpfloat_AdpfloatType_mux_27_nl;
  wire[3:0] out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_3_nl;
  wire[4:0] nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_3_nl;
  wire[0:0] out_adpfloat_AdpfloatType_and_25_nl;
  wire[0:0] not_409_nl;
  wire[0:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_13_nl;
  wire[2:0] x_max_lut_x_max_lut_or_13_nl;
  wire[2:0] x_max_lut_and_13_nl;
  wire[0:0] not_410_nl;
  wire[3:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_13_nl;
  wire[3:0] out_adpfloat_AdpfloatType_and_26_nl;
  wire[3:0] out_adpfloat_AdpfloatType_mux_28_nl;
  wire[3:0] out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_2_nl;
  wire[4:0] nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_2_nl;
  wire[0:0] out_adpfloat_AdpfloatType_and_27_nl;
  wire[0:0] not_411_nl;
  wire[0:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_14_nl;
  wire[2:0] x_max_lut_x_max_lut_or_14_nl;
  wire[2:0] x_max_lut_and_14_nl;
  wire[0:0] not_412_nl;
  wire[3:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_14_nl;
  wire[3:0] out_adpfloat_AdpfloatType_and_28_nl;
  wire[3:0] out_adpfloat_AdpfloatType_mux_29_nl;
  wire[3:0] out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_1_nl;
  wire[4:0] nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_1_nl;
  wire[0:0] out_adpfloat_AdpfloatType_and_29_nl;
  wire[0:0] not_413_nl;
  wire[0:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_15_nl;
  wire[2:0] x_max_lut_x_max_lut_or_15_nl;
  wire[2:0] x_max_lut_and_15_nl;
  wire[0:0] not_414_nl;
  wire[3:0] out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_15_nl;
  wire[3:0] out_adpfloat_AdpfloatType_and_30_nl;
  wire[3:0] out_adpfloat_AdpfloatType_mux_30_nl;
  wire[3:0] out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_nl;
  wire[4:0] nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_nl;
  wire[0:0] out_adpfloat_AdpfloatType_and_31_nl;
  wire[0:0] not_415_nl;
  wire[5:0] operator_23_true_acc_nl;
  wire[6:0] nl_operator_23_true_acc_nl;
  wire[0:0] or_5_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_15_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[0:0] ac_float_cctor_round_20_if_and_nl;
  wire[0:0] or_nl;
  wire[5:0] operator_23_true_acc_1_nl;
  wire[6:0] nl_operator_23_true_acc_1_nl;
  wire[0:0] or_11_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_14_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_1_nl;
  wire[6:0] nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_1_nl;
  wire[0:0] ac_float_cctor_round_20_if_and_1_nl;
  wire[0:0] or_6_nl;
  wire[5:0] operator_23_true_acc_2_nl;
  wire[6:0] nl_operator_23_true_acc_2_nl;
  wire[0:0] or_17_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_13_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_2_nl;
  wire[6:0] nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_2_nl;
  wire[0:0] ac_float_cctor_round_20_if_and_2_nl;
  wire[0:0] or_12_nl;
  wire[5:0] operator_23_true_acc_3_nl;
  wire[6:0] nl_operator_23_true_acc_3_nl;
  wire[0:0] or_23_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_12_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_3_nl;
  wire[6:0] nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_3_nl;
  wire[0:0] ac_float_cctor_round_20_if_and_3_nl;
  wire[0:0] or_18_nl;
  wire[5:0] operator_23_true_acc_4_nl;
  wire[6:0] nl_operator_23_true_acc_4_nl;
  wire[0:0] or_29_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_11_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_4_nl;
  wire[6:0] nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_4_nl;
  wire[0:0] ac_float_cctor_round_20_if_and_4_nl;
  wire[0:0] or_24_nl;
  wire[5:0] operator_23_true_acc_5_nl;
  wire[6:0] nl_operator_23_true_acc_5_nl;
  wire[0:0] or_35_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_10_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_5_nl;
  wire[6:0] nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_5_nl;
  wire[0:0] ac_float_cctor_round_20_if_and_5_nl;
  wire[0:0] or_30_nl;
  wire[5:0] operator_23_true_acc_6_nl;
  wire[6:0] nl_operator_23_true_acc_6_nl;
  wire[0:0] or_41_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_9_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_6_nl;
  wire[6:0] nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_6_nl;
  wire[0:0] ac_float_cctor_round_20_if_and_6_nl;
  wire[0:0] or_36_nl;
  wire[5:0] operator_23_true_acc_7_nl;
  wire[6:0] nl_operator_23_true_acc_7_nl;
  wire[0:0] or_47_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_8_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_7_nl;
  wire[6:0] nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_7_nl;
  wire[0:0] ac_float_cctor_round_20_if_and_7_nl;
  wire[0:0] or_42_nl;
  wire[5:0] operator_23_true_acc_8_nl;
  wire[6:0] nl_operator_23_true_acc_8_nl;
  wire[0:0] or_53_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_7_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_8_nl;
  wire[6:0] nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_8_nl;
  wire[0:0] ac_float_cctor_round_20_if_and_8_nl;
  wire[0:0] or_48_nl;
  wire[5:0] operator_23_true_acc_9_nl;
  wire[6:0] nl_operator_23_true_acc_9_nl;
  wire[0:0] or_59_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_6_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_9_nl;
  wire[6:0] nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_9_nl;
  wire[0:0] ac_float_cctor_round_20_if_and_9_nl;
  wire[0:0] or_54_nl;
  wire[5:0] operator_23_true_acc_10_nl;
  wire[6:0] nl_operator_23_true_acc_10_nl;
  wire[0:0] or_65_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_5_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_10_nl;
  wire[6:0] nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_10_nl;
  wire[0:0] ac_float_cctor_round_20_if_and_10_nl;
  wire[0:0] or_60_nl;
  wire[5:0] operator_23_true_acc_11_nl;
  wire[6:0] nl_operator_23_true_acc_11_nl;
  wire[0:0] or_71_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_4_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_11_nl;
  wire[6:0] nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_11_nl;
  wire[0:0] ac_float_cctor_round_20_if_and_11_nl;
  wire[0:0] or_66_nl;
  wire[5:0] operator_23_true_acc_12_nl;
  wire[6:0] nl_operator_23_true_acc_12_nl;
  wire[0:0] or_77_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_3_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_12_nl;
  wire[6:0] nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_12_nl;
  wire[0:0] ac_float_cctor_round_20_if_and_12_nl;
  wire[0:0] or_72_nl;
  wire[5:0] operator_23_true_acc_13_nl;
  wire[6:0] nl_operator_23_true_acc_13_nl;
  wire[0:0] or_83_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_2_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_13_nl;
  wire[6:0] nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_13_nl;
  wire[0:0] ac_float_cctor_round_20_if_and_13_nl;
  wire[0:0] or_78_nl;
  wire[5:0] operator_23_true_acc_14_nl;
  wire[6:0] nl_operator_23_true_acc_14_nl;
  wire[0:0] or_89_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_1_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_14_nl;
  wire[6:0] nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_14_nl;
  wire[0:0] ac_float_cctor_round_20_if_and_14_nl;
  wire[0:0] or_84_nl;
  wire[5:0] operator_23_true_acc_15_nl;
  wire[6:0] nl_operator_23_true_acc_15_nl;
  wire[0:0] or_95_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_nl;
  wire[5:0] ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_15_nl;
  wire[6:0] nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_15_nl;
  wire[0:0] ac_float_cctor_round_20_if_and_15_nl;
  wire[0:0] or_90_nl;
  wire[2:0] operator_23_true_acc_15_nl_1;
  wire[3:0] nl_operator_23_true_acc_15_nl_1;
  wire[2:0] operator_23_true_acc_14_nl_1;
  wire[3:0] nl_operator_23_true_acc_14_nl_1;
  wire[2:0] operator_23_true_acc_13_nl_1;
  wire[3:0] nl_operator_23_true_acc_13_nl_1;
  wire[2:0] operator_23_true_acc_12_nl_1;
  wire[3:0] nl_operator_23_true_acc_12_nl_1;
  wire[2:0] operator_23_true_acc_11_nl_1;
  wire[3:0] nl_operator_23_true_acc_11_nl_1;
  wire[2:0] operator_23_true_acc_10_nl_1;
  wire[3:0] nl_operator_23_true_acc_10_nl_1;
  wire[2:0] operator_23_true_acc_9_nl_1;
  wire[3:0] nl_operator_23_true_acc_9_nl_1;
  wire[2:0] operator_23_true_acc_8_nl_1;
  wire[3:0] nl_operator_23_true_acc_8_nl_1;
  wire[2:0] operator_23_true_acc_7_nl_1;
  wire[3:0] nl_operator_23_true_acc_7_nl_1;
  wire[2:0] operator_23_true_acc_6_nl_1;
  wire[3:0] nl_operator_23_true_acc_6_nl_1;
  wire[2:0] operator_23_true_acc_5_nl_1;
  wire[3:0] nl_operator_23_true_acc_5_nl_1;
  wire[2:0] operator_23_true_acc_4_nl_1;
  wire[3:0] nl_operator_23_true_acc_4_nl_1;
  wire[2:0] operator_23_true_acc_3_nl_1;
  wire[3:0] nl_operator_23_true_acc_3_nl_1;
  wire[2:0] operator_23_true_acc_2_nl_1;
  wire[3:0] nl_operator_23_true_acc_2_nl_1;
  wire[2:0] operator_23_true_acc_1_nl_1;
  wire[3:0] nl_operator_23_true_acc_1_nl_1;
  wire[2:0] operator_23_true_acc_nl_1;
  wire[3:0] nl_operator_23_true_acc_nl_1;

  // Interconnect Declarations for Component Instantiations
  wire [19:0] nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_15_rg_a;
  assign nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_15_rg_a = in_data[319:300];
  wire [19:0] nl_leading_sign_20_1_1_0_15_rg_mantissa;
  assign nl_leading_sign_20_1_1_0_15_rg_mantissa = in_data[319:300];
  wire [19:0] nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_14_rg_a;
  assign nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_14_rg_a = in_data[299:280];
  wire [19:0] nl_leading_sign_20_1_1_0_14_rg_mantissa;
  assign nl_leading_sign_20_1_1_0_14_rg_mantissa = in_data[299:280];
  wire [19:0] nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_13_rg_a;
  assign nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_13_rg_a = in_data[279:260];
  wire [19:0] nl_leading_sign_20_1_1_0_13_rg_mantissa;
  assign nl_leading_sign_20_1_1_0_13_rg_mantissa = in_data[279:260];
  wire [19:0] nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_12_rg_a;
  assign nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_12_rg_a = in_data[259:240];
  wire [19:0] nl_leading_sign_20_1_1_0_12_rg_mantissa;
  assign nl_leading_sign_20_1_1_0_12_rg_mantissa = in_data[259:240];
  wire [19:0] nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_11_rg_a;
  assign nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_11_rg_a = in_data[239:220];
  wire [19:0] nl_leading_sign_20_1_1_0_11_rg_mantissa;
  assign nl_leading_sign_20_1_1_0_11_rg_mantissa = in_data[239:220];
  wire [19:0] nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_10_rg_a;
  assign nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_10_rg_a = in_data[219:200];
  wire [19:0] nl_leading_sign_20_1_1_0_10_rg_mantissa;
  assign nl_leading_sign_20_1_1_0_10_rg_mantissa = in_data[219:200];
  wire [19:0] nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_9_rg_a;
  assign nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_9_rg_a = in_data[199:180];
  wire [19:0] nl_leading_sign_20_1_1_0_9_rg_mantissa;
  assign nl_leading_sign_20_1_1_0_9_rg_mantissa = in_data[199:180];
  wire [19:0] nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_8_rg_a;
  assign nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_8_rg_a = in_data[179:160];
  wire [19:0] nl_leading_sign_20_1_1_0_8_rg_mantissa;
  assign nl_leading_sign_20_1_1_0_8_rg_mantissa = in_data[179:160];
  wire [19:0] nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_7_rg_a;
  assign nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_7_rg_a = in_data[159:140];
  wire [19:0] nl_leading_sign_20_1_1_0_7_rg_mantissa;
  assign nl_leading_sign_20_1_1_0_7_rg_mantissa = in_data[159:140];
  wire [19:0] nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_6_rg_a;
  assign nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_6_rg_a = in_data[139:120];
  wire [19:0] nl_leading_sign_20_1_1_0_6_rg_mantissa;
  assign nl_leading_sign_20_1_1_0_6_rg_mantissa = in_data[139:120];
  wire [19:0] nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_5_rg_a;
  assign nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_5_rg_a = in_data[119:100];
  wire [19:0] nl_leading_sign_20_1_1_0_5_rg_mantissa;
  assign nl_leading_sign_20_1_1_0_5_rg_mantissa = in_data[119:100];
  wire [19:0] nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_4_rg_a;
  assign nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_4_rg_a = in_data[99:80];
  wire [19:0] nl_leading_sign_20_1_1_0_4_rg_mantissa;
  assign nl_leading_sign_20_1_1_0_4_rg_mantissa = in_data[99:80];
  wire [19:0] nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_3_rg_a;
  assign nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_3_rg_a = in_data[79:60];
  wire [19:0] nl_leading_sign_20_1_1_0_3_rg_mantissa;
  assign nl_leading_sign_20_1_1_0_3_rg_mantissa = in_data[79:60];
  wire [19:0] nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_2_rg_a;
  assign nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_2_rg_a = in_data[59:40];
  wire [19:0] nl_leading_sign_20_1_1_0_2_rg_mantissa;
  assign nl_leading_sign_20_1_1_0_2_rg_mantissa = in_data[59:40];
  wire [19:0] nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_1_rg_a;
  assign nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_1_rg_a = in_data[39:20];
  wire [19:0] nl_leading_sign_20_1_1_0_1_rg_mantissa;
  assign nl_leading_sign_20_1_1_0_1_rg_mantissa = in_data[39:20];
  wire [19:0] nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_rg_a = in_data[19:0];
  wire [19:0] nl_leading_sign_20_1_1_0_rg_mantissa;
  assign nl_leading_sign_20_1_1_0_rg_mantissa = in_data[19:0];
  ActUnit_Fixed2Adpfloat_mgc_shift_l_v5 #(.width_a(32'sd20),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd20)) operator_20_6_true_AC_TRN_AC_WRAP_lshift_15_rg (
      .a(nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_15_rg_a[19:0]),
      .s(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_48),
      .z(operator_20_6_true_AC_TRN_AC_WRAP_lshift_15_itm)
    );
  ActUnit_Fixed2Adpfloat_leading_sign_20_1_1_0  leading_sign_20_1_1_0_15_rg (
      .mantissa(nl_leading_sign_20_1_1_0_15_rg_mantissa[19:0]),
      .all_same(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_32),
      .rtn(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_48)
    );
  ActUnit_Fixed2Adpfloat_mgc_shift_l_v5 #(.width_a(32'sd20),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd20)) operator_20_6_true_AC_TRN_AC_WRAP_lshift_14_rg (
      .a(nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_14_rg_a[19:0]),
      .s(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_49),
      .z(operator_20_6_true_AC_TRN_AC_WRAP_lshift_14_itm)
    );
  ActUnit_Fixed2Adpfloat_leading_sign_20_1_1_0  leading_sign_20_1_1_0_14_rg (
      .mantissa(nl_leading_sign_20_1_1_0_14_rg_mantissa[19:0]),
      .all_same(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_33),
      .rtn(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_49)
    );
  ActUnit_Fixed2Adpfloat_mgc_shift_l_v5 #(.width_a(32'sd20),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd20)) operator_20_6_true_AC_TRN_AC_WRAP_lshift_13_rg (
      .a(nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_13_rg_a[19:0]),
      .s(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_50),
      .z(operator_20_6_true_AC_TRN_AC_WRAP_lshift_13_itm)
    );
  ActUnit_Fixed2Adpfloat_leading_sign_20_1_1_0  leading_sign_20_1_1_0_13_rg (
      .mantissa(nl_leading_sign_20_1_1_0_13_rg_mantissa[19:0]),
      .all_same(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_34),
      .rtn(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_50)
    );
  ActUnit_Fixed2Adpfloat_mgc_shift_l_v5 #(.width_a(32'sd20),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd20)) operator_20_6_true_AC_TRN_AC_WRAP_lshift_12_rg (
      .a(nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_12_rg_a[19:0]),
      .s(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_51),
      .z(operator_20_6_true_AC_TRN_AC_WRAP_lshift_12_itm)
    );
  ActUnit_Fixed2Adpfloat_leading_sign_20_1_1_0  leading_sign_20_1_1_0_12_rg (
      .mantissa(nl_leading_sign_20_1_1_0_12_rg_mantissa[19:0]),
      .all_same(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_35),
      .rtn(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_51)
    );
  ActUnit_Fixed2Adpfloat_mgc_shift_l_v5 #(.width_a(32'sd20),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd20)) operator_20_6_true_AC_TRN_AC_WRAP_lshift_11_rg (
      .a(nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_11_rg_a[19:0]),
      .s(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_52),
      .z(operator_20_6_true_AC_TRN_AC_WRAP_lshift_11_itm)
    );
  ActUnit_Fixed2Adpfloat_leading_sign_20_1_1_0  leading_sign_20_1_1_0_11_rg (
      .mantissa(nl_leading_sign_20_1_1_0_11_rg_mantissa[19:0]),
      .all_same(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_36),
      .rtn(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_52)
    );
  ActUnit_Fixed2Adpfloat_mgc_shift_l_v5 #(.width_a(32'sd20),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd20)) operator_20_6_true_AC_TRN_AC_WRAP_lshift_10_rg (
      .a(nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_10_rg_a[19:0]),
      .s(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_53),
      .z(operator_20_6_true_AC_TRN_AC_WRAP_lshift_10_itm)
    );
  ActUnit_Fixed2Adpfloat_leading_sign_20_1_1_0  leading_sign_20_1_1_0_10_rg (
      .mantissa(nl_leading_sign_20_1_1_0_10_rg_mantissa[19:0]),
      .all_same(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_37),
      .rtn(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_53)
    );
  ActUnit_Fixed2Adpfloat_mgc_shift_l_v5 #(.width_a(32'sd20),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd20)) operator_20_6_true_AC_TRN_AC_WRAP_lshift_9_rg (
      .a(nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_9_rg_a[19:0]),
      .s(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_54),
      .z(operator_20_6_true_AC_TRN_AC_WRAP_lshift_9_itm)
    );
  ActUnit_Fixed2Adpfloat_leading_sign_20_1_1_0  leading_sign_20_1_1_0_9_rg (
      .mantissa(nl_leading_sign_20_1_1_0_9_rg_mantissa[19:0]),
      .all_same(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_38),
      .rtn(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_54)
    );
  ActUnit_Fixed2Adpfloat_mgc_shift_l_v5 #(.width_a(32'sd20),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd20)) operator_20_6_true_AC_TRN_AC_WRAP_lshift_8_rg (
      .a(nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_8_rg_a[19:0]),
      .s(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_55),
      .z(operator_20_6_true_AC_TRN_AC_WRAP_lshift_8_itm)
    );
  ActUnit_Fixed2Adpfloat_leading_sign_20_1_1_0  leading_sign_20_1_1_0_8_rg (
      .mantissa(nl_leading_sign_20_1_1_0_8_rg_mantissa[19:0]),
      .all_same(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_39),
      .rtn(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_55)
    );
  ActUnit_Fixed2Adpfloat_mgc_shift_l_v5 #(.width_a(32'sd20),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd20)) operator_20_6_true_AC_TRN_AC_WRAP_lshift_7_rg (
      .a(nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_7_rg_a[19:0]),
      .s(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_56),
      .z(operator_20_6_true_AC_TRN_AC_WRAP_lshift_7_itm)
    );
  ActUnit_Fixed2Adpfloat_leading_sign_20_1_1_0  leading_sign_20_1_1_0_7_rg (
      .mantissa(nl_leading_sign_20_1_1_0_7_rg_mantissa[19:0]),
      .all_same(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_40),
      .rtn(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_56)
    );
  ActUnit_Fixed2Adpfloat_mgc_shift_l_v5 #(.width_a(32'sd20),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd20)) operator_20_6_true_AC_TRN_AC_WRAP_lshift_6_rg (
      .a(nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_6_rg_a[19:0]),
      .s(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_57),
      .z(operator_20_6_true_AC_TRN_AC_WRAP_lshift_6_itm)
    );
  ActUnit_Fixed2Adpfloat_leading_sign_20_1_1_0  leading_sign_20_1_1_0_6_rg (
      .mantissa(nl_leading_sign_20_1_1_0_6_rg_mantissa[19:0]),
      .all_same(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_41),
      .rtn(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_57)
    );
  ActUnit_Fixed2Adpfloat_mgc_shift_l_v5 #(.width_a(32'sd20),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd20)) operator_20_6_true_AC_TRN_AC_WRAP_lshift_5_rg (
      .a(nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_5_rg_a[19:0]),
      .s(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_58),
      .z(operator_20_6_true_AC_TRN_AC_WRAP_lshift_5_itm)
    );
  ActUnit_Fixed2Adpfloat_leading_sign_20_1_1_0  leading_sign_20_1_1_0_5_rg (
      .mantissa(nl_leading_sign_20_1_1_0_5_rg_mantissa[19:0]),
      .all_same(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_42),
      .rtn(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_58)
    );
  ActUnit_Fixed2Adpfloat_mgc_shift_l_v5 #(.width_a(32'sd20),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd20)) operator_20_6_true_AC_TRN_AC_WRAP_lshift_4_rg (
      .a(nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_4_rg_a[19:0]),
      .s(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_59),
      .z(operator_20_6_true_AC_TRN_AC_WRAP_lshift_4_itm)
    );
  ActUnit_Fixed2Adpfloat_leading_sign_20_1_1_0  leading_sign_20_1_1_0_4_rg (
      .mantissa(nl_leading_sign_20_1_1_0_4_rg_mantissa[19:0]),
      .all_same(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_43),
      .rtn(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_59)
    );
  ActUnit_Fixed2Adpfloat_mgc_shift_l_v5 #(.width_a(32'sd20),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd20)) operator_20_6_true_AC_TRN_AC_WRAP_lshift_3_rg (
      .a(nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_3_rg_a[19:0]),
      .s(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_60),
      .z(operator_20_6_true_AC_TRN_AC_WRAP_lshift_3_itm)
    );
  ActUnit_Fixed2Adpfloat_leading_sign_20_1_1_0  leading_sign_20_1_1_0_3_rg (
      .mantissa(nl_leading_sign_20_1_1_0_3_rg_mantissa[19:0]),
      .all_same(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_44),
      .rtn(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_60)
    );
  ActUnit_Fixed2Adpfloat_mgc_shift_l_v5 #(.width_a(32'sd20),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd20)) operator_20_6_true_AC_TRN_AC_WRAP_lshift_2_rg (
      .a(nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_2_rg_a[19:0]),
      .s(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_61),
      .z(operator_20_6_true_AC_TRN_AC_WRAP_lshift_2_itm)
    );
  ActUnit_Fixed2Adpfloat_leading_sign_20_1_1_0  leading_sign_20_1_1_0_2_rg (
      .mantissa(nl_leading_sign_20_1_1_0_2_rg_mantissa[19:0]),
      .all_same(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_45),
      .rtn(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_61)
    );
  ActUnit_Fixed2Adpfloat_mgc_shift_l_v5 #(.width_a(32'sd20),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd20)) operator_20_6_true_AC_TRN_AC_WRAP_lshift_1_rg (
      .a(nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_1_rg_a[19:0]),
      .s(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_62),
      .z(operator_20_6_true_AC_TRN_AC_WRAP_lshift_1_itm)
    );
  ActUnit_Fixed2Adpfloat_leading_sign_20_1_1_0  leading_sign_20_1_1_0_1_rg (
      .mantissa(nl_leading_sign_20_1_1_0_1_rg_mantissa[19:0]),
      .all_same(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_46),
      .rtn(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_62)
    );
  ActUnit_Fixed2Adpfloat_mgc_shift_l_v5 #(.width_a(32'sd20),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd20)) operator_20_6_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_operator_20_6_true_AC_TRN_AC_WRAP_lshift_rg_a[19:0]),
      .s(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_63),
      .z(operator_20_6_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  ActUnit_Fixed2Adpfloat_leading_sign_20_1_1_0  leading_sign_20_1_1_0_rg (
      .mantissa(nl_leading_sign_20_1_1_0_rg_mantissa[19:0]),
      .all_same(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_47),
      .rtn(libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_63)
    );
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_nl = (ac_float_cctor_round_20_if_m_1_acc_15_tmp[6])
      & and_dcpl_367;
  assign not_384_nl = ~ or_dcpl_396;
  assign x_max_lut_and_nl = MUX_v_3_2_2(3'b000, (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_mx0[2:0]),
      not_384_nl);
  assign x_max_lut_x_max_lut_or_nl = MUX_v_3_2_2(x_max_lut_and_nl, 3'b111, and_dcpl_365);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_15_nl =  -(ac_float_cctor_round_20_if_m_1_acc_15_tmp[3:0]);
  assign out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_15_nl = nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_15_nl[3:0];
  assign out_adpfloat_AdpfloatType_and_1_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_15_tmp[6]))
      & and_dcpl_367;
  assign out_adpfloat_AdpfloatType_mux_nl = MUX_v_4_2_2(out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_15_nl,
      (ac_float_cctor_round_20_if_m_1_acc_15_tmp[3:0]), out_adpfloat_AdpfloatType_and_1_nl);
  assign not_385_nl = ~ or_dcpl_396;
  assign out_adpfloat_AdpfloatType_and_nl = MUX_v_4_2_2(4'b0000, out_adpfloat_AdpfloatType_mux_nl,
      not_385_nl);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_nl = MUX_v_4_2_2(out_adpfloat_AdpfloatType_and_nl,
      4'b1111, and_dcpl_365);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_1_nl = (ac_float_cctor_round_20_if_m_1_acc_14_tmp[6])
      & and_dcpl_344;
  assign not_386_nl = ~ or_dcpl_376;
  assign x_max_lut_and_1_nl = MUX_v_3_2_2(3'b000, (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_15_mx0[2:0]),
      not_386_nl);
  assign x_max_lut_x_max_lut_or_1_nl = MUX_v_3_2_2(x_max_lut_and_1_nl, 3'b111, and_dcpl_342);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_14_nl =  -(ac_float_cctor_round_20_if_m_1_acc_14_tmp[3:0]);
  assign out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_14_nl = nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_14_nl[3:0];
  assign out_adpfloat_AdpfloatType_and_3_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_14_tmp[6]))
      & and_dcpl_344;
  assign out_adpfloat_AdpfloatType_mux_16_nl = MUX_v_4_2_2(out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_14_nl,
      (ac_float_cctor_round_20_if_m_1_acc_14_tmp[3:0]), out_adpfloat_AdpfloatType_and_3_nl);
  assign not_387_nl = ~ or_dcpl_376;
  assign out_adpfloat_AdpfloatType_and_2_nl = MUX_v_4_2_2(4'b0000, out_adpfloat_AdpfloatType_mux_16_nl,
      not_387_nl);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_1_nl = MUX_v_4_2_2(out_adpfloat_AdpfloatType_and_2_nl,
      4'b1111, and_dcpl_342);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_2_nl = (ac_float_cctor_round_20_if_m_1_acc_13_tmp[6])
      & and_dcpl_321;
  assign not_388_nl = ~ or_dcpl_356;
  assign x_max_lut_and_2_nl = MUX_v_3_2_2(3'b000, (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_14_mx0[2:0]),
      not_388_nl);
  assign x_max_lut_x_max_lut_or_2_nl = MUX_v_3_2_2(x_max_lut_and_2_nl, 3'b111, and_dcpl_319);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_13_nl =  -(ac_float_cctor_round_20_if_m_1_acc_13_tmp[3:0]);
  assign out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_13_nl = nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_13_nl[3:0];
  assign out_adpfloat_AdpfloatType_and_5_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_13_tmp[6]))
      & and_dcpl_321;
  assign out_adpfloat_AdpfloatType_mux_17_nl = MUX_v_4_2_2(out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_13_nl,
      (ac_float_cctor_round_20_if_m_1_acc_13_tmp[3:0]), out_adpfloat_AdpfloatType_and_5_nl);
  assign not_389_nl = ~ or_dcpl_356;
  assign out_adpfloat_AdpfloatType_and_4_nl = MUX_v_4_2_2(4'b0000, out_adpfloat_AdpfloatType_mux_17_nl,
      not_389_nl);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_2_nl = MUX_v_4_2_2(out_adpfloat_AdpfloatType_and_4_nl,
      4'b1111, and_dcpl_319);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_3_nl = (ac_float_cctor_round_20_if_m_1_acc_12_tmp[6])
      & and_dcpl_298;
  assign not_390_nl = ~ or_dcpl_336;
  assign x_max_lut_and_3_nl = MUX_v_3_2_2(3'b000, (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_13_mx0[2:0]),
      not_390_nl);
  assign x_max_lut_x_max_lut_or_3_nl = MUX_v_3_2_2(x_max_lut_and_3_nl, 3'b111, and_dcpl_296);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_12_nl =  -(ac_float_cctor_round_20_if_m_1_acc_12_tmp[3:0]);
  assign out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_12_nl = nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_12_nl[3:0];
  assign out_adpfloat_AdpfloatType_and_7_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_12_tmp[6]))
      & and_dcpl_298;
  assign out_adpfloat_AdpfloatType_mux_18_nl = MUX_v_4_2_2(out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_12_nl,
      (ac_float_cctor_round_20_if_m_1_acc_12_tmp[3:0]), out_adpfloat_AdpfloatType_and_7_nl);
  assign not_391_nl = ~ or_dcpl_336;
  assign out_adpfloat_AdpfloatType_and_6_nl = MUX_v_4_2_2(4'b0000, out_adpfloat_AdpfloatType_mux_18_nl,
      not_391_nl);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_3_nl = MUX_v_4_2_2(out_adpfloat_AdpfloatType_and_6_nl,
      4'b1111, and_dcpl_296);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_4_nl = (ac_float_cctor_round_20_if_m_1_acc_11_tmp[6])
      & and_dcpl_275;
  assign not_392_nl = ~ or_dcpl_316;
  assign x_max_lut_and_4_nl = MUX_v_3_2_2(3'b000, (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_12_mx0[2:0]),
      not_392_nl);
  assign x_max_lut_x_max_lut_or_4_nl = MUX_v_3_2_2(x_max_lut_and_4_nl, 3'b111, and_dcpl_273);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_11_nl =  -(ac_float_cctor_round_20_if_m_1_acc_11_tmp[3:0]);
  assign out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_11_nl = nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_11_nl[3:0];
  assign out_adpfloat_AdpfloatType_and_9_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_11_tmp[6]))
      & and_dcpl_275;
  assign out_adpfloat_AdpfloatType_mux_19_nl = MUX_v_4_2_2(out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_11_nl,
      (ac_float_cctor_round_20_if_m_1_acc_11_tmp[3:0]), out_adpfloat_AdpfloatType_and_9_nl);
  assign not_393_nl = ~ or_dcpl_316;
  assign out_adpfloat_AdpfloatType_and_8_nl = MUX_v_4_2_2(4'b0000, out_adpfloat_AdpfloatType_mux_19_nl,
      not_393_nl);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_4_nl = MUX_v_4_2_2(out_adpfloat_AdpfloatType_and_8_nl,
      4'b1111, and_dcpl_273);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_5_nl = (ac_float_cctor_round_20_if_m_1_acc_10_tmp[6])
      & and_dcpl_252;
  assign not_394_nl = ~ or_dcpl_296;
  assign x_max_lut_and_5_nl = MUX_v_3_2_2(3'b000, (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_11_mx0[2:0]),
      not_394_nl);
  assign x_max_lut_x_max_lut_or_5_nl = MUX_v_3_2_2(x_max_lut_and_5_nl, 3'b111, and_dcpl_250);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_10_nl =  -(ac_float_cctor_round_20_if_m_1_acc_10_tmp[3:0]);
  assign out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_10_nl = nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_10_nl[3:0];
  assign out_adpfloat_AdpfloatType_and_11_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_10_tmp[6]))
      & and_dcpl_252;
  assign out_adpfloat_AdpfloatType_mux_20_nl = MUX_v_4_2_2(out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_10_nl,
      (ac_float_cctor_round_20_if_m_1_acc_10_tmp[3:0]), out_adpfloat_AdpfloatType_and_11_nl);
  assign not_395_nl = ~ or_dcpl_296;
  assign out_adpfloat_AdpfloatType_and_10_nl = MUX_v_4_2_2(4'b0000, out_adpfloat_AdpfloatType_mux_20_nl,
      not_395_nl);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_5_nl = MUX_v_4_2_2(out_adpfloat_AdpfloatType_and_10_nl,
      4'b1111, and_dcpl_250);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_6_nl = (ac_float_cctor_round_20_if_m_1_acc_9_tmp[6])
      & and_dcpl_229;
  assign not_396_nl = ~ or_dcpl_276;
  assign x_max_lut_and_6_nl = MUX_v_3_2_2(3'b000, (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_10_mx0[2:0]),
      not_396_nl);
  assign x_max_lut_x_max_lut_or_6_nl = MUX_v_3_2_2(x_max_lut_and_6_nl, 3'b111, and_dcpl_227);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_9_nl =  -(ac_float_cctor_round_20_if_m_1_acc_9_tmp[3:0]);
  assign out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_9_nl = nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_9_nl[3:0];
  assign out_adpfloat_AdpfloatType_and_13_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_9_tmp[6]))
      & and_dcpl_229;
  assign out_adpfloat_AdpfloatType_mux_21_nl = MUX_v_4_2_2(out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_9_nl,
      (ac_float_cctor_round_20_if_m_1_acc_9_tmp[3:0]), out_adpfloat_AdpfloatType_and_13_nl);
  assign not_397_nl = ~ or_dcpl_276;
  assign out_adpfloat_AdpfloatType_and_12_nl = MUX_v_4_2_2(4'b0000, out_adpfloat_AdpfloatType_mux_21_nl,
      not_397_nl);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_6_nl = MUX_v_4_2_2(out_adpfloat_AdpfloatType_and_12_nl,
      4'b1111, and_dcpl_227);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_7_nl = (ac_float_cctor_round_20_if_m_1_acc_8_tmp[6])
      & and_dcpl_206;
  assign not_398_nl = ~ or_dcpl_256;
  assign x_max_lut_and_7_nl = MUX_v_3_2_2(3'b000, (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_9_mx0[2:0]),
      not_398_nl);
  assign x_max_lut_x_max_lut_or_7_nl = MUX_v_3_2_2(x_max_lut_and_7_nl, 3'b111, and_dcpl_204);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_8_nl =  -(ac_float_cctor_round_20_if_m_1_acc_8_tmp[3:0]);
  assign out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_8_nl = nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_8_nl[3:0];
  assign out_adpfloat_AdpfloatType_and_15_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_8_tmp[6]))
      & and_dcpl_206;
  assign out_adpfloat_AdpfloatType_mux_22_nl = MUX_v_4_2_2(out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_8_nl,
      (ac_float_cctor_round_20_if_m_1_acc_8_tmp[3:0]), out_adpfloat_AdpfloatType_and_15_nl);
  assign not_399_nl = ~ or_dcpl_256;
  assign out_adpfloat_AdpfloatType_and_14_nl = MUX_v_4_2_2(4'b0000, out_adpfloat_AdpfloatType_mux_22_nl,
      not_399_nl);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_7_nl = MUX_v_4_2_2(out_adpfloat_AdpfloatType_and_14_nl,
      4'b1111, and_dcpl_204);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_8_nl = (ac_float_cctor_round_20_if_m_1_acc_7_tmp[6])
      & and_dcpl_183;
  assign not_400_nl = ~ or_dcpl_236;
  assign x_max_lut_and_8_nl = MUX_v_3_2_2(3'b000, (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_8_mx0[2:0]),
      not_400_nl);
  assign x_max_lut_x_max_lut_or_8_nl = MUX_v_3_2_2(x_max_lut_and_8_nl, 3'b111, and_dcpl_181);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_7_nl =  -(ac_float_cctor_round_20_if_m_1_acc_7_tmp[3:0]);
  assign out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_7_nl = nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_7_nl[3:0];
  assign out_adpfloat_AdpfloatType_and_17_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_7_tmp[6]))
      & and_dcpl_183;
  assign out_adpfloat_AdpfloatType_mux_23_nl = MUX_v_4_2_2(out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_7_nl,
      (ac_float_cctor_round_20_if_m_1_acc_7_tmp[3:0]), out_adpfloat_AdpfloatType_and_17_nl);
  assign not_401_nl = ~ or_dcpl_236;
  assign out_adpfloat_AdpfloatType_and_16_nl = MUX_v_4_2_2(4'b0000, out_adpfloat_AdpfloatType_mux_23_nl,
      not_401_nl);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_8_nl = MUX_v_4_2_2(out_adpfloat_AdpfloatType_and_16_nl,
      4'b1111, and_dcpl_181);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_9_nl = (ac_float_cctor_round_20_if_m_1_acc_6_tmp[6])
      & and_dcpl_160;
  assign not_402_nl = ~ or_dcpl_216;
  assign x_max_lut_and_9_nl = MUX_v_3_2_2(3'b000, (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_7_mx0[2:0]),
      not_402_nl);
  assign x_max_lut_x_max_lut_or_9_nl = MUX_v_3_2_2(x_max_lut_and_9_nl, 3'b111, and_dcpl_158);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_6_nl =  -(ac_float_cctor_round_20_if_m_1_acc_6_tmp[3:0]);
  assign out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_6_nl = nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_6_nl[3:0];
  assign out_adpfloat_AdpfloatType_and_19_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_6_tmp[6]))
      & and_dcpl_160;
  assign out_adpfloat_AdpfloatType_mux_24_nl = MUX_v_4_2_2(out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_6_nl,
      (ac_float_cctor_round_20_if_m_1_acc_6_tmp[3:0]), out_adpfloat_AdpfloatType_and_19_nl);
  assign not_403_nl = ~ or_dcpl_216;
  assign out_adpfloat_AdpfloatType_and_18_nl = MUX_v_4_2_2(4'b0000, out_adpfloat_AdpfloatType_mux_24_nl,
      not_403_nl);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_9_nl = MUX_v_4_2_2(out_adpfloat_AdpfloatType_and_18_nl,
      4'b1111, and_dcpl_158);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_10_nl = (ac_float_cctor_round_20_if_m_1_acc_5_tmp[6])
      & and_dcpl_137;
  assign not_404_nl = ~ or_dcpl_196;
  assign x_max_lut_and_10_nl = MUX_v_3_2_2(3'b000, (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_6_mx0[2:0]),
      not_404_nl);
  assign x_max_lut_x_max_lut_or_10_nl = MUX_v_3_2_2(x_max_lut_and_10_nl, 3'b111,
      and_dcpl_135);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_5_nl =  -(ac_float_cctor_round_20_if_m_1_acc_5_tmp[3:0]);
  assign out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_5_nl = nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_5_nl[3:0];
  assign out_adpfloat_AdpfloatType_and_21_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_5_tmp[6]))
      & and_dcpl_137;
  assign out_adpfloat_AdpfloatType_mux_25_nl = MUX_v_4_2_2(out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_5_nl,
      (ac_float_cctor_round_20_if_m_1_acc_5_tmp[3:0]), out_adpfloat_AdpfloatType_and_21_nl);
  assign not_405_nl = ~ or_dcpl_196;
  assign out_adpfloat_AdpfloatType_and_20_nl = MUX_v_4_2_2(4'b0000, out_adpfloat_AdpfloatType_mux_25_nl,
      not_405_nl);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_10_nl = MUX_v_4_2_2(out_adpfloat_AdpfloatType_and_20_nl,
      4'b1111, and_dcpl_135);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_11_nl = (ac_float_cctor_round_20_if_m_1_acc_4_tmp[6])
      & and_dcpl_114;
  assign not_406_nl = ~ or_dcpl_176;
  assign x_max_lut_and_11_nl = MUX_v_3_2_2(3'b000, (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_5_mx0[2:0]),
      not_406_nl);
  assign x_max_lut_x_max_lut_or_11_nl = MUX_v_3_2_2(x_max_lut_and_11_nl, 3'b111,
      and_dcpl_112);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_4_nl =  -(ac_float_cctor_round_20_if_m_1_acc_4_tmp[3:0]);
  assign out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_4_nl = nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_4_nl[3:0];
  assign out_adpfloat_AdpfloatType_and_23_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_4_tmp[6]))
      & and_dcpl_114;
  assign out_adpfloat_AdpfloatType_mux_26_nl = MUX_v_4_2_2(out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_4_nl,
      (ac_float_cctor_round_20_if_m_1_acc_4_tmp[3:0]), out_adpfloat_AdpfloatType_and_23_nl);
  assign not_407_nl = ~ or_dcpl_176;
  assign out_adpfloat_AdpfloatType_and_22_nl = MUX_v_4_2_2(4'b0000, out_adpfloat_AdpfloatType_mux_26_nl,
      not_407_nl);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_11_nl = MUX_v_4_2_2(out_adpfloat_AdpfloatType_and_22_nl,
      4'b1111, and_dcpl_112);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_12_nl = (ac_float_cctor_round_20_if_m_1_acc_3_tmp[6])
      & and_dcpl_91;
  assign not_408_nl = ~ or_dcpl_156;
  assign x_max_lut_and_12_nl = MUX_v_3_2_2(3'b000, (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_4_mx0[2:0]),
      not_408_nl);
  assign x_max_lut_x_max_lut_or_12_nl = MUX_v_3_2_2(x_max_lut_and_12_nl, 3'b111,
      and_dcpl_89);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_3_nl =  -(ac_float_cctor_round_20_if_m_1_acc_3_tmp[3:0]);
  assign out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_3_nl = nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_3_nl[3:0];
  assign out_adpfloat_AdpfloatType_and_25_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_3_tmp[6]))
      & and_dcpl_91;
  assign out_adpfloat_AdpfloatType_mux_27_nl = MUX_v_4_2_2(out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_3_nl,
      (ac_float_cctor_round_20_if_m_1_acc_3_tmp[3:0]), out_adpfloat_AdpfloatType_and_25_nl);
  assign not_409_nl = ~ or_dcpl_156;
  assign out_adpfloat_AdpfloatType_and_24_nl = MUX_v_4_2_2(4'b0000, out_adpfloat_AdpfloatType_mux_27_nl,
      not_409_nl);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_12_nl = MUX_v_4_2_2(out_adpfloat_AdpfloatType_and_24_nl,
      4'b1111, and_dcpl_89);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_13_nl = (ac_float_cctor_round_20_if_m_1_acc_2_tmp[6])
      & and_dcpl_68;
  assign not_410_nl = ~ or_dcpl_136;
  assign x_max_lut_and_13_nl = MUX_v_3_2_2(3'b000, (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_3_mx0[2:0]),
      not_410_nl);
  assign x_max_lut_x_max_lut_or_13_nl = MUX_v_3_2_2(x_max_lut_and_13_nl, 3'b111,
      and_dcpl_66);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_2_nl =  -(ac_float_cctor_round_20_if_m_1_acc_2_tmp[3:0]);
  assign out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_2_nl = nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_2_nl[3:0];
  assign out_adpfloat_AdpfloatType_and_27_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_2_tmp[6]))
      & and_dcpl_68;
  assign out_adpfloat_AdpfloatType_mux_28_nl = MUX_v_4_2_2(out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_2_nl,
      (ac_float_cctor_round_20_if_m_1_acc_2_tmp[3:0]), out_adpfloat_AdpfloatType_and_27_nl);
  assign not_411_nl = ~ or_dcpl_136;
  assign out_adpfloat_AdpfloatType_and_26_nl = MUX_v_4_2_2(4'b0000, out_adpfloat_AdpfloatType_mux_28_nl,
      not_411_nl);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_13_nl = MUX_v_4_2_2(out_adpfloat_AdpfloatType_and_26_nl,
      4'b1111, and_dcpl_66);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_14_nl = (ac_float_cctor_round_20_if_m_1_acc_1_tmp[6])
      & and_dcpl_45;
  assign not_412_nl = ~ or_dcpl_116;
  assign x_max_lut_and_14_nl = MUX_v_3_2_2(3'b000, (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_2_mx0[2:0]),
      not_412_nl);
  assign x_max_lut_x_max_lut_or_14_nl = MUX_v_3_2_2(x_max_lut_and_14_nl, 3'b111,
      and_dcpl_43);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_1_nl =  -(ac_float_cctor_round_20_if_m_1_acc_1_tmp[3:0]);
  assign out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_1_nl = nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_1_nl[3:0];
  assign out_adpfloat_AdpfloatType_and_29_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_1_tmp[6]))
      & and_dcpl_45;
  assign out_adpfloat_AdpfloatType_mux_29_nl = MUX_v_4_2_2(out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_1_nl,
      (ac_float_cctor_round_20_if_m_1_acc_1_tmp[3:0]), out_adpfloat_AdpfloatType_and_29_nl);
  assign not_413_nl = ~ or_dcpl_116;
  assign out_adpfloat_AdpfloatType_and_28_nl = MUX_v_4_2_2(4'b0000, out_adpfloat_AdpfloatType_mux_29_nl,
      not_413_nl);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_14_nl = MUX_v_4_2_2(out_adpfloat_AdpfloatType_and_28_nl,
      4'b1111, and_dcpl_43);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_15_nl = (ac_float_cctor_round_20_if_m_1_acc_tmp[6])
      & and_dcpl_22;
  assign not_414_nl = ~ or_dcpl_96;
  assign x_max_lut_and_15_nl = MUX_v_3_2_2(3'b000, (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_1_mx0[2:0]),
      not_414_nl);
  assign x_max_lut_x_max_lut_or_15_nl = MUX_v_3_2_2(x_max_lut_and_15_nl, 3'b111,
      and_dcpl_20);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_nl =  -(ac_float_cctor_round_20_if_m_1_acc_tmp[3:0]);
  assign out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_nl = nl_out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_nl[3:0];
  assign out_adpfloat_AdpfloatType_and_31_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_tmp[6]))
      & and_dcpl_22;
  assign out_adpfloat_AdpfloatType_mux_30_nl = MUX_v_4_2_2(out_adpfloat_set_value_fixed_20U_14U_else_1_else_if_acc_nl,
      (ac_float_cctor_round_20_if_m_1_acc_tmp[3:0]), out_adpfloat_AdpfloatType_and_31_nl);
  assign not_415_nl = ~ or_dcpl_96;
  assign out_adpfloat_AdpfloatType_and_30_nl = MUX_v_4_2_2(4'b0000, out_adpfloat_AdpfloatType_mux_30_nl,
      not_415_nl);
  assign out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_15_nl = MUX_v_4_2_2(out_adpfloat_AdpfloatType_and_30_nl,
      4'b1111, and_dcpl_20);
  assign out_data = {out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_nl ,
      x_max_lut_x_max_lut_or_nl , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_nl
      , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_1_nl , x_max_lut_x_max_lut_or_1_nl
      , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_1_nl , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_2_nl
      , x_max_lut_x_max_lut_or_2_nl , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_2_nl
      , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_3_nl , x_max_lut_x_max_lut_or_3_nl
      , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_3_nl , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_4_nl
      , x_max_lut_x_max_lut_or_4_nl , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_4_nl
      , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_5_nl , x_max_lut_x_max_lut_or_5_nl
      , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_5_nl , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_6_nl
      , x_max_lut_x_max_lut_or_6_nl , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_6_nl
      , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_7_nl , x_max_lut_x_max_lut_or_7_nl
      , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_7_nl , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_8_nl
      , x_max_lut_x_max_lut_or_8_nl , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_8_nl
      , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_9_nl , x_max_lut_x_max_lut_or_9_nl
      , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_9_nl , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_10_nl
      , x_max_lut_x_max_lut_or_10_nl , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_10_nl
      , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_11_nl , x_max_lut_x_max_lut_or_11_nl
      , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_11_nl , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_12_nl
      , x_max_lut_x_max_lut_or_12_nl , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_12_nl
      , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_13_nl , x_max_lut_x_max_lut_or_13_nl
      , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_13_nl , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_14_nl
      , x_max_lut_x_max_lut_or_14_nl , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_14_nl
      , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_and_15_nl , x_max_lut_x_max_lut_or_15_nl
      , out_adpfloat_AdpfloatType_out_adpfloat_AdpfloatType_or_15_nl};
  assign nl_operator_24_true_operator_24_true_conc_mx0w1_5_1 = (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_16[5:1])
      + 5'b00101;
  assign operator_24_true_operator_24_true_conc_mx0w1_5_1 = nl_operator_24_true_operator_24_true_conc_mx0w1_5_1[4:0];
  assign nl_operator_23_true_acc_nl = ({operator_24_true_operator_24_true_conc_mx0w1_5_1
      , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_16[0])}) + 6'b000001;
  assign operator_23_true_acc_nl = nl_operator_23_true_acc_nl[5:0];
  assign or_5_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_tmp[6])) | (ac_float_cctor_round_20_if_m_1_acc_tmp[0])
      | (ac_float_cctor_round_20_if_m_1_acc_tmp[1]) | (ac_float_cctor_round_20_if_m_1_acc_tmp[2])
      | (ac_float_cctor_round_20_if_m_1_acc_tmp[3]) | (ac_float_cctor_round_20_if_m_1_acc_tmp[4]);
  assign out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_1_mx0 = MUX_v_6_2_2(operator_23_true_acc_nl,
      ({operator_24_true_operator_24_true_conc_mx0w1_5_1 , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_16[0])}),
      or_5_nl);
  assign ac_float_cctor_round_20_if_and_nl = (ac_float_cctor_round_20_if_m_1_acc_tmp[6:5]==2'b01);
  assign nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = ({5'b10010 , ac_float_cctor_round_20_if_and_nl}) + conv_u2s_5_6(~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_63)
      + 6'b000001;
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_nl =
      nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[5:0];
  assign or_nl = (in_data[0]) | (~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_47);
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_15_nl
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      or_nl);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_16 = ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_15_nl
      + conv_s2s_4_6({1'b1 , (~ adpfloat_bias)}) + 6'b000001;
  assign out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_16 = nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_16[5:0];
  assign nl_ac_float_cctor_round_20_if_m_1_acc_tmp = conv_s2u_6_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_itm[19:14])
      + conv_u2u_1_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_itm[13]);
  assign ac_float_cctor_round_20_if_m_1_acc_tmp = nl_ac_float_cctor_round_20_if_m_1_acc_tmp[6:0];
  assign nl_operator_24_true_operator_24_true_conc_3_mx0w1_5_1 = (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_17[5:1])
      + 5'b00101;
  assign operator_24_true_operator_24_true_conc_3_mx0w1_5_1 = nl_operator_24_true_operator_24_true_conc_3_mx0w1_5_1[4:0];
  assign nl_operator_23_true_acc_1_nl = ({operator_24_true_operator_24_true_conc_3_mx0w1_5_1
      , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_17[0])}) + 6'b000001;
  assign operator_23_true_acc_1_nl = nl_operator_23_true_acc_1_nl[5:0];
  assign or_11_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_1_tmp[6])) | (ac_float_cctor_round_20_if_m_1_acc_1_tmp[0])
      | (ac_float_cctor_round_20_if_m_1_acc_1_tmp[1]) | (ac_float_cctor_round_20_if_m_1_acc_1_tmp[2])
      | (ac_float_cctor_round_20_if_m_1_acc_1_tmp[3]) | (ac_float_cctor_round_20_if_m_1_acc_1_tmp[4]);
  assign out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_2_mx0 = MUX_v_6_2_2(operator_23_true_acc_1_nl,
      ({operator_24_true_operator_24_true_conc_3_mx0w1_5_1 , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_17[0])}),
      or_11_nl);
  assign ac_float_cctor_round_20_if_and_1_nl = (ac_float_cctor_round_20_if_m_1_acc_1_tmp[6:5]==2'b01);
  assign nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_1_nl
      = ({5'b10010 , ac_float_cctor_round_20_if_and_1_nl}) + conv_u2s_5_6(~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_62)
      + 6'b000001;
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_1_nl
      = nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_1_nl[5:0];
  assign or_6_nl = (in_data[20]) | (~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_46);
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_14_nl
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_1_nl,
      or_6_nl);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_17 = ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_14_nl
      + conv_s2s_4_6({1'b1 , (~ adpfloat_bias)}) + 6'b000001;
  assign out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_17 = nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_17[5:0];
  assign nl_ac_float_cctor_round_20_if_m_1_acc_1_tmp = conv_s2u_6_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_1_itm[19:14])
      + conv_u2u_1_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_1_itm[13]);
  assign ac_float_cctor_round_20_if_m_1_acc_1_tmp = nl_ac_float_cctor_round_20_if_m_1_acc_1_tmp[6:0];
  assign nl_operator_24_true_operator_24_true_conc_5_mx0w1_5_1 = (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_18[5:1])
      + 5'b00101;
  assign operator_24_true_operator_24_true_conc_5_mx0w1_5_1 = nl_operator_24_true_operator_24_true_conc_5_mx0w1_5_1[4:0];
  assign nl_operator_23_true_acc_2_nl = ({operator_24_true_operator_24_true_conc_5_mx0w1_5_1
      , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_18[0])}) + 6'b000001;
  assign operator_23_true_acc_2_nl = nl_operator_23_true_acc_2_nl[5:0];
  assign or_17_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_2_tmp[6])) | (ac_float_cctor_round_20_if_m_1_acc_2_tmp[0])
      | (ac_float_cctor_round_20_if_m_1_acc_2_tmp[1]) | (ac_float_cctor_round_20_if_m_1_acc_2_tmp[2])
      | (ac_float_cctor_round_20_if_m_1_acc_2_tmp[3]) | (ac_float_cctor_round_20_if_m_1_acc_2_tmp[4]);
  assign out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_3_mx0 = MUX_v_6_2_2(operator_23_true_acc_2_nl,
      ({operator_24_true_operator_24_true_conc_5_mx0w1_5_1 , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_18[0])}),
      or_17_nl);
  assign ac_float_cctor_round_20_if_and_2_nl = (ac_float_cctor_round_20_if_m_1_acc_2_tmp[6:5]==2'b01);
  assign nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_2_nl
      = ({5'b10010 , ac_float_cctor_round_20_if_and_2_nl}) + conv_u2s_5_6(~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_61)
      + 6'b000001;
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_2_nl
      = nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_2_nl[5:0];
  assign or_12_nl = (in_data[40]) | (~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_45);
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_13_nl
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_2_nl,
      or_12_nl);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_18 = ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_13_nl
      + conv_s2s_4_6({1'b1 , (~ adpfloat_bias)}) + 6'b000001;
  assign out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_18 = nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_18[5:0];
  assign nl_ac_float_cctor_round_20_if_m_1_acc_2_tmp = conv_s2u_6_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_2_itm[19:14])
      + conv_u2u_1_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_2_itm[13]);
  assign ac_float_cctor_round_20_if_m_1_acc_2_tmp = nl_ac_float_cctor_round_20_if_m_1_acc_2_tmp[6:0];
  assign nl_operator_24_true_operator_24_true_conc_7_mx0w1_5_1 = (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_19[5:1])
      + 5'b00101;
  assign operator_24_true_operator_24_true_conc_7_mx0w1_5_1 = nl_operator_24_true_operator_24_true_conc_7_mx0w1_5_1[4:0];
  assign nl_operator_23_true_acc_3_nl = ({operator_24_true_operator_24_true_conc_7_mx0w1_5_1
      , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_19[0])}) + 6'b000001;
  assign operator_23_true_acc_3_nl = nl_operator_23_true_acc_3_nl[5:0];
  assign or_23_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_3_tmp[6])) | (ac_float_cctor_round_20_if_m_1_acc_3_tmp[0])
      | (ac_float_cctor_round_20_if_m_1_acc_3_tmp[1]) | (ac_float_cctor_round_20_if_m_1_acc_3_tmp[2])
      | (ac_float_cctor_round_20_if_m_1_acc_3_tmp[3]) | (ac_float_cctor_round_20_if_m_1_acc_3_tmp[4]);
  assign out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_4_mx0 = MUX_v_6_2_2(operator_23_true_acc_3_nl,
      ({operator_24_true_operator_24_true_conc_7_mx0w1_5_1 , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_19[0])}),
      or_23_nl);
  assign ac_float_cctor_round_20_if_and_3_nl = (ac_float_cctor_round_20_if_m_1_acc_3_tmp[6:5]==2'b01);
  assign nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_3_nl
      = ({5'b10010 , ac_float_cctor_round_20_if_and_3_nl}) + conv_u2s_5_6(~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_60)
      + 6'b000001;
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_3_nl
      = nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_3_nl[5:0];
  assign or_18_nl = (in_data[60]) | (~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_44);
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_12_nl
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_3_nl,
      or_18_nl);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_19 = ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_12_nl
      + conv_s2s_4_6({1'b1 , (~ adpfloat_bias)}) + 6'b000001;
  assign out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_19 = nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_19[5:0];
  assign nl_ac_float_cctor_round_20_if_m_1_acc_3_tmp = conv_s2u_6_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_3_itm[19:14])
      + conv_u2u_1_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_3_itm[13]);
  assign ac_float_cctor_round_20_if_m_1_acc_3_tmp = nl_ac_float_cctor_round_20_if_m_1_acc_3_tmp[6:0];
  assign nl_operator_24_true_operator_24_true_conc_9_mx0w1_5_1 = (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_20[5:1])
      + 5'b00101;
  assign operator_24_true_operator_24_true_conc_9_mx0w1_5_1 = nl_operator_24_true_operator_24_true_conc_9_mx0w1_5_1[4:0];
  assign nl_operator_23_true_acc_4_nl = ({operator_24_true_operator_24_true_conc_9_mx0w1_5_1
      , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_20[0])}) + 6'b000001;
  assign operator_23_true_acc_4_nl = nl_operator_23_true_acc_4_nl[5:0];
  assign or_29_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_4_tmp[6])) | (ac_float_cctor_round_20_if_m_1_acc_4_tmp[0])
      | (ac_float_cctor_round_20_if_m_1_acc_4_tmp[1]) | (ac_float_cctor_round_20_if_m_1_acc_4_tmp[2])
      | (ac_float_cctor_round_20_if_m_1_acc_4_tmp[3]) | (ac_float_cctor_round_20_if_m_1_acc_4_tmp[4]);
  assign out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_5_mx0 = MUX_v_6_2_2(operator_23_true_acc_4_nl,
      ({operator_24_true_operator_24_true_conc_9_mx0w1_5_1 , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_20[0])}),
      or_29_nl);
  assign ac_float_cctor_round_20_if_and_4_nl = (ac_float_cctor_round_20_if_m_1_acc_4_tmp[6:5]==2'b01);
  assign nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_4_nl
      = ({5'b10010 , ac_float_cctor_round_20_if_and_4_nl}) + conv_u2s_5_6(~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_59)
      + 6'b000001;
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_4_nl
      = nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_4_nl[5:0];
  assign or_24_nl = (in_data[80]) | (~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_43);
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_11_nl
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_4_nl,
      or_24_nl);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_20 = ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_11_nl
      + conv_s2s_4_6({1'b1 , (~ adpfloat_bias)}) + 6'b000001;
  assign out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_20 = nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_20[5:0];
  assign nl_ac_float_cctor_round_20_if_m_1_acc_4_tmp = conv_s2u_6_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_4_itm[19:14])
      + conv_u2u_1_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_4_itm[13]);
  assign ac_float_cctor_round_20_if_m_1_acc_4_tmp = nl_ac_float_cctor_round_20_if_m_1_acc_4_tmp[6:0];
  assign nl_operator_24_true_operator_24_true_conc_11_mx0w1_5_1 = (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_21[5:1])
      + 5'b00101;
  assign operator_24_true_operator_24_true_conc_11_mx0w1_5_1 = nl_operator_24_true_operator_24_true_conc_11_mx0w1_5_1[4:0];
  assign nl_operator_23_true_acc_5_nl = ({operator_24_true_operator_24_true_conc_11_mx0w1_5_1
      , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_21[0])}) + 6'b000001;
  assign operator_23_true_acc_5_nl = nl_operator_23_true_acc_5_nl[5:0];
  assign or_35_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_5_tmp[6])) | (ac_float_cctor_round_20_if_m_1_acc_5_tmp[0])
      | (ac_float_cctor_round_20_if_m_1_acc_5_tmp[1]) | (ac_float_cctor_round_20_if_m_1_acc_5_tmp[2])
      | (ac_float_cctor_round_20_if_m_1_acc_5_tmp[3]) | (ac_float_cctor_round_20_if_m_1_acc_5_tmp[4]);
  assign out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_6_mx0 = MUX_v_6_2_2(operator_23_true_acc_5_nl,
      ({operator_24_true_operator_24_true_conc_11_mx0w1_5_1 , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_21[0])}),
      or_35_nl);
  assign ac_float_cctor_round_20_if_and_5_nl = (ac_float_cctor_round_20_if_m_1_acc_5_tmp[6:5]==2'b01);
  assign nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_5_nl
      = ({5'b10010 , ac_float_cctor_round_20_if_and_5_nl}) + conv_u2s_5_6(~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_58)
      + 6'b000001;
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_5_nl
      = nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_5_nl[5:0];
  assign or_30_nl = (in_data[100]) | (~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_42);
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_10_nl
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_5_nl,
      or_30_nl);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_21 = ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_10_nl
      + conv_s2s_4_6({1'b1 , (~ adpfloat_bias)}) + 6'b000001;
  assign out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_21 = nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_21[5:0];
  assign nl_ac_float_cctor_round_20_if_m_1_acc_5_tmp = conv_s2u_6_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_5_itm[19:14])
      + conv_u2u_1_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_5_itm[13]);
  assign ac_float_cctor_round_20_if_m_1_acc_5_tmp = nl_ac_float_cctor_round_20_if_m_1_acc_5_tmp[6:0];
  assign nl_operator_24_true_operator_24_true_conc_13_mx0w1_5_1 = (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_22[5:1])
      + 5'b00101;
  assign operator_24_true_operator_24_true_conc_13_mx0w1_5_1 = nl_operator_24_true_operator_24_true_conc_13_mx0w1_5_1[4:0];
  assign nl_operator_23_true_acc_6_nl = ({operator_24_true_operator_24_true_conc_13_mx0w1_5_1
      , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_22[0])}) + 6'b000001;
  assign operator_23_true_acc_6_nl = nl_operator_23_true_acc_6_nl[5:0];
  assign or_41_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_6_tmp[6])) | (ac_float_cctor_round_20_if_m_1_acc_6_tmp[0])
      | (ac_float_cctor_round_20_if_m_1_acc_6_tmp[1]) | (ac_float_cctor_round_20_if_m_1_acc_6_tmp[2])
      | (ac_float_cctor_round_20_if_m_1_acc_6_tmp[3]) | (ac_float_cctor_round_20_if_m_1_acc_6_tmp[4]);
  assign out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_7_mx0 = MUX_v_6_2_2(operator_23_true_acc_6_nl,
      ({operator_24_true_operator_24_true_conc_13_mx0w1_5_1 , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_22[0])}),
      or_41_nl);
  assign ac_float_cctor_round_20_if_and_6_nl = (ac_float_cctor_round_20_if_m_1_acc_6_tmp[6:5]==2'b01);
  assign nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_6_nl
      = ({5'b10010 , ac_float_cctor_round_20_if_and_6_nl}) + conv_u2s_5_6(~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_57)
      + 6'b000001;
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_6_nl
      = nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_6_nl[5:0];
  assign or_36_nl = (in_data[120]) | (~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_41);
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_9_nl
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_6_nl,
      or_36_nl);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_22 = ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_9_nl
      + conv_s2s_4_6({1'b1 , (~ adpfloat_bias)}) + 6'b000001;
  assign out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_22 = nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_22[5:0];
  assign nl_ac_float_cctor_round_20_if_m_1_acc_6_tmp = conv_s2u_6_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_6_itm[19:14])
      + conv_u2u_1_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_6_itm[13]);
  assign ac_float_cctor_round_20_if_m_1_acc_6_tmp = nl_ac_float_cctor_round_20_if_m_1_acc_6_tmp[6:0];
  assign nl_operator_24_true_operator_24_true_conc_15_mx0w1_5_1 = (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_23[5:1])
      + 5'b00101;
  assign operator_24_true_operator_24_true_conc_15_mx0w1_5_1 = nl_operator_24_true_operator_24_true_conc_15_mx0w1_5_1[4:0];
  assign nl_operator_23_true_acc_7_nl = ({operator_24_true_operator_24_true_conc_15_mx0w1_5_1
      , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_23[0])}) + 6'b000001;
  assign operator_23_true_acc_7_nl = nl_operator_23_true_acc_7_nl[5:0];
  assign or_47_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_7_tmp[6])) | (ac_float_cctor_round_20_if_m_1_acc_7_tmp[0])
      | (ac_float_cctor_round_20_if_m_1_acc_7_tmp[1]) | (ac_float_cctor_round_20_if_m_1_acc_7_tmp[2])
      | (ac_float_cctor_round_20_if_m_1_acc_7_tmp[3]) | (ac_float_cctor_round_20_if_m_1_acc_7_tmp[4]);
  assign out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_8_mx0 = MUX_v_6_2_2(operator_23_true_acc_7_nl,
      ({operator_24_true_operator_24_true_conc_15_mx0w1_5_1 , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_23[0])}),
      or_47_nl);
  assign ac_float_cctor_round_20_if_and_7_nl = (ac_float_cctor_round_20_if_m_1_acc_7_tmp[6:5]==2'b01);
  assign nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_7_nl
      = ({5'b10010 , ac_float_cctor_round_20_if_and_7_nl}) + conv_u2s_5_6(~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_56)
      + 6'b000001;
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_7_nl
      = nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_7_nl[5:0];
  assign or_42_nl = (in_data[140]) | (~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_40);
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_8_nl
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_7_nl,
      or_42_nl);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_23 = ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_8_nl
      + conv_s2s_4_6({1'b1 , (~ adpfloat_bias)}) + 6'b000001;
  assign out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_23 = nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_23[5:0];
  assign nl_ac_float_cctor_round_20_if_m_1_acc_7_tmp = conv_s2u_6_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_7_itm[19:14])
      + conv_u2u_1_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_7_itm[13]);
  assign ac_float_cctor_round_20_if_m_1_acc_7_tmp = nl_ac_float_cctor_round_20_if_m_1_acc_7_tmp[6:0];
  assign nl_operator_24_true_operator_24_true_conc_17_mx0w1_5_1 = (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_24[5:1])
      + 5'b00101;
  assign operator_24_true_operator_24_true_conc_17_mx0w1_5_1 = nl_operator_24_true_operator_24_true_conc_17_mx0w1_5_1[4:0];
  assign nl_operator_23_true_acc_8_nl = ({operator_24_true_operator_24_true_conc_17_mx0w1_5_1
      , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_24[0])}) + 6'b000001;
  assign operator_23_true_acc_8_nl = nl_operator_23_true_acc_8_nl[5:0];
  assign or_53_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_8_tmp[6])) | (ac_float_cctor_round_20_if_m_1_acc_8_tmp[0])
      | (ac_float_cctor_round_20_if_m_1_acc_8_tmp[1]) | (ac_float_cctor_round_20_if_m_1_acc_8_tmp[2])
      | (ac_float_cctor_round_20_if_m_1_acc_8_tmp[3]) | (ac_float_cctor_round_20_if_m_1_acc_8_tmp[4]);
  assign out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_9_mx0 = MUX_v_6_2_2(operator_23_true_acc_8_nl,
      ({operator_24_true_operator_24_true_conc_17_mx0w1_5_1 , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_24[0])}),
      or_53_nl);
  assign ac_float_cctor_round_20_if_and_8_nl = (ac_float_cctor_round_20_if_m_1_acc_8_tmp[6:5]==2'b01);
  assign nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_8_nl
      = ({5'b10010 , ac_float_cctor_round_20_if_and_8_nl}) + conv_u2s_5_6(~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_55)
      + 6'b000001;
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_8_nl
      = nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_8_nl[5:0];
  assign or_48_nl = (in_data[160]) | (~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_39);
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_7_nl
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_8_nl,
      or_48_nl);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_24 = ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_7_nl
      + conv_s2s_4_6({1'b1 , (~ adpfloat_bias)}) + 6'b000001;
  assign out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_24 = nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_24[5:0];
  assign nl_ac_float_cctor_round_20_if_m_1_acc_8_tmp = conv_s2u_6_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_8_itm[19:14])
      + conv_u2u_1_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_8_itm[13]);
  assign ac_float_cctor_round_20_if_m_1_acc_8_tmp = nl_ac_float_cctor_round_20_if_m_1_acc_8_tmp[6:0];
  assign nl_operator_24_true_operator_24_true_conc_19_mx0w1_5_1 = (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_25[5:1])
      + 5'b00101;
  assign operator_24_true_operator_24_true_conc_19_mx0w1_5_1 = nl_operator_24_true_operator_24_true_conc_19_mx0w1_5_1[4:0];
  assign nl_operator_23_true_acc_9_nl = ({operator_24_true_operator_24_true_conc_19_mx0w1_5_1
      , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_25[0])}) + 6'b000001;
  assign operator_23_true_acc_9_nl = nl_operator_23_true_acc_9_nl[5:0];
  assign or_59_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_9_tmp[6])) | (ac_float_cctor_round_20_if_m_1_acc_9_tmp[0])
      | (ac_float_cctor_round_20_if_m_1_acc_9_tmp[1]) | (ac_float_cctor_round_20_if_m_1_acc_9_tmp[2])
      | (ac_float_cctor_round_20_if_m_1_acc_9_tmp[3]) | (ac_float_cctor_round_20_if_m_1_acc_9_tmp[4]);
  assign out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_10_mx0 = MUX_v_6_2_2(operator_23_true_acc_9_nl,
      ({operator_24_true_operator_24_true_conc_19_mx0w1_5_1 , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_25[0])}),
      or_59_nl);
  assign ac_float_cctor_round_20_if_and_9_nl = (ac_float_cctor_round_20_if_m_1_acc_9_tmp[6:5]==2'b01);
  assign nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_9_nl
      = ({5'b10010 , ac_float_cctor_round_20_if_and_9_nl}) + conv_u2s_5_6(~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_54)
      + 6'b000001;
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_9_nl
      = nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_9_nl[5:0];
  assign or_54_nl = (in_data[180]) | (~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_38);
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_6_nl
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_9_nl,
      or_54_nl);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_25 = ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_6_nl
      + conv_s2s_4_6({1'b1 , (~ adpfloat_bias)}) + 6'b000001;
  assign out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_25 = nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_25[5:0];
  assign nl_ac_float_cctor_round_20_if_m_1_acc_9_tmp = conv_s2u_6_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_9_itm[19:14])
      + conv_u2u_1_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_9_itm[13]);
  assign ac_float_cctor_round_20_if_m_1_acc_9_tmp = nl_ac_float_cctor_round_20_if_m_1_acc_9_tmp[6:0];
  assign nl_operator_24_true_operator_24_true_conc_21_mx0w1_5_1 = (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_26[5:1])
      + 5'b00101;
  assign operator_24_true_operator_24_true_conc_21_mx0w1_5_1 = nl_operator_24_true_operator_24_true_conc_21_mx0w1_5_1[4:0];
  assign nl_operator_23_true_acc_10_nl = ({operator_24_true_operator_24_true_conc_21_mx0w1_5_1
      , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_26[0])}) + 6'b000001;
  assign operator_23_true_acc_10_nl = nl_operator_23_true_acc_10_nl[5:0];
  assign or_65_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_10_tmp[6])) | (ac_float_cctor_round_20_if_m_1_acc_10_tmp[0])
      | (ac_float_cctor_round_20_if_m_1_acc_10_tmp[1]) | (ac_float_cctor_round_20_if_m_1_acc_10_tmp[2])
      | (ac_float_cctor_round_20_if_m_1_acc_10_tmp[3]) | (ac_float_cctor_round_20_if_m_1_acc_10_tmp[4]);
  assign out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_11_mx0 = MUX_v_6_2_2(operator_23_true_acc_10_nl,
      ({operator_24_true_operator_24_true_conc_21_mx0w1_5_1 , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_26[0])}),
      or_65_nl);
  assign ac_float_cctor_round_20_if_and_10_nl = (ac_float_cctor_round_20_if_m_1_acc_10_tmp[6:5]==2'b01);
  assign nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_10_nl
      = ({5'b10010 , ac_float_cctor_round_20_if_and_10_nl}) + conv_u2s_5_6(~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_53)
      + 6'b000001;
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_10_nl
      = nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_10_nl[5:0];
  assign or_60_nl = (in_data[200]) | (~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_37);
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_5_nl
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_10_nl,
      or_60_nl);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_26 = ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_5_nl
      + conv_s2s_4_6({1'b1 , (~ adpfloat_bias)}) + 6'b000001;
  assign out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_26 = nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_26[5:0];
  assign nl_ac_float_cctor_round_20_if_m_1_acc_10_tmp = conv_s2u_6_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_10_itm[19:14])
      + conv_u2u_1_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_10_itm[13]);
  assign ac_float_cctor_round_20_if_m_1_acc_10_tmp = nl_ac_float_cctor_round_20_if_m_1_acc_10_tmp[6:0];
  assign nl_operator_24_true_operator_24_true_conc_23_mx0w1_5_1 = (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_27[5:1])
      + 5'b00101;
  assign operator_24_true_operator_24_true_conc_23_mx0w1_5_1 = nl_operator_24_true_operator_24_true_conc_23_mx0w1_5_1[4:0];
  assign nl_operator_23_true_acc_11_nl = ({operator_24_true_operator_24_true_conc_23_mx0w1_5_1
      , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_27[0])}) + 6'b000001;
  assign operator_23_true_acc_11_nl = nl_operator_23_true_acc_11_nl[5:0];
  assign or_71_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_11_tmp[6])) | (ac_float_cctor_round_20_if_m_1_acc_11_tmp[0])
      | (ac_float_cctor_round_20_if_m_1_acc_11_tmp[1]) | (ac_float_cctor_round_20_if_m_1_acc_11_tmp[2])
      | (ac_float_cctor_round_20_if_m_1_acc_11_tmp[3]) | (ac_float_cctor_round_20_if_m_1_acc_11_tmp[4]);
  assign out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_12_mx0 = MUX_v_6_2_2(operator_23_true_acc_11_nl,
      ({operator_24_true_operator_24_true_conc_23_mx0w1_5_1 , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_27[0])}),
      or_71_nl);
  assign ac_float_cctor_round_20_if_and_11_nl = (ac_float_cctor_round_20_if_m_1_acc_11_tmp[6:5]==2'b01);
  assign nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_11_nl
      = ({5'b10010 , ac_float_cctor_round_20_if_and_11_nl}) + conv_u2s_5_6(~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_52)
      + 6'b000001;
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_11_nl
      = nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_11_nl[5:0];
  assign or_66_nl = (in_data[220]) | (~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_36);
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_4_nl
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_11_nl,
      or_66_nl);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_27 = ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_4_nl
      + conv_s2s_4_6({1'b1 , (~ adpfloat_bias)}) + 6'b000001;
  assign out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_27 = nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_27[5:0];
  assign nl_ac_float_cctor_round_20_if_m_1_acc_11_tmp = conv_s2u_6_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_11_itm[19:14])
      + conv_u2u_1_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_11_itm[13]);
  assign ac_float_cctor_round_20_if_m_1_acc_11_tmp = nl_ac_float_cctor_round_20_if_m_1_acc_11_tmp[6:0];
  assign nl_operator_24_true_operator_24_true_conc_25_mx0w1_5_1 = (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_28[5:1])
      + 5'b00101;
  assign operator_24_true_operator_24_true_conc_25_mx0w1_5_1 = nl_operator_24_true_operator_24_true_conc_25_mx0w1_5_1[4:0];
  assign nl_operator_23_true_acc_12_nl = ({operator_24_true_operator_24_true_conc_25_mx0w1_5_1
      , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_28[0])}) + 6'b000001;
  assign operator_23_true_acc_12_nl = nl_operator_23_true_acc_12_nl[5:0];
  assign or_77_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_12_tmp[6])) | (ac_float_cctor_round_20_if_m_1_acc_12_tmp[0])
      | (ac_float_cctor_round_20_if_m_1_acc_12_tmp[1]) | (ac_float_cctor_round_20_if_m_1_acc_12_tmp[2])
      | (ac_float_cctor_round_20_if_m_1_acc_12_tmp[3]) | (ac_float_cctor_round_20_if_m_1_acc_12_tmp[4]);
  assign out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_13_mx0 = MUX_v_6_2_2(operator_23_true_acc_12_nl,
      ({operator_24_true_operator_24_true_conc_25_mx0w1_5_1 , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_28[0])}),
      or_77_nl);
  assign ac_float_cctor_round_20_if_and_12_nl = (ac_float_cctor_round_20_if_m_1_acc_12_tmp[6:5]==2'b01);
  assign nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_12_nl
      = ({5'b10010 , ac_float_cctor_round_20_if_and_12_nl}) + conv_u2s_5_6(~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_51)
      + 6'b000001;
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_12_nl
      = nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_12_nl[5:0];
  assign or_72_nl = (in_data[240]) | (~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_35);
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_3_nl
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_12_nl,
      or_72_nl);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_28 = ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_3_nl
      + conv_s2s_4_6({1'b1 , (~ adpfloat_bias)}) + 6'b000001;
  assign out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_28 = nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_28[5:0];
  assign nl_ac_float_cctor_round_20_if_m_1_acc_12_tmp = conv_s2u_6_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_12_itm[19:14])
      + conv_u2u_1_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_12_itm[13]);
  assign ac_float_cctor_round_20_if_m_1_acc_12_tmp = nl_ac_float_cctor_round_20_if_m_1_acc_12_tmp[6:0];
  assign nl_operator_24_true_operator_24_true_conc_27_mx0w1_5_1 = (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_29[5:1])
      + 5'b00101;
  assign operator_24_true_operator_24_true_conc_27_mx0w1_5_1 = nl_operator_24_true_operator_24_true_conc_27_mx0w1_5_1[4:0];
  assign nl_operator_23_true_acc_13_nl = ({operator_24_true_operator_24_true_conc_27_mx0w1_5_1
      , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_29[0])}) + 6'b000001;
  assign operator_23_true_acc_13_nl = nl_operator_23_true_acc_13_nl[5:0];
  assign or_83_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_13_tmp[6])) | (ac_float_cctor_round_20_if_m_1_acc_13_tmp[0])
      | (ac_float_cctor_round_20_if_m_1_acc_13_tmp[1]) | (ac_float_cctor_round_20_if_m_1_acc_13_tmp[2])
      | (ac_float_cctor_round_20_if_m_1_acc_13_tmp[3]) | (ac_float_cctor_round_20_if_m_1_acc_13_tmp[4]);
  assign out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_14_mx0 = MUX_v_6_2_2(operator_23_true_acc_13_nl,
      ({operator_24_true_operator_24_true_conc_27_mx0w1_5_1 , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_29[0])}),
      or_83_nl);
  assign ac_float_cctor_round_20_if_and_13_nl = (ac_float_cctor_round_20_if_m_1_acc_13_tmp[6:5]==2'b01);
  assign nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_13_nl
      = ({5'b10010 , ac_float_cctor_round_20_if_and_13_nl}) + conv_u2s_5_6(~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_50)
      + 6'b000001;
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_13_nl
      = nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_13_nl[5:0];
  assign or_78_nl = (in_data[260]) | (~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_34);
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_2_nl
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_13_nl,
      or_78_nl);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_29 = ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_2_nl
      + conv_s2s_4_6({1'b1 , (~ adpfloat_bias)}) + 6'b000001;
  assign out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_29 = nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_29[5:0];
  assign nl_ac_float_cctor_round_20_if_m_1_acc_13_tmp = conv_s2u_6_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_13_itm[19:14])
      + conv_u2u_1_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_13_itm[13]);
  assign ac_float_cctor_round_20_if_m_1_acc_13_tmp = nl_ac_float_cctor_round_20_if_m_1_acc_13_tmp[6:0];
  assign nl_operator_24_true_operator_24_true_conc_29_mx0w1_5_1 = (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_30[5:1])
      + 5'b00101;
  assign operator_24_true_operator_24_true_conc_29_mx0w1_5_1 = nl_operator_24_true_operator_24_true_conc_29_mx0w1_5_1[4:0];
  assign nl_operator_23_true_acc_14_nl = ({operator_24_true_operator_24_true_conc_29_mx0w1_5_1
      , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_30[0])}) + 6'b000001;
  assign operator_23_true_acc_14_nl = nl_operator_23_true_acc_14_nl[5:0];
  assign or_89_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_14_tmp[6])) | (ac_float_cctor_round_20_if_m_1_acc_14_tmp[0])
      | (ac_float_cctor_round_20_if_m_1_acc_14_tmp[1]) | (ac_float_cctor_round_20_if_m_1_acc_14_tmp[2])
      | (ac_float_cctor_round_20_if_m_1_acc_14_tmp[3]) | (ac_float_cctor_round_20_if_m_1_acc_14_tmp[4]);
  assign out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_15_mx0 = MUX_v_6_2_2(operator_23_true_acc_14_nl,
      ({operator_24_true_operator_24_true_conc_29_mx0w1_5_1 , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_30[0])}),
      or_89_nl);
  assign ac_float_cctor_round_20_if_and_14_nl = (ac_float_cctor_round_20_if_m_1_acc_14_tmp[6:5]==2'b01);
  assign nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_14_nl
      = ({5'b10010 , ac_float_cctor_round_20_if_and_14_nl}) + conv_u2s_5_6(~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_49)
      + 6'b000001;
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_14_nl
      = nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_14_nl[5:0];
  assign or_84_nl = (in_data[280]) | (~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_33);
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_1_nl
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_14_nl,
      or_84_nl);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_30 = ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_1_nl
      + conv_s2s_4_6({1'b1 , (~ adpfloat_bias)}) + 6'b000001;
  assign out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_30 = nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_30[5:0];
  assign nl_ac_float_cctor_round_20_if_m_1_acc_14_tmp = conv_s2u_6_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_14_itm[19:14])
      + conv_u2u_1_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_14_itm[13]);
  assign ac_float_cctor_round_20_if_m_1_acc_14_tmp = nl_ac_float_cctor_round_20_if_m_1_acc_14_tmp[6:0];
  assign nl_operator_24_true_operator_24_true_conc_31_mx0w1_5_1 = (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_31[5:1])
      + 5'b00101;
  assign operator_24_true_operator_24_true_conc_31_mx0w1_5_1 = nl_operator_24_true_operator_24_true_conc_31_mx0w1_5_1[4:0];
  assign nl_operator_23_true_acc_15_nl = ({operator_24_true_operator_24_true_conc_31_mx0w1_5_1
      , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_31[0])}) + 6'b000001;
  assign operator_23_true_acc_15_nl = nl_operator_23_true_acc_15_nl[5:0];
  assign or_95_nl = (~ (ac_float_cctor_round_20_if_m_1_acc_15_tmp[6])) | (ac_float_cctor_round_20_if_m_1_acc_15_tmp[0])
      | (ac_float_cctor_round_20_if_m_1_acc_15_tmp[1]) | (ac_float_cctor_round_20_if_m_1_acc_15_tmp[2])
      | (ac_float_cctor_round_20_if_m_1_acc_15_tmp[3]) | (ac_float_cctor_round_20_if_m_1_acc_15_tmp[4]);
  assign out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_mx0 = MUX_v_6_2_2(operator_23_true_acc_15_nl,
      ({operator_24_true_operator_24_true_conc_31_mx0w1_5_1 , (out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_31[0])}),
      or_95_nl);
  assign ac_float_cctor_round_20_if_and_15_nl = (ac_float_cctor_round_20_if_m_1_acc_15_tmp[6:5]==2'b01);
  assign nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_15_nl
      = ({5'b10010 , ac_float_cctor_round_20_if_and_15_nl}) + conv_u2s_5_6(~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_48)
      + 6'b000001;
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_15_nl
      = nl_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_15_nl[5:0];
  assign or_90_nl = (in_data[300]) | (~ libraries_leading_sign_20_1_1_0_76b0da59e271ffee6fadead7366344fb6166_32);
  assign ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_nl
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_else_1_qelse_acc_15_nl,
      or_90_nl);
  assign nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_31 = ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_ac_float_cctor_assign_from_0_0_20_6_AC_TRN_AC_WRAP_qif_and_nl
      + conv_s2s_4_6({1'b1 , (~ adpfloat_bias)}) + 6'b000001;
  assign out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_31 = nl_out_adpfloat_set_value_fixed_20U_14U_acc_psp_5_0_31[5:0];
  assign nl_ac_float_cctor_round_20_if_m_1_acc_15_tmp = conv_s2u_6_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_15_itm[19:14])
      + conv_u2u_1_7(operator_20_6_true_AC_TRN_AC_WRAP_lshift_15_itm[13]);
  assign ac_float_cctor_round_20_if_m_1_acc_15_tmp = nl_ac_float_cctor_round_20_if_m_1_acc_15_tmp[6:0];
  assign nl_operator_23_true_acc_15_nl_1 = (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_mx0[5:3])
      + 3'b111;
  assign operator_23_true_acc_15_nl_1 = nl_operator_23_true_acc_15_nl_1[2:0];
  assign operator_23_true_acc_15_itm_2_1 = readslicef_3_1_2(operator_23_true_acc_15_nl_1);
  assign nl_operator_23_true_acc_14_nl_1 = (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_15_mx0[5:3])
      + 3'b111;
  assign operator_23_true_acc_14_nl_1 = nl_operator_23_true_acc_14_nl_1[2:0];
  assign operator_23_true_acc_14_itm_2_1 = readslicef_3_1_2(operator_23_true_acc_14_nl_1);
  assign nl_operator_23_true_acc_13_nl_1 = (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_14_mx0[5:3])
      + 3'b111;
  assign operator_23_true_acc_13_nl_1 = nl_operator_23_true_acc_13_nl_1[2:0];
  assign operator_23_true_acc_13_itm_2_1 = readslicef_3_1_2(operator_23_true_acc_13_nl_1);
  assign nl_operator_23_true_acc_12_nl_1 = (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_13_mx0[5:3])
      + 3'b111;
  assign operator_23_true_acc_12_nl_1 = nl_operator_23_true_acc_12_nl_1[2:0];
  assign operator_23_true_acc_12_itm_2_1 = readslicef_3_1_2(operator_23_true_acc_12_nl_1);
  assign nl_operator_23_true_acc_11_nl_1 = (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_12_mx0[5:3])
      + 3'b111;
  assign operator_23_true_acc_11_nl_1 = nl_operator_23_true_acc_11_nl_1[2:0];
  assign operator_23_true_acc_11_itm_2_1 = readslicef_3_1_2(operator_23_true_acc_11_nl_1);
  assign nl_operator_23_true_acc_10_nl_1 = (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_11_mx0[5:3])
      + 3'b111;
  assign operator_23_true_acc_10_nl_1 = nl_operator_23_true_acc_10_nl_1[2:0];
  assign operator_23_true_acc_10_itm_2_1 = readslicef_3_1_2(operator_23_true_acc_10_nl_1);
  assign nl_operator_23_true_acc_9_nl_1 = (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_10_mx0[5:3])
      + 3'b111;
  assign operator_23_true_acc_9_nl_1 = nl_operator_23_true_acc_9_nl_1[2:0];
  assign operator_23_true_acc_9_itm_2_1 = readslicef_3_1_2(operator_23_true_acc_9_nl_1);
  assign nl_operator_23_true_acc_8_nl_1 = (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_9_mx0[5:3])
      + 3'b111;
  assign operator_23_true_acc_8_nl_1 = nl_operator_23_true_acc_8_nl_1[2:0];
  assign operator_23_true_acc_8_itm_2_1 = readslicef_3_1_2(operator_23_true_acc_8_nl_1);
  assign nl_operator_23_true_acc_7_nl_1 = (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_8_mx0[5:3])
      + 3'b111;
  assign operator_23_true_acc_7_nl_1 = nl_operator_23_true_acc_7_nl_1[2:0];
  assign operator_23_true_acc_7_itm_2_1 = readslicef_3_1_2(operator_23_true_acc_7_nl_1);
  assign nl_operator_23_true_acc_6_nl_1 = (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_7_mx0[5:3])
      + 3'b111;
  assign operator_23_true_acc_6_nl_1 = nl_operator_23_true_acc_6_nl_1[2:0];
  assign operator_23_true_acc_6_itm_2_1 = readslicef_3_1_2(operator_23_true_acc_6_nl_1);
  assign nl_operator_23_true_acc_5_nl_1 = (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_6_mx0[5:3])
      + 3'b111;
  assign operator_23_true_acc_5_nl_1 = nl_operator_23_true_acc_5_nl_1[2:0];
  assign operator_23_true_acc_5_itm_2_1 = readslicef_3_1_2(operator_23_true_acc_5_nl_1);
  assign nl_operator_23_true_acc_4_nl_1 = (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_5_mx0[5:3])
      + 3'b111;
  assign operator_23_true_acc_4_nl_1 = nl_operator_23_true_acc_4_nl_1[2:0];
  assign operator_23_true_acc_4_itm_2_1 = readslicef_3_1_2(operator_23_true_acc_4_nl_1);
  assign nl_operator_23_true_acc_3_nl_1 = (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_4_mx0[5:3])
      + 3'b111;
  assign operator_23_true_acc_3_nl_1 = nl_operator_23_true_acc_3_nl_1[2:0];
  assign operator_23_true_acc_3_itm_2_1 = readslicef_3_1_2(operator_23_true_acc_3_nl_1);
  assign nl_operator_23_true_acc_2_nl_1 = (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_3_mx0[5:3])
      + 3'b111;
  assign operator_23_true_acc_2_nl_1 = nl_operator_23_true_acc_2_nl_1[2:0];
  assign operator_23_true_acc_2_itm_2_1 = readslicef_3_1_2(operator_23_true_acc_2_nl_1);
  assign nl_operator_23_true_acc_1_nl_1 = (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_2_mx0[5:3])
      + 3'b111;
  assign operator_23_true_acc_1_nl_1 = nl_operator_23_true_acc_1_nl_1[2:0];
  assign operator_23_true_acc_1_itm_2_1 = readslicef_3_1_2(operator_23_true_acc_1_nl_1);
  assign nl_operator_23_true_acc_nl_1 = (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_1_mx0[5:3])
      + 3'b111;
  assign operator_23_true_acc_nl_1 = nl_operator_23_true_acc_nl_1[2:0];
  assign operator_23_true_acc_itm_2_1 = readslicef_3_1_2(operator_23_true_acc_nl_1);
  assign or_dcpl_96 = ((in_data[19:0]==20'b00000000000000000000)) | (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_1_mx0[5]);
  assign or_dcpl_115 = (in_data[19:0]!=20'b00000000000000000000);
  assign and_dcpl_20 = or_dcpl_115 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_1_mx0[5]))
      & (~ operator_23_true_acc_itm_2_1);
  assign and_dcpl_22 = or_dcpl_115 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_1_mx0[5]))
      & operator_23_true_acc_itm_2_1;
  assign or_dcpl_116 = ((in_data[39:20]==20'b00000000000000000000)) | (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_2_mx0[5]);
  assign or_dcpl_135 = (in_data[39:20]!=20'b00000000000000000000);
  assign and_dcpl_43 = or_dcpl_135 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_2_mx0[5]))
      & (~ operator_23_true_acc_1_itm_2_1);
  assign and_dcpl_45 = or_dcpl_135 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_2_mx0[5]))
      & operator_23_true_acc_1_itm_2_1;
  assign or_dcpl_136 = ((in_data[59:40]==20'b00000000000000000000)) | (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_3_mx0[5]);
  assign or_dcpl_155 = (in_data[59:40]!=20'b00000000000000000000);
  assign and_dcpl_66 = or_dcpl_155 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_3_mx0[5]))
      & (~ operator_23_true_acc_2_itm_2_1);
  assign and_dcpl_68 = or_dcpl_155 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_3_mx0[5]))
      & operator_23_true_acc_2_itm_2_1;
  assign or_dcpl_156 = ((in_data[79:60]==20'b00000000000000000000)) | (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_4_mx0[5]);
  assign or_dcpl_175 = (in_data[79:60]!=20'b00000000000000000000);
  assign and_dcpl_89 = or_dcpl_175 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_4_mx0[5]))
      & (~ operator_23_true_acc_3_itm_2_1);
  assign and_dcpl_91 = or_dcpl_175 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_4_mx0[5]))
      & operator_23_true_acc_3_itm_2_1;
  assign or_dcpl_176 = ((in_data[99:80]==20'b00000000000000000000)) | (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_5_mx0[5]);
  assign or_dcpl_195 = (in_data[99:80]!=20'b00000000000000000000);
  assign and_dcpl_112 = or_dcpl_195 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_5_mx0[5]))
      & (~ operator_23_true_acc_4_itm_2_1);
  assign and_dcpl_114 = or_dcpl_195 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_5_mx0[5]))
      & operator_23_true_acc_4_itm_2_1;
  assign or_dcpl_196 = ((in_data[119:100]==20'b00000000000000000000)) | (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_6_mx0[5]);
  assign or_dcpl_215 = (in_data[119:100]!=20'b00000000000000000000);
  assign and_dcpl_135 = or_dcpl_215 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_6_mx0[5]))
      & (~ operator_23_true_acc_5_itm_2_1);
  assign and_dcpl_137 = or_dcpl_215 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_6_mx0[5]))
      & operator_23_true_acc_5_itm_2_1;
  assign or_dcpl_216 = ((in_data[139:120]==20'b00000000000000000000)) | (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_7_mx0[5]);
  assign or_dcpl_235 = (in_data[139:120]!=20'b00000000000000000000);
  assign and_dcpl_158 = or_dcpl_235 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_7_mx0[5]))
      & (~ operator_23_true_acc_6_itm_2_1);
  assign and_dcpl_160 = or_dcpl_235 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_7_mx0[5]))
      & operator_23_true_acc_6_itm_2_1;
  assign or_dcpl_236 = ((in_data[159:140]==20'b00000000000000000000)) | (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_8_mx0[5]);
  assign or_dcpl_255 = (in_data[159:140]!=20'b00000000000000000000);
  assign and_dcpl_181 = or_dcpl_255 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_8_mx0[5]))
      & (~ operator_23_true_acc_7_itm_2_1);
  assign and_dcpl_183 = or_dcpl_255 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_8_mx0[5]))
      & operator_23_true_acc_7_itm_2_1;
  assign or_dcpl_256 = ((in_data[179:160]==20'b00000000000000000000)) | (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_9_mx0[5]);
  assign or_dcpl_275 = (in_data[179:160]!=20'b00000000000000000000);
  assign and_dcpl_204 = or_dcpl_275 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_9_mx0[5]))
      & (~ operator_23_true_acc_8_itm_2_1);
  assign and_dcpl_206 = or_dcpl_275 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_9_mx0[5]))
      & operator_23_true_acc_8_itm_2_1;
  assign or_dcpl_276 = ((in_data[199:180]==20'b00000000000000000000)) | (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_10_mx0[5]);
  assign or_dcpl_295 = (in_data[199:180]!=20'b00000000000000000000);
  assign and_dcpl_227 = or_dcpl_295 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_10_mx0[5]))
      & (~ operator_23_true_acc_9_itm_2_1);
  assign and_dcpl_229 = or_dcpl_295 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_10_mx0[5]))
      & operator_23_true_acc_9_itm_2_1;
  assign or_dcpl_296 = ((in_data[219:200]==20'b00000000000000000000)) | (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_11_mx0[5]);
  assign or_dcpl_315 = (in_data[219:200]!=20'b00000000000000000000);
  assign and_dcpl_250 = or_dcpl_315 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_11_mx0[5]))
      & (~ operator_23_true_acc_10_itm_2_1);
  assign and_dcpl_252 = or_dcpl_315 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_11_mx0[5]))
      & operator_23_true_acc_10_itm_2_1;
  assign or_dcpl_316 = ((in_data[239:220]==20'b00000000000000000000)) | (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_12_mx0[5]);
  assign or_dcpl_335 = (in_data[239:220]!=20'b00000000000000000000);
  assign and_dcpl_273 = or_dcpl_335 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_12_mx0[5]))
      & (~ operator_23_true_acc_11_itm_2_1);
  assign and_dcpl_275 = or_dcpl_335 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_12_mx0[5]))
      & operator_23_true_acc_11_itm_2_1;
  assign or_dcpl_336 = ((in_data[259:240]==20'b00000000000000000000)) | (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_13_mx0[5]);
  assign or_dcpl_355 = (in_data[259:240]!=20'b00000000000000000000);
  assign and_dcpl_296 = or_dcpl_355 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_13_mx0[5]))
      & (~ operator_23_true_acc_12_itm_2_1);
  assign and_dcpl_298 = or_dcpl_355 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_13_mx0[5]))
      & operator_23_true_acc_12_itm_2_1;
  assign or_dcpl_356 = ((in_data[279:260]==20'b00000000000000000000)) | (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_14_mx0[5]);
  assign or_dcpl_375 = (in_data[279:260]!=20'b00000000000000000000);
  assign and_dcpl_319 = or_dcpl_375 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_14_mx0[5]))
      & (~ operator_23_true_acc_13_itm_2_1);
  assign and_dcpl_321 = or_dcpl_375 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_14_mx0[5]))
      & operator_23_true_acc_13_itm_2_1;
  assign or_dcpl_376 = ((in_data[299:280]==20'b00000000000000000000)) | (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_15_mx0[5]);
  assign or_dcpl_395 = (in_data[299:280]!=20'b00000000000000000000);
  assign and_dcpl_342 = or_dcpl_395 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_15_mx0[5]))
      & (~ operator_23_true_acc_14_itm_2_1);
  assign and_dcpl_344 = or_dcpl_395 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_15_mx0[5]))
      & operator_23_true_acc_14_itm_2_1;
  assign or_dcpl_396 = ((in_data[319:300]==20'b00000000000000000000)) | (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_mx0[5]);
  assign or_dcpl_415 = (in_data[319:300]!=20'b00000000000000000000);
  assign and_dcpl_365 = or_dcpl_415 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_mx0[5]))
      & (~ operator_23_true_acc_15_itm_2_1);
  assign and_dcpl_367 = or_dcpl_415 & (~ (out_adpfloat_set_value_fixed_20U_14U_exp_tmp_5_0_mx0[5]))
      & operator_23_true_acc_15_itm_2_1;

  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_3_1_2;
    input [2:0] vector;
    reg [2:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_3_1_2 = tmp[0:0];
  end
  endfunction


  function automatic [5:0] conv_s2s_4_6 ;
    input [3:0]  vector ;
  begin
    conv_s2s_4_6 = {{2{vector[3]}}, vector};
  end
  endfunction


  function automatic [6:0] conv_s2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_s2u_6_7 = {vector[5], vector};
  end
  endfunction


  function automatic [5:0] conv_u2s_5_6 ;
    input [4:0]  vector ;
  begin
    conv_u2s_5_6 =  {1'b0, vector};
  end
  endfunction


  function automatic [6:0] conv_u2u_1_7 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_7 = {{6{1'b0}}, vector};
  end
  endfunction

endmodule




//------> ./ActUnit.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
// 
//  Generated by:   huaixil@sat8
//  Generated date: Fri Apr  8 23:14:40 2022
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_ActUnitRun_fsm
//  FSM Module
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_ActUnitRun_fsm (
  clk, rst, ActUnitRun_wen, fsm_output
);
  input clk;
  input rst;
  input ActUnitRun_wen;
  output [2:0] fsm_output;
  reg [2:0] fsm_output;


  // FSM State Type Declaration for ActUnit_ActUnit_ActUnitRun_ActUnitRun_fsm_1
  parameter
    ActUnitRun_rlp_C_0 = 2'd0,
    while_C_0 = 2'd1,
    while_C_1 = 2'd2;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : ActUnit_ActUnit_ActUnitRun_ActUnitRun_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 3'b010;
        state_var_NS = while_C_1;
      end
      while_C_1 : begin
        fsm_output = 3'b100;
        state_var_NS = while_C_0;
      end
      // ActUnitRun_rlp_C_0
      default : begin
        fsm_output = 3'b001;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk ) begin
    if ( ~ rst ) begin
      state_var <= ActUnitRun_rlp_C_0;
    end
    else if ( ActUnitRun_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_staller
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_staller (
  clk, rst, ActUnitRun_wen, ActUnitRun_wten, rva_out_Push_mioi_wen_comp, output_port_Push_mioi_wen_comp,
      done_Push_mioi_wen_comp
);
  input clk;
  input rst;
  output ActUnitRun_wen;
  output ActUnitRun_wten;
  input rva_out_Push_mioi_wen_comp;
  input output_port_Push_mioi_wen_comp;
  input done_Push_mioi_wen_comp;


  // Interconnect Declarations
  reg ActUnitRun_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign ActUnitRun_wen = rva_out_Push_mioi_wen_comp & output_port_Push_mioi_wen_comp
      & done_Push_mioi_wen_comp;
  assign ActUnitRun_wten = ActUnitRun_wten_reg;
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      ActUnitRun_wten_reg <= 1'b0;
    end
    else begin
      ActUnitRun_wten_reg <= ~ ActUnitRun_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_done_Push_mioi_done_Push_mio_wait_dp
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_done_Push_mioi_done_Push_mio_wait_dp (
  clk, rst, done_Push_mioi_oswt, done_Push_mioi_wen_comp, done_Push_mioi_biwt, done_Push_mioi_bdwt,
      done_Push_mioi_bcwt
);
  input clk;
  input rst;
  input done_Push_mioi_oswt;
  output done_Push_mioi_wen_comp;
  input done_Push_mioi_biwt;
  input done_Push_mioi_bdwt;
  output done_Push_mioi_bcwt;
  reg done_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign done_Push_mioi_wen_comp = (~ done_Push_mioi_oswt) | done_Push_mioi_biwt
      | done_Push_mioi_bcwt;
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      done_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      done_Push_mioi_bcwt <= ~((~(done_Push_mioi_bcwt | done_Push_mioi_biwt)) | done_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_done_Push_mioi_done_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_done_Push_mioi_done_Push_mio_wait_ctrl (
  ActUnitRun_wen, done_Push_mioi_oswt, done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct,
      done_Push_mioi_biwt, done_Push_mioi_bdwt, done_Push_mioi_bcwt, done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct,
      done_Push_mioi_ccs_ccore_done_sync_vld
);
  input ActUnitRun_wen;
  input done_Push_mioi_oswt;
  input done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct;
  output done_Push_mioi_biwt;
  output done_Push_mioi_bdwt;
  input done_Push_mioi_bcwt;
  output done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct;
  input done_Push_mioi_ccs_ccore_done_sync_vld;



  // Interconnect Declarations for Component Instantiations 
  assign done_Push_mioi_bdwt = done_Push_mioi_oswt & ActUnitRun_wen;
  assign done_Push_mioi_biwt = done_Push_mioi_oswt & (~ done_Push_mioi_bcwt) & done_Push_mioi_ccs_ccore_done_sync_vld;
  assign done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct = done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct
      & ActUnitRun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_output_port_Push_mioi_output_port_Push_mio_wait_dp
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_output_port_Push_mioi_output_port_Push_mio_wait_dp
    (
  clk, rst, output_port_Push_mioi_oswt, output_port_Push_mioi_wen_comp, output_port_Push_mioi_biwt,
      output_port_Push_mioi_bdwt, output_port_Push_mioi_bcwt
);
  input clk;
  input rst;
  input output_port_Push_mioi_oswt;
  output output_port_Push_mioi_wen_comp;
  input output_port_Push_mioi_biwt;
  input output_port_Push_mioi_bdwt;
  output output_port_Push_mioi_bcwt;
  reg output_port_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign output_port_Push_mioi_wen_comp = (~ output_port_Push_mioi_oswt) | output_port_Push_mioi_biwt
      | output_port_Push_mioi_bcwt;
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      output_port_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      output_port_Push_mioi_bcwt <= ~((~(output_port_Push_mioi_bcwt | output_port_Push_mioi_biwt))
          | output_port_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_output_port_Push_mioi_output_port_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_output_port_Push_mioi_output_port_Push_mio_wait_ctrl
    (
  ActUnitRun_wen, output_port_Push_mioi_oswt, output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct,
      output_port_Push_mioi_biwt, output_port_Push_mioi_bdwt, output_port_Push_mioi_bcwt,
      output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct, output_port_Push_mioi_ccs_ccore_done_sync_vld
);
  input ActUnitRun_wen;
  input output_port_Push_mioi_oswt;
  input output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct;
  output output_port_Push_mioi_biwt;
  output output_port_Push_mioi_bdwt;
  input output_port_Push_mioi_bcwt;
  output output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct;
  input output_port_Push_mioi_ccs_ccore_done_sync_vld;



  // Interconnect Declarations for Component Instantiations 
  assign output_port_Push_mioi_bdwt = output_port_Push_mioi_oswt & ActUnitRun_wen;
  assign output_port_Push_mioi_biwt = output_port_Push_mioi_oswt & (~ output_port_Push_mioi_bcwt)
      & output_port_Push_mioi_ccs_ccore_done_sync_vld;
  assign output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct = output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct
      & ActUnitRun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_start_PopNB_mioi_start_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_start_PopNB_mioi_start_PopNB_mio_wait_dp (
  clk, rst, start_PopNB_mioi_data_rsc_z_mxwt, start_PopNB_mioi_return_rsc_z_mxwt,
      start_PopNB_mioi_data_rsc_z, start_PopNB_mioi_biwt, start_PopNB_mioi_bdwt,
      start_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output start_PopNB_mioi_data_rsc_z_mxwt;
  output start_PopNB_mioi_return_rsc_z_mxwt;
  input start_PopNB_mioi_data_rsc_z;
  input start_PopNB_mioi_biwt;
  input start_PopNB_mioi_bdwt;
  input start_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg start_PopNB_mioi_bcwt;
  reg start_PopNB_mioi_data_rsc_z_bfwt;
  reg start_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign start_PopNB_mioi_data_rsc_z_mxwt = MUX_s_1_2_2(start_PopNB_mioi_data_rsc_z,
      start_PopNB_mioi_data_rsc_z_bfwt, start_PopNB_mioi_bcwt);
  assign start_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(start_PopNB_mioi_return_rsc_z,
      start_PopNB_mioi_return_rsc_z_bfwt, start_PopNB_mioi_bcwt);
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      start_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      start_PopNB_mioi_bcwt <= ~((~(start_PopNB_mioi_bcwt | start_PopNB_mioi_biwt))
          | start_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      start_PopNB_mioi_data_rsc_z_bfwt <= 1'b0;
      start_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( start_PopNB_mioi_biwt ) begin
      start_PopNB_mioi_data_rsc_z_bfwt <= start_PopNB_mioi_data_rsc_z;
      start_PopNB_mioi_return_rsc_z_bfwt <= start_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl (
  ActUnitRun_wen, ActUnitRun_wten, start_PopNB_mioi_oswt, start_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct,
      start_PopNB_mioi_biwt, start_PopNB_mioi_bdwt, start_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct
);
  input ActUnitRun_wen;
  input ActUnitRun_wten;
  input start_PopNB_mioi_oswt;
  input start_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct;
  output start_PopNB_mioi_biwt;
  output start_PopNB_mioi_bdwt;
  output start_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct;



  // Interconnect Declarations for Component Instantiations 
  assign start_PopNB_mioi_bdwt = start_PopNB_mioi_oswt & ActUnitRun_wen;
  assign start_PopNB_mioi_biwt = (~ ActUnitRun_wten) & start_PopNB_mioi_oswt;
  assign start_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct = start_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct
      & ActUnitRun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp (
  clk, rst, rva_out_Push_mioi_oswt, rva_out_Push_mioi_wen_comp, rva_out_Push_mioi_biwt,
      rva_out_Push_mioi_bdwt, rva_out_Push_mioi_bcwt
);
  input clk;
  input rst;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_wen_comp;
  input rva_out_Push_mioi_biwt;
  input rva_out_Push_mioi_bdwt;
  output rva_out_Push_mioi_bcwt;
  reg rva_out_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign rva_out_Push_mioi_wen_comp = (~ rva_out_Push_mioi_oswt) | rva_out_Push_mioi_biwt
      | rva_out_Push_mioi_bcwt;
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      rva_out_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      rva_out_Push_mioi_bcwt <= ~((~(rva_out_Push_mioi_bcwt | rva_out_Push_mioi_biwt))
          | rva_out_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl (
  ActUnitRun_wen, rva_out_Push_mioi_oswt, rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct,
      rva_out_Push_mioi_biwt, rva_out_Push_mioi_bdwt, rva_out_Push_mioi_bcwt, rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct,
      rva_out_Push_mioi_ccs_ccore_done_sync_vld
);
  input ActUnitRun_wen;
  input rva_out_Push_mioi_oswt;
  input rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct;
  output rva_out_Push_mioi_biwt;
  output rva_out_Push_mioi_bdwt;
  input rva_out_Push_mioi_bcwt;
  output rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct;
  input rva_out_Push_mioi_ccs_ccore_done_sync_vld;



  // Interconnect Declarations for Component Instantiations 
  assign rva_out_Push_mioi_bdwt = rva_out_Push_mioi_oswt & ActUnitRun_wen;
  assign rva_out_Push_mioi_biwt = rva_out_Push_mioi_oswt & (~ rva_out_Push_mioi_bcwt)
      & rva_out_Push_mioi_ccs_ccore_done_sync_vld;
  assign rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct = rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct
      & ActUnitRun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_act_port_PopNB_mioi_act_port_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_act_port_PopNB_mioi_act_port_PopNB_mio_wait_dp
    (
  clk, rst, act_port_PopNB_mioi_data_data_rsc_z_mxwt, act_port_PopNB_mioi_return_rsc_z_mxwt,
      act_port_PopNB_mioi_data_data_rsc_z, act_port_PopNB_mioi_biwt, act_port_PopNB_mioi_bdwt,
      act_port_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [319:0] act_port_PopNB_mioi_data_data_rsc_z_mxwt;
  output act_port_PopNB_mioi_return_rsc_z_mxwt;
  input [319:0] act_port_PopNB_mioi_data_data_rsc_z;
  input act_port_PopNB_mioi_biwt;
  input act_port_PopNB_mioi_bdwt;
  input act_port_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg act_port_PopNB_mioi_bcwt;
  reg [319:0] act_port_PopNB_mioi_data_data_rsc_z_bfwt;
  reg act_port_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign act_port_PopNB_mioi_data_data_rsc_z_mxwt = MUX_v_320_2_2(act_port_PopNB_mioi_data_data_rsc_z,
      act_port_PopNB_mioi_data_data_rsc_z_bfwt, act_port_PopNB_mioi_bcwt);
  assign act_port_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(act_port_PopNB_mioi_return_rsc_z,
      act_port_PopNB_mioi_return_rsc_z_bfwt, act_port_PopNB_mioi_bcwt);
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_port_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      act_port_PopNB_mioi_bcwt <= ~((~(act_port_PopNB_mioi_bcwt | act_port_PopNB_mioi_biwt))
          | act_port_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_port_PopNB_mioi_data_data_rsc_z_bfwt <= 320'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      act_port_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( act_port_PopNB_mioi_biwt ) begin
      act_port_PopNB_mioi_data_data_rsc_z_bfwt <= act_port_PopNB_mioi_data_data_rsc_z;
      act_port_PopNB_mioi_return_rsc_z_bfwt <= act_port_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [319:0] MUX_v_320_2_2;
    input [319:0] input_0;
    input [319:0] input_1;
    input [0:0] sel;
    reg [319:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_320_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_act_port_PopNB_mioi_act_port_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_act_port_PopNB_mioi_act_port_PopNB_mio_wait_ctrl
    (
  ActUnitRun_wen, ActUnitRun_wten, act_port_PopNB_mioi_oswt, act_port_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct,
      act_port_PopNB_mioi_biwt, act_port_PopNB_mioi_bdwt, act_port_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct
);
  input ActUnitRun_wen;
  input ActUnitRun_wten;
  input act_port_PopNB_mioi_oswt;
  input act_port_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct;
  output act_port_PopNB_mioi_biwt;
  output act_port_PopNB_mioi_bdwt;
  output act_port_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct;



  // Interconnect Declarations for Component Instantiations 
  assign act_port_PopNB_mioi_bdwt = act_port_PopNB_mioi_oswt & ActUnitRun_wen;
  assign act_port_PopNB_mioi_biwt = (~ ActUnitRun_wten) & act_port_PopNB_mioi_oswt;
  assign act_port_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct = act_port_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct
      & ActUnitRun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp (
  clk, rst, rva_in_PopNB_mioi_data_data_rsc_z_mxwt, rva_in_PopNB_mioi_data_addr_rsc_z_mxwt,
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt, rva_in_PopNB_mioi_return_rsc_z_mxwt,
      rva_in_PopNB_mioi_data_data_rsc_z, rva_in_PopNB_mioi_biwt, rva_in_PopNB_mioi_bdwt,
      rva_in_PopNB_mioi_data_addr_rsc_z, rva_in_PopNB_mioi_data_rw_rsc_z, rva_in_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [127:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  output [11:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  output rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  output rva_in_PopNB_mioi_return_rsc_z_mxwt;
  input [127:0] rva_in_PopNB_mioi_data_data_rsc_z;
  input rva_in_PopNB_mioi_biwt;
  input rva_in_PopNB_mioi_bdwt;
  input [23:0] rva_in_PopNB_mioi_data_addr_rsc_z;
  input rva_in_PopNB_mioi_data_rw_rsc_z;
  input rva_in_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg rva_in_PopNB_mioi_bcwt;
  reg [127:0] rva_in_PopNB_mioi_data_data_rsc_z_bfwt;
  reg rva_in_PopNB_mioi_data_rw_rsc_z_bfwt;
  reg rva_in_PopNB_mioi_return_rsc_z_bfwt;
  wire [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst;
  reg [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4;


  // Interconnect Declarations for Component Instantiations 
  assign rva_in_PopNB_mioi_data_data_rsc_z_mxwt = MUX_v_128_2_2(rva_in_PopNB_mioi_data_data_rsc_z,
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_data_rw_rsc_z_mxwt = MUX_s_1_2_2(rva_in_PopNB_mioi_data_rw_rsc_z,
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(rva_in_PopNB_mioi_return_rsc_z,
      rva_in_PopNB_mioi_return_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst = MUX_v_20_2_2((rva_in_PopNB_mioi_data_addr_rsc_z[23:4]),
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_data_addr_rsc_z_mxwt = {(rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst[19:16])
      , (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst[7:0])};
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      rva_in_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      rva_in_PopNB_mioi_bcwt <= ~((~(rva_in_PopNB_mioi_bcwt | rva_in_PopNB_mioi_biwt))
          | rva_in_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4 <= 20'b00000000000000000000;
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt <= 1'b0;
      rva_in_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( rva_in_PopNB_mioi_biwt ) begin
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt <= rva_in_PopNB_mioi_data_data_rsc_z;
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4 <= rva_in_PopNB_mioi_data_addr_rsc_z[23:4];
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt <= rva_in_PopNB_mioi_data_rw_rsc_z;
      rva_in_PopNB_mioi_return_rsc_z_bfwt <= rva_in_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input [0:0] sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction


  function automatic [19:0] MUX_v_20_2_2;
    input [19:0] input_0;
    input [19:0] input_1;
    input [0:0] sel;
    reg [19:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_20_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl (
  ActUnitRun_wen, rva_in_PopNB_mioi_oswt, ActUnitRun_wten, rva_in_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct,
      rva_in_PopNB_mioi_biwt, rva_in_PopNB_mioi_bdwt, rva_in_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct
);
  input ActUnitRun_wen;
  input rva_in_PopNB_mioi_oswt;
  input ActUnitRun_wten;
  input rva_in_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct;
  output rva_in_PopNB_mioi_biwt;
  output rva_in_PopNB_mioi_bdwt;
  output rva_in_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct;



  // Interconnect Declarations for Component Instantiations 
  assign rva_in_PopNB_mioi_bdwt = rva_in_PopNB_mioi_oswt & ActUnitRun_wen;
  assign rva_in_PopNB_mioi_biwt = (~ ActUnitRun_wten) & rva_in_PopNB_mioi_oswt;
  assign rva_in_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct = rva_in_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct
      & ActUnitRun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_done_Push_mioi
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_done_Push_mioi (
  clk, rst, done_val, done_rdy, done_msg, ActUnitRun_wen, done_Push_mioi_oswt, done_Push_mioi_wen_comp,
      done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct
);
  input clk;
  input rst;
  output done_val;
  input done_rdy;
  output done_msg;
  input ActUnitRun_wen;
  input done_Push_mioi_oswt;
  output done_Push_mioi_wen_comp;
  input done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct;


  // Interconnect Declarations
  wire done_Push_mioi_biwt;
  wire done_Push_mioi_bdwt;
  wire done_Push_mioi_bcwt;
  wire done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct;
  wire done_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  ActUnit_Connections_OutBlocking_bool_Connections_SYN_PORT_Push  done_Push_mioi
      (
      .this_val(done_val),
      .this_rdy(done_rdy),
      .this_msg(done_msg),
      .ccs_ccore_start_rsc_dat(done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct),
      .ccs_ccore_done_sync_vld(done_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  ActUnit_ActUnit_ActUnitRun_done_Push_mioi_done_Push_mio_wait_ctrl ActUnit_ActUnitRun_done_Push_mioi_done_Push_mio_wait_ctrl_inst
      (
      .ActUnitRun_wen(ActUnitRun_wen),
      .done_Push_mioi_oswt(done_Push_mioi_oswt),
      .done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct(done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct),
      .done_Push_mioi_biwt(done_Push_mioi_biwt),
      .done_Push_mioi_bdwt(done_Push_mioi_bdwt),
      .done_Push_mioi_bcwt(done_Push_mioi_bcwt),
      .done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct(done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct),
      .done_Push_mioi_ccs_ccore_done_sync_vld(done_Push_mioi_ccs_ccore_done_sync_vld)
    );
  ActUnit_ActUnit_ActUnitRun_done_Push_mioi_done_Push_mio_wait_dp ActUnit_ActUnitRun_done_Push_mioi_done_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .done_Push_mioi_oswt(done_Push_mioi_oswt),
      .done_Push_mioi_wen_comp(done_Push_mioi_wen_comp),
      .done_Push_mioi_biwt(done_Push_mioi_biwt),
      .done_Push_mioi_bdwt(done_Push_mioi_bdwt),
      .done_Push_mioi_bcwt(done_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_output_port_Push_mioi
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_output_port_Push_mioi (
  clk, rst, output_port_val, output_port_rdy, output_port_msg, ActUnitRun_wen, output_port_Push_mioi_oswt,
      output_port_Push_mioi_wen_comp, output_port_Push_mioi_m_data_data_rsc_dat_ActUnitRun,
      output_port_Push_mioi_m_logical_addr_rsc_dat_ActUnitRun, output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct
);
  input clk;
  input rst;
  output output_port_val;
  input output_port_rdy;
  output [137:0] output_port_msg;
  input ActUnitRun_wen;
  input output_port_Push_mioi_oswt;
  output output_port_Push_mioi_wen_comp;
  input [127:0] output_port_Push_mioi_m_data_data_rsc_dat_ActUnitRun;
  input [7:0] output_port_Push_mioi_m_logical_addr_rsc_dat_ActUnitRun;
  input output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct;


  // Interconnect Declarations
  wire output_port_Push_mioi_biwt;
  wire output_port_Push_mioi_bdwt;
  wire output_port_Push_mioi_bcwt;
  wire output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct;
  wire output_port_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  ActUnit_Connections_OutBlocking_spec_StreamType_Connections_SYN_PORT_Push  output_port_Push_mioi
      (
      .this_val(output_port_val),
      .this_rdy(output_port_rdy),
      .this_msg(output_port_msg),
      .m_data_data_rsc_dat(output_port_Push_mioi_m_data_data_rsc_dat_ActUnitRun),
      .m_logical_addr_rsc_dat(output_port_Push_mioi_m_logical_addr_rsc_dat_ActUnitRun),
      .ccs_ccore_start_rsc_dat(output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct),
      .ccs_ccore_done_sync_vld(output_port_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  ActUnit_ActUnit_ActUnitRun_output_port_Push_mioi_output_port_Push_mio_wait_ctrl
      ActUnit_ActUnitRun_output_port_Push_mioi_output_port_Push_mio_wait_ctrl_inst
      (
      .ActUnitRun_wen(ActUnitRun_wen),
      .output_port_Push_mioi_oswt(output_port_Push_mioi_oswt),
      .output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct(output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct),
      .output_port_Push_mioi_biwt(output_port_Push_mioi_biwt),
      .output_port_Push_mioi_bdwt(output_port_Push_mioi_bdwt),
      .output_port_Push_mioi_bcwt(output_port_Push_mioi_bcwt),
      .output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct(output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct),
      .output_port_Push_mioi_ccs_ccore_done_sync_vld(output_port_Push_mioi_ccs_ccore_done_sync_vld)
    );
  ActUnit_ActUnit_ActUnitRun_output_port_Push_mioi_output_port_Push_mio_wait_dp ActUnit_ActUnitRun_output_port_Push_mioi_output_port_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .output_port_Push_mioi_oswt(output_port_Push_mioi_oswt),
      .output_port_Push_mioi_wen_comp(output_port_Push_mioi_wen_comp),
      .output_port_Push_mioi_biwt(output_port_Push_mioi_biwt),
      .output_port_Push_mioi_bdwt(output_port_Push_mioi_bdwt),
      .output_port_Push_mioi_bcwt(output_port_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_start_PopNB_mioi
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_start_PopNB_mioi (
  clk, rst, start_val, start_rdy, start_msg, ActUnitRun_wen, ActUnitRun_wten, start_PopNB_mioi_oswt,
      start_PopNB_mioi_data_rsc_z_mxwt, start_PopNB_mioi_return_rsc_z_mxwt, start_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct
);
  input clk;
  input rst;
  input start_val;
  output start_rdy;
  input start_msg;
  input ActUnitRun_wen;
  input ActUnitRun_wten;
  input start_PopNB_mioi_oswt;
  output start_PopNB_mioi_data_rsc_z_mxwt;
  output start_PopNB_mioi_return_rsc_z_mxwt;
  input start_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct;


  // Interconnect Declarations
  wire start_PopNB_mioi_data_rsc_z;
  wire start_PopNB_mioi_biwt;
  wire start_PopNB_mioi_bdwt;
  wire start_PopNB_mioi_return_rsc_z;
  wire start_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct;


  // Interconnect Declarations for Component Instantiations 
  ActUnit_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB  start_PopNB_mioi
      (
      .this_val(start_val),
      .this_rdy(start_rdy),
      .this_msg(start_msg),
      .data_rsc_z(start_PopNB_mioi_data_rsc_z),
      .return_rsc_z(start_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(start_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  ActUnit_ActUnit_ActUnitRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl ActUnit_ActUnitRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl_inst
      (
      .ActUnitRun_wen(ActUnitRun_wen),
      .ActUnitRun_wten(ActUnitRun_wten),
      .start_PopNB_mioi_oswt(start_PopNB_mioi_oswt),
      .start_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct(start_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct),
      .start_PopNB_mioi_biwt(start_PopNB_mioi_biwt),
      .start_PopNB_mioi_bdwt(start_PopNB_mioi_bdwt),
      .start_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct(start_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct)
    );
  ActUnit_ActUnit_ActUnitRun_start_PopNB_mioi_start_PopNB_mio_wait_dp ActUnit_ActUnitRun_start_PopNB_mioi_start_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .start_PopNB_mioi_data_rsc_z_mxwt(start_PopNB_mioi_data_rsc_z_mxwt),
      .start_PopNB_mioi_return_rsc_z_mxwt(start_PopNB_mioi_return_rsc_z_mxwt),
      .start_PopNB_mioi_data_rsc_z(start_PopNB_mioi_data_rsc_z),
      .start_PopNB_mioi_biwt(start_PopNB_mioi_biwt),
      .start_PopNB_mioi_bdwt(start_PopNB_mioi_bdwt),
      .start_PopNB_mioi_return_rsc_z(start_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_rva_out_Push_mioi
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_rva_out_Push_mioi (
  clk, rst, rva_out_val, rva_out_rdy, rva_out_msg, ActUnitRun_wen, rva_out_Push_mioi_oswt,
      rva_out_Push_mioi_wen_comp, rva_out_Push_mioi_m_data_rsc_dat_ActUnitRun, rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct
);
  input clk;
  input rst;
  output rva_out_val;
  input rva_out_rdy;
  output [127:0] rva_out_msg;
  input ActUnitRun_wen;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_wen_comp;
  input [127:0] rva_out_Push_mioi_m_data_rsc_dat_ActUnitRun;
  input rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct;


  // Interconnect Declarations
  wire rva_out_Push_mioi_biwt;
  wire rva_out_Push_mioi_bdwt;
  wire rva_out_Push_mioi_bcwt;
  wire rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct;
  wire rva_out_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  ActUnit_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
      rva_out_Push_mioi (
      .this_val(rva_out_val),
      .this_rdy(rva_out_rdy),
      .this_msg(rva_out_msg),
      .m_data_rsc_dat(rva_out_Push_mioi_m_data_rsc_dat_ActUnitRun),
      .ccs_ccore_start_rsc_dat(rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct),
      .ccs_ccore_done_sync_vld(rva_out_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  ActUnit_ActUnit_ActUnitRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl ActUnit_ActUnitRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl_inst
      (
      .ActUnitRun_wen(ActUnitRun_wen),
      .rva_out_Push_mioi_oswt(rva_out_Push_mioi_oswt),
      .rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct(rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct),
      .rva_out_Push_mioi_biwt(rva_out_Push_mioi_biwt),
      .rva_out_Push_mioi_bdwt(rva_out_Push_mioi_bdwt),
      .rva_out_Push_mioi_bcwt(rva_out_Push_mioi_bcwt),
      .rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct(rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct),
      .rva_out_Push_mioi_ccs_ccore_done_sync_vld(rva_out_Push_mioi_ccs_ccore_done_sync_vld)
    );
  ActUnit_ActUnit_ActUnitRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp ActUnit_ActUnitRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_out_Push_mioi_oswt(rva_out_Push_mioi_oswt),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp),
      .rva_out_Push_mioi_biwt(rva_out_Push_mioi_biwt),
      .rva_out_Push_mioi_bdwt(rva_out_Push_mioi_bdwt),
      .rva_out_Push_mioi_bcwt(rva_out_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_act_port_PopNB_mioi
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_act_port_PopNB_mioi (
  clk, rst, act_port_val, act_port_rdy, act_port_msg, ActUnitRun_wen, ActUnitRun_wten,
      act_port_PopNB_mioi_oswt, act_port_PopNB_mioi_data_data_rsc_z_mxwt, act_port_PopNB_mioi_return_rsc_z_mxwt,
      act_port_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct
);
  input clk;
  input rst;
  input act_port_val;
  output act_port_rdy;
  input [319:0] act_port_msg;
  input ActUnitRun_wen;
  input ActUnitRun_wten;
  input act_port_PopNB_mioi_oswt;
  output [319:0] act_port_PopNB_mioi_data_data_rsc_z_mxwt;
  output act_port_PopNB_mioi_return_rsc_z_mxwt;
  input act_port_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct;


  // Interconnect Declarations
  wire [319:0] act_port_PopNB_mioi_data_data_rsc_z;
  wire act_port_PopNB_mioi_biwt;
  wire act_port_PopNB_mioi_bdwt;
  wire act_port_PopNB_mioi_return_rsc_z;
  wire act_port_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct;


  // Interconnect Declarations for Component Instantiations 
  ActUnit_Connections_InBlocking_spec_ActVectorType_Connections_SYN_PORT_PopNB  act_port_PopNB_mioi
      (
      .this_val(act_port_val),
      .this_rdy(act_port_rdy),
      .this_msg(act_port_msg),
      .data_data_rsc_z(act_port_PopNB_mioi_data_data_rsc_z),
      .return_rsc_z(act_port_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(act_port_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  ActUnit_ActUnit_ActUnitRun_act_port_PopNB_mioi_act_port_PopNB_mio_wait_ctrl ActUnit_ActUnitRun_act_port_PopNB_mioi_act_port_PopNB_mio_wait_ctrl_inst
      (
      .ActUnitRun_wen(ActUnitRun_wen),
      .ActUnitRun_wten(ActUnitRun_wten),
      .act_port_PopNB_mioi_oswt(act_port_PopNB_mioi_oswt),
      .act_port_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct(act_port_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct),
      .act_port_PopNB_mioi_biwt(act_port_PopNB_mioi_biwt),
      .act_port_PopNB_mioi_bdwt(act_port_PopNB_mioi_bdwt),
      .act_port_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct(act_port_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct)
    );
  ActUnit_ActUnit_ActUnitRun_act_port_PopNB_mioi_act_port_PopNB_mio_wait_dp ActUnit_ActUnitRun_act_port_PopNB_mioi_act_port_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .act_port_PopNB_mioi_data_data_rsc_z_mxwt(act_port_PopNB_mioi_data_data_rsc_z_mxwt),
      .act_port_PopNB_mioi_return_rsc_z_mxwt(act_port_PopNB_mioi_return_rsc_z_mxwt),
      .act_port_PopNB_mioi_data_data_rsc_z(act_port_PopNB_mioi_data_data_rsc_z),
      .act_port_PopNB_mioi_biwt(act_port_PopNB_mioi_biwt),
      .act_port_PopNB_mioi_bdwt(act_port_PopNB_mioi_bdwt),
      .act_port_PopNB_mioi_return_rsc_z(act_port_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_rva_in_PopNB_mioi
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_rva_in_PopNB_mioi (
  clk, rst, rva_in_val, rva_in_rdy, rva_in_msg, ActUnitRun_wen, rva_in_PopNB_mioi_oswt,
      ActUnitRun_wten, rva_in_PopNB_mioi_data_data_rsc_z_mxwt, rva_in_PopNB_mioi_data_addr_rsc_z_mxwt,
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt, rva_in_PopNB_mioi_return_rsc_z_mxwt,
      rva_in_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct
);
  input clk;
  input rst;
  input rva_in_val;
  output rva_in_rdy;
  input [168:0] rva_in_msg;
  input ActUnitRun_wen;
  input rva_in_PopNB_mioi_oswt;
  input ActUnitRun_wten;
  output [127:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  output [11:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  output rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  output rva_in_PopNB_mioi_return_rsc_z_mxwt;
  input rva_in_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct;


  // Interconnect Declarations
  wire [127:0] rva_in_PopNB_mioi_data_data_rsc_z;
  wire rva_in_PopNB_mioi_biwt;
  wire rva_in_PopNB_mioi_bdwt;
  wire [23:0] rva_in_PopNB_mioi_data_addr_rsc_z;
  wire [15:0] rva_in_PopNB_mioi_data_wstrb_rsc_z;
  wire rva_in_PopNB_mioi_data_rw_rsc_z;
  wire rva_in_PopNB_mioi_return_rsc_z;
  wire rva_in_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct;
  wire [11:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  ActUnit_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
      rva_in_PopNB_mioi (
      .this_val(rva_in_val),
      .this_rdy(rva_in_rdy),
      .this_msg(rva_in_msg),
      .data_data_rsc_z(rva_in_PopNB_mioi_data_data_rsc_z),
      .data_addr_rsc_z(rva_in_PopNB_mioi_data_addr_rsc_z),
      .data_wstrb_rsc_z(rva_in_PopNB_mioi_data_wstrb_rsc_z),
      .data_rw_rsc_z(rva_in_PopNB_mioi_data_rw_rsc_z),
      .return_rsc_z(rva_in_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(rva_in_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  ActUnit_ActUnit_ActUnitRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl ActUnit_ActUnitRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl_inst
      (
      .ActUnitRun_wen(ActUnitRun_wen),
      .rva_in_PopNB_mioi_oswt(rva_in_PopNB_mioi_oswt),
      .ActUnitRun_wten(ActUnitRun_wten),
      .rva_in_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct(rva_in_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct),
      .rva_in_PopNB_mioi_biwt(rva_in_PopNB_mioi_biwt),
      .rva_in_PopNB_mioi_bdwt(rva_in_PopNB_mioi_bdwt),
      .rva_in_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct(rva_in_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct)
    );
  ActUnit_ActUnit_ActUnitRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp ActUnit_ActUnitRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_in_PopNB_mioi_data_data_rsc_z_mxwt(rva_in_PopNB_mioi_data_data_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_addr_rsc_z_mxwt(rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst),
      .rva_in_PopNB_mioi_data_rw_rsc_z_mxwt(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt),
      .rva_in_PopNB_mioi_return_rsc_z_mxwt(rva_in_PopNB_mioi_return_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_data_rsc_z(rva_in_PopNB_mioi_data_data_rsc_z),
      .rva_in_PopNB_mioi_biwt(rva_in_PopNB_mioi_biwt),
      .rva_in_PopNB_mioi_bdwt(rva_in_PopNB_mioi_bdwt),
      .rva_in_PopNB_mioi_data_addr_rsc_z(rva_in_PopNB_mioi_data_addr_rsc_z),
      .rva_in_PopNB_mioi_data_rw_rsc_z(rva_in_PopNB_mioi_data_rw_rsc_z),
      .rva_in_PopNB_mioi_return_rsc_z(rva_in_PopNB_mioi_return_rsc_z)
    );
  assign rva_in_PopNB_mioi_data_addr_rsc_z_mxwt = rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun (
  clk, rst, start_val, start_rdy, start_msg, act_port_val, act_port_rdy, act_port_msg,
      rva_in_val, rva_in_rdy, rva_in_msg, rva_out_val, rva_out_rdy, rva_out_msg,
      output_port_val, output_port_rdy, output_port_msg, done_val, done_rdy, done_msg
);
  input clk;
  input rst;
  input start_val;
  output start_rdy;
  input start_msg;
  input act_port_val;
  output act_port_rdy;
  input [319:0] act_port_msg;
  input rva_in_val;
  output rva_in_rdy;
  input [168:0] rva_in_msg;
  output rva_out_val;
  input rva_out_rdy;
  output [127:0] rva_out_msg;
  output output_port_val;
  input output_port_rdy;
  output [137:0] output_port_msg;
  output done_val;
  input done_rdy;
  output done_msg;


  // Interconnect Declarations
  wire ActUnitRun_wen;
  wire ActUnitRun_wten;
  wire [127:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  wire [11:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  wire rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  wire rva_in_PopNB_mioi_return_rsc_z_mxwt;
  wire [319:0] act_port_PopNB_mioi_data_data_rsc_z_mxwt;
  wire act_port_PopNB_mioi_return_rsc_z_mxwt;
  wire rva_out_Push_mioi_wen_comp;
  wire start_PopNB_mioi_data_rsc_z_mxwt;
  wire start_PopNB_mioi_return_rsc_z_mxwt;
  wire output_port_Push_mioi_wen_comp;
  wire done_Push_mioi_wen_comp;
  wire [2:0] fsm_output;
  wire act_config_InstIncr_if_if_unequal_tmp;
  wire [8:0] operator_8_false_acc_tmp;
  wire [9:0] nl_operator_8_false_acc_tmp;
  wire act_config_InstIncr_if_equal_1_tmp;
  wire [6:0] operator_6_false_acc_tmp;
  wire [7:0] nl_operator_6_false_acc_tmp;
  wire ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_1_tmp;
  wire [7:0] act_config_in_InstFetch_mux_tmp;
  wire [4:0] while_mux_125_tmp;
  wire mux_tmp_1;
  wire and_dcpl;
  wire and_dcpl_1;
  wire and_dcpl_5;
  wire and_dcpl_8;
  wire and_dcpl_11;
  wire or_dcpl_8;
  wire or_dcpl_9;
  wire and_dcpl_31;
  wire nor_tmp_6;
  wire mux_tmp_16;
  wire or_dcpl_13;
  wire or_dcpl_15;
  wire or_dcpl_22;
  wire not_tmp_34;
  wire or_dcpl_27;
  wire and_dcpl_45;
  wire or_dcpl_33;
  wire or_dcpl_34;
  wire or_dcpl_35;
  wire or_dcpl_38;
  wire or_dcpl_41;
  wire or_dcpl_44;
  wire or_dcpl_47;
  wire or_dcpl_56;
  wire or_dcpl_57;
  wire or_dcpl_66;
  wire or_dcpl_75;
  wire or_dcpl_76;
  wire or_dcpl_85;
  wire or_dcpl_94;
  wire or_dcpl_95;
  wire or_dcpl_104;
  wire or_dcpl_116;
  wire and_dcpl_65;
  wire or_tmp_61;
  wire and_158_cse;
  wire act_config_InstIncr_if_act_config_InstIncr_if_if_act_config_InstIncr_if_if_nor_mdf_sva_1;
  wire act_config_InstIncr_act_config_InstIncr_if_and_svs_1;
  wire act_config_ActConfigRead_else_unequal_tmp_1;
  wire act_config_ActConfigRead_unequal_tmp_1;
  wire ActUnit_RunInst_switch_lp_and_66_tmp_1;
  reg ActUnit_RunInst_switch_lp_equal_tmp_2;
  reg is_start_sva;
  wire ActUnit_RunInst_switch_lp_equal_tmp_20;
  reg ActUnit_RunInst_switch_lp_equal_tmp_1;
  reg ActUnit_RunInst_switch_lp_equal_tmp_3;
  reg ActUnit_RunInst_switch_lp_nor_tmp;
  reg ActUnit_RunInst_switch_lp_equal_tmp_4;
  reg ActUnit_RunInst_switch_lp_equal_tmp_5;
  reg ActUnit_RunInst_switch_lp_equal_tmp_6;
  reg ActUnit_RunInst_switch_lp_equal_tmp_7;
  reg ActUnit_RunInst_switch_lp_equal_tmp_8;
  reg ActUnit_RunInst_switch_lp_equal_tmp_9;
  reg ActUnit_RunInst_switch_lp_equal_tmp_10;
  wire ActUnit_RunInst_switch_lp_and_ssc_sva_1;
  wire ActUnit_RunInst_switch_lp_and_50_tmp_1;
  wire ActUnit_RunInst_switch_lp_and_ssc_1_sva_1;
  wire ActUnit_RunInst_switch_lp_and_34_tmp_1;
  wire ActUnit_RunInst_switch_lp_and_ssc_2_sva_1;
  wire ActUnit_RunInst_switch_lp_and_18_tmp_1;
  wire ActUnit_RunInst_switch_lp_nor_ssc_sva_1;
  wire ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0;
  wire ActUnit_RunInst_switch_lp_equal_tmp_11;
  wire ActUnit_RunInst_switch_lp_equal_tmp_12;
  wire ActUnit_RunInst_switch_lp_equal_tmp_13;
  wire ActUnit_RunInst_switch_lp_equal_tmp_14;
  wire ActUnit_RunInst_switch_lp_equal_tmp_15;
  wire ActUnit_RunInst_switch_lp_equal_tmp_16;
  wire ActUnit_RunInst_switch_lp_equal_tmp_17;
  wire ActUnit_RunInst_switch_lp_equal_tmp_18;
  wire ActUnit_RunInst_switch_lp_equal_tmp_19;
  wire ActUnit_RunInst_switch_lp_nor_tmp_1;
  wire is_incr_lpi_1_dfm_2;
  wire ActUnit_RunLoad_if_else_and_ssc_sva_1;
  wire ActUnit_PushOutput_and_tmp_1;
  wire act_config_is_zero_first_sva_dfm_4_mx0;
  wire ActUnit_RunLoad_if_else_and_ssc_1_sva_1;
  wire ActUnit_RunLoad_if_else_and_ssc_2_sva_1;
  wire ActUnit_RunLoad_if_else_nor_ssc_sva_1;
  reg ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_cse;
  reg [4:0] act_config_inst_counter_sva;
  wire [7:0] ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_23_4_mx1_tmp_7_0;
  reg act_config_is_valid_sva;
  wire ActUnit_DecodeAxiRead_unequal_tmp_1;
  wire [1:0] nvhls_get_slc_2U_NVUINT8_return_3_sva_1;
  reg [7:0] act_config_inst_regs_0_sva_dfm_5;
  reg [7:0] act_config_inst_regs_1_sva_dfm_5;
  reg [7:0] act_config_inst_regs_2_sva_dfm_5;
  reg [7:0] act_config_inst_regs_3_sva_dfm_5;
  reg [7:0] act_config_inst_regs_4_sva_dfm_5;
  reg [7:0] act_config_inst_regs_5_sva_dfm_5;
  reg [7:0] act_config_inst_regs_6_sva_dfm_5;
  reg [7:0] act_config_inst_regs_7_sva_dfm_5;
  reg [7:0] act_config_inst_regs_8_sva_dfm_5;
  reg [7:0] act_config_inst_regs_9_sva_dfm_5;
  reg [7:0] act_config_inst_regs_10_sva_dfm_5;
  reg [7:0] act_config_inst_regs_11_sva_dfm_5;
  reg [7:0] act_config_inst_regs_12_sva_dfm_5;
  reg [7:0] act_config_inst_regs_13_sva_dfm_5;
  reg [7:0] act_config_inst_regs_14_sva_dfm_5;
  reg [7:0] act_config_inst_regs_15_sva_dfm_5;
  reg [7:0] act_config_inst_regs_16_sva_dfm_6;
  reg [7:0] act_config_inst_regs_17_sva_dfm_6;
  reg [7:0] act_config_inst_regs_18_sva_dfm_6;
  reg [7:0] act_config_inst_regs_19_sva_dfm_6;
  reg [7:0] act_config_inst_regs_20_sva_dfm_6;
  reg [7:0] act_config_inst_regs_21_sva_dfm_6;
  reg [7:0] act_config_inst_regs_22_sva_dfm_6;
  reg [7:0] act_config_inst_regs_23_sva_dfm_6;
  reg [7:0] act_config_inst_regs_24_sva_dfm_6;
  reg [7:0] act_config_inst_regs_25_sva_dfm_6;
  reg [7:0] act_config_inst_regs_26_sva_dfm_6;
  reg [7:0] act_config_inst_regs_27_sva_dfm_6;
  reg [7:0] act_config_inst_regs_28_sva_dfm_6;
  reg [7:0] act_config_inst_regs_29_sva_dfm_6;
  reg [7:0] act_config_inst_regs_30_sva_dfm_6;
  reg [7:0] act_config_inst_regs_31_sva_dfm_6;
  reg [7:0] reg_ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_23_4_ftd_12;
  wire act_mem_banks_write_if_for_if_mux_cse;
  wire act_mem_banks_write_if_for_if_mux_1_cse;
  wire act_mem_banks_read_for_mux_16_cse;
  wire act_mem_banks_read_for_mux_17_cse;
  wire ActUnit_DecodeAxiRead_and_9_cse;
  wire ActUnit_DecodeAxiRead_and_10_cse;
  reg reg_done_Push_mioi_iswt0_cse;
  reg reg_output_port_Push_mioi_iswt0_cse;
  reg reg_start_PopNB_mioi_iswt0_cse;
  reg reg_rva_out_Push_mioi_iswt0_cse;
  reg reg_act_port_PopNB_mioi_iswt0_cse;
  reg reg_rva_in_PopNB_mioi_iswt0_cse;
  wire act_regs_data_and_cse;
  wire act_config_adpfloat_bias_and_cse;
  wire act_config_inst_regs_and_cse;
  wire act_config_inst_regs_and_16_cse;
  wire act_mem_banks_bank_array_impl_data0_and_cse;
  wire act_mem_banks_bank_array_impl_data0_and_1_cse;
  wire act_mem_banks_bank_array_impl_data0_and_2_cse;
  wire act_mem_banks_bank_array_impl_data0_and_3_cse;
  wire act_mem_banks_bank_array_impl_data0_and_4_cse;
  wire act_mem_banks_bank_array_impl_data0_and_5_cse;
  wire act_mem_banks_bank_array_impl_data0_and_6_cse;
  wire act_mem_banks_bank_array_impl_data0_and_7_cse;
  wire act_mem_banks_bank_array_impl_data0_and_8_cse;
  wire act_mem_banks_bank_array_impl_data0_and_9_cse;
  wire act_mem_banks_bank_array_impl_data0_and_10_cse;
  wire act_mem_banks_bank_array_impl_data0_and_11_cse;
  wire act_mem_banks_bank_array_impl_data0_and_12_cse;
  wire act_mem_banks_bank_array_impl_data0_and_13_cse;
  wire act_mem_banks_bank_array_impl_data0_and_14_cse;
  wire act_mem_banks_bank_array_impl_data0_and_15_cse;
  wire act_mem_banks_bank_array_impl_data0_and_16_cse;
  wire act_mem_banks_bank_array_impl_data0_and_17_cse;
  wire act_mem_banks_bank_array_impl_data0_and_18_cse;
  wire act_mem_banks_bank_array_impl_data0_and_19_cse;
  wire act_mem_banks_bank_array_impl_data0_and_20_cse;
  wire act_mem_banks_bank_array_impl_data0_and_21_cse;
  wire act_mem_banks_bank_array_impl_data0_and_22_cse;
  wire act_mem_banks_bank_array_impl_data0_and_23_cse;
  wire act_mem_banks_bank_array_impl_data0_and_24_cse;
  wire act_mem_banks_bank_array_impl_data0_and_25_cse;
  wire act_mem_banks_bank_array_impl_data0_and_26_cse;
  wire act_mem_banks_bank_array_impl_data0_and_27_cse;
  wire act_mem_banks_bank_array_impl_data0_and_28_cse;
  wire act_mem_banks_bank_array_impl_data0_and_29_cse;
  wire act_mem_banks_bank_array_impl_data0_and_30_cse;
  wire act_mem_banks_bank_array_impl_data0_and_31_cse;
  wire act_mem_banks_read_read_data_and_cse;
  wire or_55_cse;
  wire or_58_cse;
  wire ActUnit_CheckStart_if_ActUnit_CheckStart_if_and_1_cse;
  wire ActUnit_RunInst_switch_lp_nor_13_cse;
  wire or_16_cse;
  wire mux_5_cse;
  wire act_port_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct_mx0;
  wire rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct_mx0;
  reg [7:0] act_config_output_counter_sva;
  reg [7:0] act_config_output_addr_base_sva;
  wire output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct_mx0;
  wire done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct_mx0;
  wire [7:0] act_mem_banks_read_for_mux_mx0w0;
  wire act_config_ActConfigRead_else_else_not_22;
  wire [7:0] act_mem_banks_read_for_mux_1_mx0w0;
  wire [7:0] act_mem_banks_read_for_mux_2_mx0w0;
  wire [7:0] act_mem_banks_read_for_mux_3_mx0w0;
  wire [7:0] act_mem_banks_read_for_mux_4_mx0w0;
  wire [7:0] act_mem_banks_read_for_mux_5_mx0w0;
  wire [7:0] act_mem_banks_read_for_mux_6_mx0w0;
  wire [7:0] act_mem_banks_read_for_mux_7_mx0w0;
  wire ActUnit_DecodeAxiRead_and_cse_1;
  wire [7:0] act_mem_banks_read_for_mux_8_mx0w0;
  wire [7:0] act_mem_banks_read_for_mux_9_mx0w0;
  reg [4:0] act_config_buffer_addr_base_sva;
  wire [7:0] act_mem_banks_read_for_mux_10_mx0w0;
  wire [7:0] act_mem_banks_read_for_mux_11_mx0w0;
  reg [7:0] act_config_num_output_sva;
  wire [7:0] act_mem_banks_read_for_mux_12_mx0w0;
  reg [5:0] act_config_num_inst_sva;
  wire [7:0] act_mem_banks_read_for_mux_13_mx0w0;
  reg [2:0] act_config_adpfloat_bias_sva;
  wire [7:0] act_mem_banks_read_for_mux_14_mx0w0;
  reg act_config_is_zero_first_sva;
  reg act_config_inst_regs_1_sva_0;
  reg act_config_inst_regs_17_sva_0;
  wire [7:0] act_mem_banks_read_for_mux_15_mx0w0;
  reg ActUnit_RunInst_switch_lp_nor_7_itm;
  reg act_config_inst_regs_16_sva_0;
  wire or_dcpl;
  wire or_dcpl_122;
  wire or_dcpl_123;
  wire or_dcpl_124;
  wire and_tmp;
  wire and_dcpl_73;
  wire while_asn_1364;
  wire while_asn_1378;
  wire [19:0] act_regs_data_0_15_sva_dfm_3;
  wire while_asn_1374;
  wire [19:0] act_regs_data_1_15_sva_dfm_3;
  wire while_asn_1370;
  wire [19:0] act_regs_data_2_15_sva_dfm_3;
  wire while_asn_1366;
  wire [19:0] act_regs_data_3_15_sva_dfm_3;
  wire [19:0] act_regs_data_0_14_sva_dfm_3;
  wire [19:0] act_regs_data_1_14_sva_dfm_3;
  wire [19:0] act_regs_data_2_14_sva_dfm_3;
  wire [19:0] act_regs_data_3_14_sva_dfm_3;
  wire [19:0] act_regs_data_0_13_sva_dfm_3;
  wire [19:0] act_regs_data_1_13_sva_dfm_3;
  wire [19:0] act_regs_data_2_13_sva_dfm_3;
  wire [19:0] act_regs_data_3_13_sva_dfm_3;
  wire [19:0] act_regs_data_0_12_sva_dfm_3;
  wire [19:0] act_regs_data_1_12_sva_dfm_3;
  wire [19:0] act_regs_data_2_12_sva_dfm_3;
  wire [19:0] act_regs_data_3_12_sva_dfm_3;
  wire [19:0] act_regs_data_0_11_sva_dfm_3;
  wire [19:0] act_regs_data_1_11_sva_dfm_3;
  wire [19:0] act_regs_data_2_11_sva_dfm_3;
  wire [19:0] act_regs_data_3_11_sva_dfm_3;
  wire [19:0] act_regs_data_0_10_sva_dfm_3;
  wire [19:0] act_regs_data_1_10_sva_dfm_3;
  wire [19:0] act_regs_data_2_10_sva_dfm_3;
  wire [19:0] act_regs_data_3_10_sva_dfm_3;
  wire [19:0] act_regs_data_0_9_sva_dfm_3;
  wire [19:0] act_regs_data_1_9_sva_dfm_3;
  wire [19:0] act_regs_data_2_9_sva_dfm_3;
  wire [19:0] act_regs_data_3_9_sva_dfm_3;
  wire [19:0] act_regs_data_0_8_sva_dfm_3;
  wire [19:0] act_regs_data_1_8_sva_dfm_3;
  wire [19:0] act_regs_data_2_8_sva_dfm_3;
  wire [19:0] act_regs_data_3_8_sva_dfm_3;
  wire [19:0] act_regs_data_0_7_sva_dfm_3;
  wire [19:0] act_regs_data_1_7_sva_dfm_3;
  wire [19:0] act_regs_data_2_7_sva_dfm_3;
  wire [19:0] act_regs_data_3_7_sva_dfm_3;
  wire [19:0] act_regs_data_0_6_sva_dfm_3;
  wire [19:0] act_regs_data_1_6_sva_dfm_3;
  wire [19:0] act_regs_data_2_6_sva_dfm_3;
  wire [19:0] act_regs_data_3_6_sva_dfm_3;
  wire [19:0] act_regs_data_0_5_sva_dfm_3;
  wire [19:0] act_regs_data_1_5_sva_dfm_3;
  wire [19:0] act_regs_data_2_5_sva_dfm_3;
  wire [19:0] act_regs_data_3_5_sva_dfm_3;
  wire [19:0] act_regs_data_0_4_sva_dfm_3;
  wire [19:0] act_regs_data_1_4_sva_dfm_3;
  wire [19:0] act_regs_data_2_4_sva_dfm_3;
  wire [19:0] act_regs_data_3_4_sva_dfm_3;
  wire [19:0] act_regs_data_0_3_sva_dfm_3;
  wire [19:0] act_regs_data_1_3_sva_dfm_3;
  wire [19:0] act_regs_data_2_3_sva_dfm_3;
  wire [19:0] act_regs_data_3_3_sva_dfm_3;
  wire [19:0] act_regs_data_0_2_sva_dfm_3;
  wire [19:0] act_regs_data_1_2_sva_dfm_3;
  wire [19:0] act_regs_data_2_2_sva_dfm_3;
  wire [19:0] act_regs_data_3_2_sva_dfm_3;
  wire [19:0] act_regs_data_0_1_sva_dfm_3;
  wire [19:0] act_regs_data_1_1_sva_dfm_3;
  wire [19:0] act_regs_data_2_1_sva_dfm_3;
  wire [19:0] act_regs_data_3_1_sva_dfm_3;
  wire [19:0] act_regs_data_0_0_sva_dfm_3;
  wire [19:0] act_regs_data_1_0_sva_dfm_3;
  wire [19:0] act_regs_data_2_0_sva_dfm_3;
  wire [19:0] act_regs_data_3_0_sva_dfm_3;
  wire act_config_output_counter_sva_mx0c1;
  wire or_887_tmp;
  reg [319:0] ActUnit_RunInst_case_8_EAdd_act_regs_data_sva;
  reg [319:0] ActUnit_RunInst_case_9_EMul_act_regs_data_sva;
  reg [319:0] ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva;
  reg [319:0] ActUnit_RunInst_case_11_Tanh_act_regs_data_sva;
  reg [319:0] ActUnit_RunInst_case_12_Relu_act_regs_data_sva;
  reg [319:0] ActUnit_RunInst_case_13_OneX_act_regs_data_sva;
  wire and_1551_tmp;
  wire nor_18_cse;
  wire nor_19_cse;
  wire nor_20_cse;
  wire nor_21_cse;
  wire or_884_itm;
  wire [127:0] out_data_out;
  wire or_tmp_756;
  reg [19:0] act_regs_data_1_15_sva;
  reg [19:0] act_regs_data_2_0_sva;
  reg [19:0] act_regs_data_1_14_sva;
  reg [19:0] act_regs_data_2_1_sva;
  reg [19:0] act_regs_data_1_13_sva;
  reg [19:0] act_regs_data_2_2_sva;
  reg [19:0] act_regs_data_1_12_sva;
  reg [19:0] act_regs_data_2_3_sva;
  reg [19:0] act_regs_data_1_11_sva;
  reg [19:0] act_regs_data_2_4_sva;
  reg [19:0] act_regs_data_1_10_sva;
  reg [19:0] act_regs_data_2_5_sva;
  reg [19:0] act_regs_data_1_9_sva;
  reg [19:0] act_regs_data_2_6_sva;
  reg [19:0] act_regs_data_1_8_sva;
  reg [19:0] act_regs_data_2_7_sva;
  reg [19:0] act_regs_data_1_7_sva;
  reg [19:0] act_regs_data_2_8_sva;
  reg [19:0] act_regs_data_1_6_sva;
  reg [19:0] act_regs_data_2_9_sva;
  reg [19:0] act_regs_data_1_5_sva;
  reg [19:0] act_regs_data_2_10_sva;
  reg [19:0] act_regs_data_1_4_sva;
  reg [19:0] act_regs_data_2_11_sva;
  reg [19:0] act_regs_data_1_3_sva;
  reg [19:0] act_regs_data_2_12_sva;
  reg [19:0] act_regs_data_1_2_sva;
  reg [19:0] act_regs_data_2_13_sva;
  reg [19:0] act_regs_data_1_1_sva;
  reg [19:0] act_regs_data_2_14_sva;
  reg [19:0] act_regs_data_1_0_sva;
  reg [19:0] act_regs_data_2_15_sva;
  reg [19:0] act_regs_data_0_15_sva;
  reg [19:0] act_regs_data_3_0_sva;
  reg [19:0] act_regs_data_0_14_sva;
  reg [19:0] act_regs_data_3_1_sva;
  reg [19:0] act_regs_data_0_13_sva;
  reg [19:0] act_regs_data_3_2_sva;
  reg [19:0] act_regs_data_0_12_sva;
  reg [19:0] act_regs_data_3_3_sva;
  reg [19:0] act_regs_data_0_11_sva;
  reg [19:0] act_regs_data_3_4_sva;
  reg [19:0] act_regs_data_0_10_sva;
  reg [19:0] act_regs_data_3_5_sva;
  reg [19:0] act_regs_data_0_9_sva;
  reg [19:0] act_regs_data_3_6_sva;
  reg [19:0] act_regs_data_0_8_sva;
  reg [19:0] act_regs_data_3_7_sva;
  reg [19:0] act_regs_data_0_7_sva;
  reg [19:0] act_regs_data_3_8_sva;
  reg [19:0] act_regs_data_0_6_sva;
  reg [19:0] act_regs_data_3_9_sva;
  reg [19:0] act_regs_data_0_5_sva;
  reg [19:0] act_regs_data_3_10_sva;
  reg [19:0] act_regs_data_0_4_sva;
  reg [19:0] act_regs_data_3_11_sva;
  reg [19:0] act_regs_data_0_3_sva;
  reg [19:0] act_regs_data_3_12_sva;
  reg [19:0] act_regs_data_0_2_sva;
  reg [19:0] act_regs_data_3_13_sva;
  reg [19:0] act_regs_data_0_1_sva;
  reg [19:0] act_regs_data_3_14_sva;
  reg [19:0] act_regs_data_0_0_sva;
  reg [19:0] act_regs_data_3_15_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva;
  reg [4:0] act_read_addrs_lpi_1_dfm_5;
  reg [7:0] act_write_data_data_0_0_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_1_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_2_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_3_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_4_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_5_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_6_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_7_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_8_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_9_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_10_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_11_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_12_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_13_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_14_lpi_1_dfm_4;
  reg [7:0] act_write_data_data_0_15_lpi_1_dfm_4;
  reg [4:0] act_write_addrs_lpi_1_dfm_5;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_0_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_1_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_2_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_3_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_4_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_5_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_6_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_7_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_8_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_9_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_10_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_11_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_12_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_13_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_14_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_15_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_16_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_17_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_18_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_19_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_20_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_21_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_22_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_23_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_24_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_25_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_26_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_27_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_28_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_29_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_30_7_0_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_127_120_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_119_112_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_111_104_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_103_96_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_95_88_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_87_80_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_79_72_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_71_64_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_63_56_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_55_48_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_47_40_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_39_32_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_31_24_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_23_16_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_15_8_sva_dfm;
  reg [7:0] act_mem_banks_bank_array_impl_data0_31_7_0_sva_dfm;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_127_120;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_119_112;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_111_104;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_103_96;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_95_88;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_87_80;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_79_72;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_71_64;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_63_56;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_55_48;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_47_40;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_39_32;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_31_24;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_23_16;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_15_8;
  reg [7:0] act_mem_banks_read_read_data_lpi_1_dfm_1_7_0;
  wire act_config_is_valid_sva_mx0c0;
  wire ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0;
  wire is_start_sva_mx0c1;
  wire [4:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_3_mx0w2;
  wire act_write_addrs_lpi_1_dfm_5_mx0c2;
  wire ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_cse_1;
  wire ActUnit_RunInst_switch_lp_nor_7_itm_mx0w0;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [19:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
  wire [4:0] while_mux_124_ssc_mx0;
  wire [4:0] act_read_addrs_lpi_1_dfm_9;
  wire [7:0] act_write_data_data_0_0_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_1_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_2_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_3_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_4_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_5_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_6_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_7_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_8_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_9_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_10_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_11_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_12_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_13_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_14_lpi_1_dfm_5_mx0;
  wire [7:0] act_write_data_data_0_15_lpi_1_dfm_5_mx0;
  wire while_asn_1290;
  wire while_asn_1292;
  wire while_asn_1294;
  wire while_asn_1296;
  wire while_asn_1298;
  wire while_asn_1300;
  wire while_asn_1302;
  wire while_asn_1304;
  wire while_asn_1306;
  wire while_asn_1308;
  wire while_asn_1310;
  wire while_asn_1312;
  wire while_asn_1314;
  wire while_asn_1316;
  wire while_asn_1318;
  wire while_asn_1320;
  wire while_asn_1322;
  wire while_asn_1324;
  wire while_asn_1326;
  wire while_asn_1328;
  wire while_asn_1330;
  wire while_asn_1332;
  wire while_asn_1334;
  wire while_asn_1336;
  wire while_asn_1338;
  wire while_asn_1340;
  wire while_asn_1342;
  wire while_asn_1344;
  wire while_asn_1346;
  wire while_asn_1348;
  wire while_asn_1350;
  wire while_asn_1352;
  wire while_asn_1354;
  wire while_asn_1356;
  wire while_asn_1358;
  wire while_asn_1360;
  wire [319:0] libraries_EAdd_0d1aed8b807329bc366abb192bb53bb66056_1;
  wire [319:0] libraries_EMul_50466378fb684d7351699b7bf1bdec8c6525_1;
  wire [319:0] libraries_Sigmoid_6ea22cc51ee279163d827d3cc5db43491cd81_1;
  wire [319:0] libraries_Tanh_0c47cc570305d1d8c1a9dd465101e61217b26_1;
  wire [319:0] libraries_Relu_29d7978308309996bcf6431af85e65007d30_1;
  wire [319:0] libraries_OneX_6a9c88d8c3af0ca712acdf3bbda5530a55e7_1;
  wire [319:0] libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1;
  reg [2:0] act_config_in_InstFetch_return_sva_4_2;
  wire mux_10_cse;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_cse;
  wire act_write_data_data_and_cse;
  wire ActUnit_PushAxiRsp_if_and_cse;
  wire ActUnit_PushAxiRsp_if_and_1_cse;
  wire mux_tmp_118;
  wire not_tmp_67;
  wire or_tmp_791;
  wire or_958_cse;
  wire or_957_cse;
  wire or_956_cse;
  wire or_955_cse;
  wire or_954_cse;
  wire or_953_cse;
  wire or_952_cse;
  wire or_951_cse;
  wire or_950_cse;
  wire or_949_cse;
  wire or_948_cse;
  wire or_947_cse;
  wire or_946_cse;
  wire or_945_cse;
  wire or_944_cse;
  wire or_943_cse;
  wire or_942_cse;
  wire or_941_cse;
  wire or_940_cse;
  wire or_939_cse;
  wire or_938_cse;
  wire or_937_cse;
  wire or_936_cse;
  wire or_935_cse;
  wire or_934_cse;
  wire or_933_cse;
  wire or_932_cse;
  wire or_931_cse;
  wire or_930_cse;
  wire or_929_cse;
  wire or_928_cse;
  wire or_925_cse;
  reg reg_act_regs_data_3_15_enexo;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo;
  reg reg_act_config_inst_counter_enexo;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_1;
  reg reg_act_regs_data_1_14_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_1;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_2;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_2;
  reg reg_act_regs_data_1_13_enexo;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_3;
  reg reg_act_regs_data_0_12_enexo;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_4;
  reg reg_act_regs_data_0_11_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_4;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_5;
  reg reg_act_regs_data_0_10_enexo;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_6;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_6;
  reg reg_act_regs_data_3_9_enexo;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_7;
  reg reg_act_regs_data_2_8_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_7;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_8;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_8;
  reg reg_act_regs_data_0_7_enexo;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_9;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_9;
  reg reg_act_regs_data_1_6_enexo;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_10;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_10;
  reg reg_act_regs_data_3_5_enexo;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_11;
  reg reg_act_regs_data_2_4_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_11;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_12;
  reg reg_act_regs_data_3_3_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_12;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_13;
  reg reg_act_regs_data_1_2_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_13;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_14;
  reg reg_act_regs_data_0_1_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_14;
  reg reg_act_config_inst_regs_19_sva_dfm_6_enexo_15;
  reg reg_act_regs_data_1_0_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_15;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_18_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_19_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_20_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_21_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_22_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_23_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_24_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_25_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_26_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_27_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_28_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_29_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_30_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_31_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_32_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_33_enex5;
  wire [19:0] nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [19:0] nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [7:0] z_out_7_0;
  wire [8:0] nl_z_out_7_0;

  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_prb;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_prb;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb;
  wire[0:0] pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb;
  wire[0:0] pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb;
  wire[0:0] nor_12_nl;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1;
  wire[0:0] act_config_InstIncr_if_act_config_InstIncr_if_and_1_nl;
  wire[0:0] ActUnit_DecodeAxi_mux_88_nl;
  wire[0:0] ActUnit_DecodeAxi_if_mux_82_nl;
  wire[0:0] ActUnit_DecodeAxiWrite_mux_36_nl;
  wire[0:0] act_config_ActConfigWrite_mux_33_nl;
  wire[7:0] mux_91_nl;
  wire[0:0] and_1557_nl;
  wire[0:0] not_235_nl;
  wire[4:0] and_1554_nl;
  wire[4:0] while_while_while_or_nl;
  wire[0:0] while_while_not_nl;
  wire[0:0] mux_19_nl;
  wire[0:0] nand_6_nl;
  wire[0:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_2_nl;
  wire[0:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_33_nl;
  wire[0:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_5_nl;
  wire[0:0] mux_158_nl;
  wire[0:0] or_960_nl;
  wire[0:0] mux_157_nl;
  wire[0:0] mux_156_nl;
  wire[0:0] mux_155_nl;
  wire[0:0] mux_154_nl;
  wire[0:0] mux_153_nl;
  wire[0:0] mux_152_nl;
  wire[0:0] mux_151_nl;
  wire[0:0] mux_150_nl;
  wire[0:0] mux_149_nl;
  wire[0:0] and_1734_nl;
  wire[0:0] and_1733_nl;
  wire[0:0] mux_148_nl;
  wire[0:0] and_1732_nl;
  wire[0:0] and_1731_nl;
  wire[0:0] mux_147_nl;
  wire[0:0] mux_146_nl;
  wire[0:0] and_1730_nl;
  wire[0:0] and_1729_nl;
  wire[0:0] mux_145_nl;
  wire[0:0] and_1728_nl;
  wire[0:0] and_1727_nl;
  wire[0:0] mux_144_nl;
  wire[0:0] mux_143_nl;
  wire[0:0] mux_142_nl;
  wire[0:0] and_1726_nl;
  wire[0:0] and_1725_nl;
  wire[0:0] mux_141_nl;
  wire[0:0] and_1724_nl;
  wire[0:0] and_1723_nl;
  wire[0:0] mux_140_nl;
  wire[0:0] mux_139_nl;
  wire[0:0] and_1722_nl;
  wire[0:0] and_1721_nl;
  wire[0:0] mux_138_nl;
  wire[0:0] and_1720_nl;
  wire[0:0] and_1719_nl;
  wire[0:0] mux_137_nl;
  wire[0:0] mux_136_nl;
  wire[0:0] mux_135_nl;
  wire[0:0] mux_134_nl;
  wire[0:0] and_1718_nl;
  wire[0:0] and_1717_nl;
  wire[0:0] mux_133_nl;
  wire[0:0] and_1716_nl;
  wire[0:0] and_1715_nl;
  wire[0:0] mux_132_nl;
  wire[0:0] mux_131_nl;
  wire[0:0] and_1714_nl;
  wire[0:0] and_1713_nl;
  wire[0:0] mux_130_nl;
  wire[0:0] and_1712_nl;
  wire[0:0] and_1711_nl;
  wire[0:0] mux_129_nl;
  wire[0:0] mux_128_nl;
  wire[0:0] mux_127_nl;
  wire[0:0] and_1710_nl;
  wire[0:0] and_1709_nl;
  wire[0:0] mux_126_nl;
  wire[0:0] and_1708_nl;
  wire[0:0] and_1707_nl;
  wire[0:0] mux_125_nl;
  wire[0:0] mux_124_nl;
  wire[0:0] and_1706_nl;
  wire[0:0] and_1705_nl;
  wire[0:0] mux_123_nl;
  wire[0:0] and_1704_nl;
  wire[0:0] and_1703_nl;
  wire[0:0] nand_nl;
  wire[0:0] while_else_1_while_else_1_nand_nl;
  wire[0:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_31_nl;
  wire[0:0] mux_4_nl;
  wire[0:0] nor_16_nl;
  wire[0:0] or_1_nl;
  wire[4:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_21_nl;
  wire[0:0] ActUnit_DecodeAxiWrite_else_not_17_nl;
  wire[1:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_1_nl;
  wire[1:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_4_nl;
  wire[1:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_7_nl;
  wire[1:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_9_nl;
  wire[1:0] act_config_ActConfigWrite_if_mux_3_nl;
  wire[1:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_11_nl;
  wire[1:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_13_nl;
  wire[1:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_15_nl;
  wire[1:0] act_config_ActConfigWrite_if_mux_5_nl;
  wire[1:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_17_nl;
  wire[1:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_19_nl;
  wire[1:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_21_nl;
  wire[1:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_23_nl;
  wire[1:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_25_nl;
  wire[1:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_27_nl;
  wire[1:0] nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_29_nl;
  wire[0:0] ActUnit_DecodeAxi_mux_89_nl;
  wire[0:0] ActUnit_DecodeAxi_if_mux_83_nl;
  wire[0:0] ActUnit_DecodeAxiWrite_mux_37_nl;
  wire[0:0] act_config_ActConfigWrite_mux_34_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_22_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_23_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_24_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_25_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_26_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_27_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_28_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_29_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_30_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_31_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_32_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_33_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_34_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_35_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_36_nl;
  wire[7:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_37_nl;
  wire[4:0] ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_and_1_nl;
  wire[0:0] mux_nl;
  wire[0:0] nor_14_nl;
  wire[0:0] mux_15_nl;
  wire[0:0] or_64_nl;
  wire[0:0] mux_121_nl;
  wire[0:0] mux_120_nl;
  wire[0:0] mux_119_nl;
  wire[0:0] mux_118_nl;
  wire[0:0] mux_117_nl;
  wire[0:0] mux_116_nl;
  wire[0:0] mux_115_nl;
  wire[0:0] mux_114_nl;
  wire[0:0] mux_113_nl;
  wire[0:0] mux_112_nl;
  wire[0:0] mux_111_nl;
  wire[0:0] mux_110_nl;
  wire[0:0] mux_109_nl;
  wire[0:0] mux_108_nl;
  wire[0:0] mux_107_nl;
  wire[0:0] mux_106_nl;
  wire[0:0] mux_105_nl;
  wire[0:0] mux_104_nl;
  wire[0:0] mux_103_nl;
  wire[0:0] mux_102_nl;
  wire[0:0] mux_101_nl;
  wire[0:0] mux_100_nl;
  wire[0:0] mux_99_nl;
  wire[0:0] mux_98_nl;
  wire[0:0] mux_97_nl;
  wire[0:0] mux_96_nl;
  wire[0:0] mux_95_nl;
  wire[0:0] mux_94_nl;
  wire[0:0] mux_93_nl;
  wire[0:0] mux_92_nl;
  wire[2:0] operator_8_false_operator_8_false_and_1_nl;
  wire[0:0] operator_8_false_nor_1_nl;
  wire[4:0] operator_8_false_operator_8_false_mux_2_nl;
  wire[4:0] operator_8_false_operator_8_false_mux_3_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [319:0] nl_EAdd_rg_in_1_data;
  assign nl_EAdd_rg_in_1_data = {nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1};
  wire [319:0] nl_EAdd_rg_in_2_data;
  assign nl_EAdd_rg_in_2_data = {nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm};
  wire [319:0] nl_EMul_rg_in_1_data;
  assign nl_EMul_rg_in_1_data = {nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      , nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1};
  wire [319:0] nl_EMul_rg_in_2_data;
  assign nl_EMul_rg_in_2_data = {nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm};
  wire [319:0] nl_Sigmoid_rg_in_data;
  assign nl_Sigmoid_rg_in_data = {nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm};
  wire [319:0] nl_Tanh_rg_in_data;
  assign nl_Tanh_rg_in_data = {nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm};
  wire [319:0] nl_Relu_rg_in_data;
  assign nl_Relu_rg_in_data = {nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm};
  wire [319:0] nl_OneX_rg_in_data;
  assign nl_OneX_rg_in_data = {nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm};
  wire[7:0] act_mem_banks_read_for_mux_22_nl;
  wire[7:0] act_mem_banks_read_for_mux_28_nl;
  wire[7:0] act_mem_banks_read_for_mux_31_nl;
  wire[7:0] act_mem_banks_read_for_mux_37_nl;
  wire[7:0] act_mem_banks_read_for_mux_40_nl;
  wire[7:0] act_mem_banks_read_for_mux_46_nl;
  wire[7:0] act_mem_banks_read_for_mux_49_nl;
  wire[7:0] act_mem_banks_read_for_mux_55_nl;
  wire[7:0] act_mem_banks_read_for_mux_58_nl;
  wire[7:0] act_mem_banks_read_for_mux_64_nl;
  wire[7:0] act_mem_banks_read_for_mux_67_nl;
  wire[7:0] act_mem_banks_read_for_mux_61_nl;
  wire[7:0] act_mem_banks_read_for_mux_52_nl;
  wire[7:0] act_mem_banks_read_for_mux_43_nl;
  wire[7:0] act_mem_banks_read_for_mux_34_nl;
  wire[7:0] act_mem_banks_read_for_mux_25_nl;
  wire [127:0] nl_Adpfloat2Fixed_1_rg_in_data;
  assign act_mem_banks_read_for_mux_22_nl = MUX_v_8_2_2(act_mem_banks_read_read_data_lpi_1_dfm_1_127_120,
      act_mem_banks_read_for_mux_mx0w0, ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_1_tmp);
  assign act_mem_banks_read_for_mux_28_nl = MUX_v_8_2_2(act_mem_banks_read_read_data_lpi_1_dfm_1_119_112,
      act_mem_banks_read_for_mux_1_mx0w0, ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_1_tmp);
  assign act_mem_banks_read_for_mux_31_nl = MUX_v_8_2_2(act_mem_banks_read_read_data_lpi_1_dfm_1_111_104,
      act_mem_banks_read_for_mux_2_mx0w0, ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_1_tmp);
  assign act_mem_banks_read_for_mux_37_nl = MUX_v_8_2_2(act_mem_banks_read_read_data_lpi_1_dfm_1_103_96,
      act_mem_banks_read_for_mux_3_mx0w0, ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_1_tmp);
  assign act_mem_banks_read_for_mux_40_nl = MUX_v_8_2_2(act_mem_banks_read_read_data_lpi_1_dfm_1_95_88,
      act_mem_banks_read_for_mux_4_mx0w0, ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_1_tmp);
  assign act_mem_banks_read_for_mux_46_nl = MUX_v_8_2_2(act_mem_banks_read_read_data_lpi_1_dfm_1_87_80,
      act_mem_banks_read_for_mux_5_mx0w0, ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_1_tmp);
  assign act_mem_banks_read_for_mux_49_nl = MUX_v_8_2_2(act_mem_banks_read_read_data_lpi_1_dfm_1_79_72,
      act_mem_banks_read_for_mux_6_mx0w0, ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_1_tmp);
  assign act_mem_banks_read_for_mux_55_nl = MUX_v_8_2_2(act_mem_banks_read_read_data_lpi_1_dfm_1_71_64,
      act_mem_banks_read_for_mux_7_mx0w0, ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_1_tmp);
  assign act_mem_banks_read_for_mux_58_nl = MUX_v_8_2_2(act_mem_banks_read_read_data_lpi_1_dfm_1_63_56,
      act_mem_banks_read_for_mux_8_mx0w0, ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_1_tmp);
  assign act_mem_banks_read_for_mux_64_nl = MUX_v_8_2_2(act_mem_banks_read_read_data_lpi_1_dfm_1_55_48,
      act_mem_banks_read_for_mux_9_mx0w0, ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_1_tmp);
  assign act_mem_banks_read_for_mux_67_nl = MUX_v_8_2_2(act_mem_banks_read_read_data_lpi_1_dfm_1_47_40,
      act_mem_banks_read_for_mux_10_mx0w0, ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_1_tmp);
  assign act_mem_banks_read_for_mux_61_nl = MUX_v_8_2_2(act_mem_banks_read_read_data_lpi_1_dfm_1_39_32,
      act_mem_banks_read_for_mux_11_mx0w0, ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_1_tmp);
  assign act_mem_banks_read_for_mux_52_nl = MUX_v_8_2_2(act_mem_banks_read_read_data_lpi_1_dfm_1_31_24,
      act_mem_banks_read_for_mux_12_mx0w0, ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_1_tmp);
  assign act_mem_banks_read_for_mux_43_nl = MUX_v_8_2_2(act_mem_banks_read_read_data_lpi_1_dfm_1_23_16,
      act_mem_banks_read_for_mux_13_mx0w0, ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_1_tmp);
  assign act_mem_banks_read_for_mux_34_nl = MUX_v_8_2_2(act_mem_banks_read_read_data_lpi_1_dfm_1_15_8,
      act_mem_banks_read_for_mux_14_mx0w0, ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_1_tmp);
  assign act_mem_banks_read_for_mux_25_nl = MUX_v_8_2_2(act_mem_banks_read_read_data_lpi_1_dfm_1_7_0,
      act_mem_banks_read_for_mux_15_mx0w0, ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_1_tmp);
  assign nl_Adpfloat2Fixed_1_rg_in_data = {act_mem_banks_read_for_mux_22_nl , act_mem_banks_read_for_mux_28_nl
      , act_mem_banks_read_for_mux_31_nl , act_mem_banks_read_for_mux_37_nl , act_mem_banks_read_for_mux_40_nl
      , act_mem_banks_read_for_mux_46_nl , act_mem_banks_read_for_mux_49_nl , act_mem_banks_read_for_mux_55_nl
      , act_mem_banks_read_for_mux_58_nl , act_mem_banks_read_for_mux_64_nl , act_mem_banks_read_for_mux_67_nl
      , act_mem_banks_read_for_mux_61_nl , act_mem_banks_read_for_mux_52_nl , act_mem_banks_read_for_mux_43_nl
      , act_mem_banks_read_for_mux_34_nl , act_mem_banks_read_for_mux_25_nl};
  wire[19:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_nl;
  wire[0:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_nl;
  wire[0:0] ActUnit_PushOutput_if_and_1_nl;
  wire[0:0] ActUnit_PushOutput_if_and_2_nl;
  wire[0:0] ActUnit_PushOutput_if_and_3_nl;
  wire[19:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_1_nl;
  wire[0:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_16_nl;
  wire[0:0] ActUnit_PushOutput_if_and_5_nl;
  wire[0:0] ActUnit_PushOutput_if_and_6_nl;
  wire[0:0] ActUnit_PushOutput_if_and_7_nl;
  wire[19:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_2_nl;
  wire[0:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_17_nl;
  wire[0:0] ActUnit_PushOutput_if_and_9_nl;
  wire[0:0] ActUnit_PushOutput_if_and_10_nl;
  wire[0:0] ActUnit_PushOutput_if_and_11_nl;
  wire[19:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_3_nl;
  wire[0:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_18_nl;
  wire[0:0] ActUnit_PushOutput_if_and_13_nl;
  wire[0:0] ActUnit_PushOutput_if_and_14_nl;
  wire[0:0] ActUnit_PushOutput_if_and_15_nl;
  wire[19:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_4_nl;
  wire[0:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_19_nl;
  wire[0:0] ActUnit_PushOutput_if_and_17_nl;
  wire[0:0] ActUnit_PushOutput_if_and_18_nl;
  wire[0:0] ActUnit_PushOutput_if_and_19_nl;
  wire[19:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_5_nl;
  wire[0:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_20_nl;
  wire[0:0] ActUnit_PushOutput_if_and_21_nl;
  wire[0:0] ActUnit_PushOutput_if_and_22_nl;
  wire[0:0] ActUnit_PushOutput_if_and_23_nl;
  wire[19:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_6_nl;
  wire[0:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_21_nl;
  wire[0:0] ActUnit_PushOutput_if_and_25_nl;
  wire[0:0] ActUnit_PushOutput_if_and_26_nl;
  wire[0:0] ActUnit_PushOutput_if_and_27_nl;
  wire[19:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_7_nl;
  wire[0:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_22_nl;
  wire[0:0] ActUnit_PushOutput_if_and_29_nl;
  wire[0:0] ActUnit_PushOutput_if_and_30_nl;
  wire[0:0] ActUnit_PushOutput_if_and_31_nl;
  wire[19:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_8_nl;
  wire[0:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_23_nl;
  wire[0:0] ActUnit_PushOutput_if_and_33_nl;
  wire[0:0] ActUnit_PushOutput_if_and_34_nl;
  wire[0:0] ActUnit_PushOutput_if_and_35_nl;
  wire[19:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_9_nl;
  wire[0:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_24_nl;
  wire[0:0] ActUnit_PushOutput_if_and_37_nl;
  wire[0:0] ActUnit_PushOutput_if_and_38_nl;
  wire[0:0] ActUnit_PushOutput_if_and_39_nl;
  wire[19:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_10_nl;
  wire[0:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_25_nl;
  wire[0:0] ActUnit_PushOutput_if_and_41_nl;
  wire[0:0] ActUnit_PushOutput_if_and_42_nl;
  wire[0:0] ActUnit_PushOutput_if_and_43_nl;
  wire[19:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_11_nl;
  wire[0:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_26_nl;
  wire[0:0] ActUnit_PushOutput_if_and_45_nl;
  wire[0:0] ActUnit_PushOutput_if_and_46_nl;
  wire[0:0] ActUnit_PushOutput_if_and_47_nl;
  wire[19:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_12_nl;
  wire[0:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_27_nl;
  wire[0:0] ActUnit_PushOutput_if_and_49_nl;
  wire[0:0] ActUnit_PushOutput_if_and_50_nl;
  wire[0:0] ActUnit_PushOutput_if_and_51_nl;
  wire[19:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_13_nl;
  wire[0:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_28_nl;
  wire[0:0] ActUnit_PushOutput_if_and_53_nl;
  wire[0:0] ActUnit_PushOutput_if_and_54_nl;
  wire[0:0] ActUnit_PushOutput_if_and_55_nl;
  wire[19:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_14_nl;
  wire[0:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_29_nl;
  wire[0:0] ActUnit_PushOutput_if_and_57_nl;
  wire[0:0] ActUnit_PushOutput_if_and_58_nl;
  wire[0:0] ActUnit_PushOutput_if_and_59_nl;
  wire[19:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_15_nl;
  wire[0:0] ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_30_nl;
  wire[0:0] ActUnit_PushOutput_if_and_61_nl;
  wire[0:0] ActUnit_PushOutput_if_and_62_nl;
  wire[0:0] ActUnit_PushOutput_if_and_63_nl;
  wire [319:0] nl_Fixed2Adpfloat_rg_in_data;
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_nl = ~((nvhls_get_slc_2U_NVUINT8_return_3_sva_1!=2'b00)
      | (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_1_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b01)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_2_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b10)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_3_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b11)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_nl = MUX1HOT_v_20_5_2(act_regs_data_0_15_sva_dfm_3,
      act_regs_data_1_15_sva_dfm_3, act_regs_data_2_15_sva_dfm_3, act_regs_data_3_15_sva_dfm_3,
      nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm,
      {ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_nl , ActUnit_PushOutput_if_and_1_nl
      , ActUnit_PushOutput_if_and_2_nl , ActUnit_PushOutput_if_and_3_nl , (fsm_output[1])});
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_16_nl = ~((nvhls_get_slc_2U_NVUINT8_return_3_sva_1!=2'b00)
      | (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_5_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b01)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_6_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b10)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_7_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b11)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_1_nl = MUX1HOT_v_20_5_2(act_regs_data_0_14_sva_dfm_3,
      act_regs_data_1_14_sva_dfm_3, act_regs_data_2_14_sva_dfm_3, act_regs_data_3_14_sva_dfm_3,
      nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm,
      {ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_16_nl , ActUnit_PushOutput_if_and_5_nl
      , ActUnit_PushOutput_if_and_6_nl , ActUnit_PushOutput_if_and_7_nl , (fsm_output[1])});
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_17_nl = ~((nvhls_get_slc_2U_NVUINT8_return_3_sva_1!=2'b00)
      | (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_9_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b01)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_10_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b10)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_11_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b11)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_2_nl = MUX1HOT_v_20_5_2(act_regs_data_0_13_sva_dfm_3,
      act_regs_data_1_13_sva_dfm_3, act_regs_data_2_13_sva_dfm_3, act_regs_data_3_13_sva_dfm_3,
      nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm,
      {ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_17_nl , ActUnit_PushOutput_if_and_9_nl
      , ActUnit_PushOutput_if_and_10_nl , ActUnit_PushOutput_if_and_11_nl , (fsm_output[1])});
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_18_nl = ~((nvhls_get_slc_2U_NVUINT8_return_3_sva_1!=2'b00)
      | (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_13_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b01)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_14_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b10)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_15_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b11)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_3_nl = MUX1HOT_v_20_5_2(act_regs_data_0_12_sva_dfm_3,
      act_regs_data_1_12_sva_dfm_3, act_regs_data_2_12_sva_dfm_3, act_regs_data_3_12_sva_dfm_3,
      nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm,
      {ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_18_nl , ActUnit_PushOutput_if_and_13_nl
      , ActUnit_PushOutput_if_and_14_nl , ActUnit_PushOutput_if_and_15_nl , (fsm_output[1])});
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_19_nl = ~((nvhls_get_slc_2U_NVUINT8_return_3_sva_1!=2'b00)
      | (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_17_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b01)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_18_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b10)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_19_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b11)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_4_nl = MUX1HOT_v_20_5_2(act_regs_data_0_11_sva_dfm_3,
      act_regs_data_1_11_sva_dfm_3, act_regs_data_2_11_sva_dfm_3, act_regs_data_3_11_sva_dfm_3,
      nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm,
      {ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_19_nl , ActUnit_PushOutput_if_and_17_nl
      , ActUnit_PushOutput_if_and_18_nl , ActUnit_PushOutput_if_and_19_nl , (fsm_output[1])});
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_20_nl = ~((nvhls_get_slc_2U_NVUINT8_return_3_sva_1!=2'b00)
      | (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_21_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b01)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_22_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b10)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_23_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b11)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_5_nl = MUX1HOT_v_20_5_2(act_regs_data_0_10_sva_dfm_3,
      act_regs_data_1_10_sva_dfm_3, act_regs_data_2_10_sva_dfm_3, act_regs_data_3_10_sva_dfm_3,
      nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm,
      {ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_20_nl , ActUnit_PushOutput_if_and_21_nl
      , ActUnit_PushOutput_if_and_22_nl , ActUnit_PushOutput_if_and_23_nl , (fsm_output[1])});
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_21_nl = ~((nvhls_get_slc_2U_NVUINT8_return_3_sva_1!=2'b00)
      | (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_25_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b01)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_26_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b10)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_27_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b11)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_6_nl = MUX1HOT_v_20_5_2(act_regs_data_0_9_sva_dfm_3,
      act_regs_data_1_9_sva_dfm_3, act_regs_data_2_9_sva_dfm_3, act_regs_data_3_9_sva_dfm_3,
      nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm,
      {ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_21_nl , ActUnit_PushOutput_if_and_25_nl
      , ActUnit_PushOutput_if_and_26_nl , ActUnit_PushOutput_if_and_27_nl , (fsm_output[1])});
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_22_nl = ~((nvhls_get_slc_2U_NVUINT8_return_3_sva_1!=2'b00)
      | (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_29_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b01)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_30_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b10)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_31_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b11)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_7_nl = MUX1HOT_v_20_5_2(act_regs_data_0_8_sva_dfm_3,
      act_regs_data_1_8_sva_dfm_3, act_regs_data_2_8_sva_dfm_3, act_regs_data_3_8_sva_dfm_3,
      nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm,
      {ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_22_nl , ActUnit_PushOutput_if_and_29_nl
      , ActUnit_PushOutput_if_and_30_nl , ActUnit_PushOutput_if_and_31_nl , (fsm_output[1])});
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_23_nl = ~((nvhls_get_slc_2U_NVUINT8_return_3_sva_1!=2'b00)
      | (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_33_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b01)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_34_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b10)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_35_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b11)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_8_nl = MUX1HOT_v_20_5_2(act_regs_data_0_7_sva_dfm_3,
      act_regs_data_1_7_sva_dfm_3, act_regs_data_2_7_sva_dfm_3, act_regs_data_3_7_sva_dfm_3,
      nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm,
      {ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_23_nl , ActUnit_PushOutput_if_and_33_nl
      , ActUnit_PushOutput_if_and_34_nl , ActUnit_PushOutput_if_and_35_nl , (fsm_output[1])});
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_24_nl = ~((nvhls_get_slc_2U_NVUINT8_return_3_sva_1!=2'b00)
      | (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_37_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b01)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_38_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b10)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_39_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b11)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_9_nl = MUX1HOT_v_20_5_2(act_regs_data_0_6_sva_dfm_3,
      act_regs_data_1_6_sva_dfm_3, act_regs_data_2_6_sva_dfm_3, act_regs_data_3_6_sva_dfm_3,
      nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm,
      {ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_24_nl , ActUnit_PushOutput_if_and_37_nl
      , ActUnit_PushOutput_if_and_38_nl , ActUnit_PushOutput_if_and_39_nl , (fsm_output[1])});
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_25_nl = ~((nvhls_get_slc_2U_NVUINT8_return_3_sva_1!=2'b00)
      | (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_41_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b01)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_42_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b10)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_43_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b11)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_10_nl = MUX1HOT_v_20_5_2(act_regs_data_0_5_sva_dfm_3,
      act_regs_data_1_5_sva_dfm_3, act_regs_data_2_5_sva_dfm_3, act_regs_data_3_5_sva_dfm_3,
      nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm,
      {ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_25_nl , ActUnit_PushOutput_if_and_41_nl
      , ActUnit_PushOutput_if_and_42_nl , ActUnit_PushOutput_if_and_43_nl , (fsm_output[1])});
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_26_nl = ~((nvhls_get_slc_2U_NVUINT8_return_3_sva_1!=2'b00)
      | (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_45_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b01)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_46_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b10)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_47_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b11)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_11_nl = MUX1HOT_v_20_5_2(act_regs_data_0_4_sva_dfm_3,
      act_regs_data_1_4_sva_dfm_3, act_regs_data_2_4_sva_dfm_3, act_regs_data_3_4_sva_dfm_3,
      nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm,
      {ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_26_nl , ActUnit_PushOutput_if_and_45_nl
      , ActUnit_PushOutput_if_and_46_nl , ActUnit_PushOutput_if_and_47_nl , (fsm_output[1])});
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_27_nl = ~((nvhls_get_slc_2U_NVUINT8_return_3_sva_1!=2'b00)
      | (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_49_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b01)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_50_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b10)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_51_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b11)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_12_nl = MUX1HOT_v_20_5_2(act_regs_data_0_3_sva_dfm_3,
      act_regs_data_1_3_sva_dfm_3, act_regs_data_2_3_sva_dfm_3, act_regs_data_3_3_sva_dfm_3,
      nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm,
      {ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_27_nl , ActUnit_PushOutput_if_and_49_nl
      , ActUnit_PushOutput_if_and_50_nl , ActUnit_PushOutput_if_and_51_nl , (fsm_output[1])});
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_28_nl = ~((nvhls_get_slc_2U_NVUINT8_return_3_sva_1!=2'b00)
      | (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_53_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b01)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_54_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b10)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_55_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b11)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_13_nl = MUX1HOT_v_20_5_2(act_regs_data_0_2_sva_dfm_3,
      act_regs_data_1_2_sva_dfm_3, act_regs_data_2_2_sva_dfm_3, act_regs_data_3_2_sva_dfm_3,
      nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm,
      {ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_28_nl , ActUnit_PushOutput_if_and_53_nl
      , ActUnit_PushOutput_if_and_54_nl , ActUnit_PushOutput_if_and_55_nl , (fsm_output[1])});
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_29_nl = ~((nvhls_get_slc_2U_NVUINT8_return_3_sva_1!=2'b00)
      | (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_57_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b01)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_58_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b10)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_59_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b11)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_14_nl = MUX1HOT_v_20_5_2(act_regs_data_0_1_sva_dfm_3,
      act_regs_data_1_1_sva_dfm_3, act_regs_data_2_1_sva_dfm_3, act_regs_data_3_1_sva_dfm_3,
      nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm,
      {ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_29_nl , ActUnit_PushOutput_if_and_57_nl
      , ActUnit_PushOutput_if_and_58_nl , ActUnit_PushOutput_if_and_59_nl , (fsm_output[1])});
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_30_nl = ~((nvhls_get_slc_2U_NVUINT8_return_3_sva_1!=2'b00)
      | (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_61_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b01)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_62_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b10)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_and_63_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b11)
      & (~ (fsm_output[1]));
  assign ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_15_nl = MUX1HOT_v_20_5_2(act_regs_data_0_0_sva_dfm_3,
      act_regs_data_1_0_sva_dfm_3, act_regs_data_2_0_sva_dfm_3, act_regs_data_3_0_sva_dfm_3,
      nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm,
      {ActUnit_PushOutput_if_ActUnit_PushOutput_if_nor_30_nl , ActUnit_PushOutput_if_and_61_nl
      , ActUnit_PushOutput_if_and_62_nl , ActUnit_PushOutput_if_and_63_nl , (fsm_output[1])});
  assign nl_Fixed2Adpfloat_rg_in_data = {ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_nl
      , ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_1_nl , ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_2_nl
      , ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_3_nl , ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_4_nl
      , ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_5_nl , ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_6_nl
      , ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_7_nl , ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_8_nl
      , ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_9_nl , ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_10_nl
      , ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_11_nl , ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_12_nl
      , ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_13_nl , ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_14_nl
      , ActUnit_PushOutput_if_ActUnit_PushOutput_if_mux1h_15_nl};
  wire[7:0] ActUnit_PushAxiRsp_if_mux_10_nl;
  wire[7:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_47_nl;
  wire[7:0] act_config_ActConfigRead_else_else_mux_18_nl;
  wire[7:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_40_nl;
  wire[7:0] ActUnit_PushAxiRsp_if_mux_9_nl;
  wire[7:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_45_nl;
  wire[7:0] act_config_ActConfigRead_else_else_mux_17_nl;
  wire[7:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_39_nl;
  wire[7:0] ActUnit_PushAxiRsp_if_mux_8_nl;
  wire[7:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_43_nl;
  wire[7:0] act_config_ActConfigRead_else_else_mux_16_nl;
  wire[7:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_38_nl;
  wire[7:0] ActUnit_PushAxiRsp_if_mux_7_nl;
  wire[7:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_41_nl;
  wire[7:0] act_config_ActConfigRead_else_else_mux_15_nl;
  wire[7:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_37_nl;
  wire[7:0] ActUnit_PushAxiRsp_if_mux_6_nl;
  wire[7:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_39_nl;
  wire[7:0] act_config_ActConfigRead_else_else_mux_14_nl;
  wire[7:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_36_nl;
  wire[7:0] ActUnit_PushAxiRsp_if_mux_5_nl;
  wire[7:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_37_nl;
  wire[7:0] act_config_ActConfigRead_else_else_mux_13_nl;
  wire[7:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_35_nl;
  wire[7:0] ActUnit_PushAxiRsp_if_mux_4_nl;
  wire[7:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_35_nl;
  wire[7:0] act_config_ActConfigRead_else_else_mux_12_nl;
  wire[7:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_34_nl;
  wire[7:0] and_1686_nl;
  wire[7:0] mux1h_65_nl;
  wire[0:0] not_366_nl;
  wire[7:0] ActUnit_PushAxiRsp_if_mux_2_nl;
  wire[7:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_33_nl;
  wire[7:0] act_config_ActConfigRead_else_else_mux_11_nl;
  wire[7:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_33_nl;
  wire[2:0] act_mem_banks_read_read_data_mux_9_nl;
  wire[2:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_31_nl;
  wire[2:0] act_config_ActConfigRead_else_else_mux_10_nl;
  wire[2:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_32_nl;
  wire[4:0] and_1687_nl;
  wire[4:0] mux1h_66_nl;
  wire[0:0] not_370_nl;
  wire[7:0] ActUnit_PushAxiRsp_if_mux_1_nl;
  wire[7:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_29_nl;
  wire[7:0] act_config_ActConfigRead_else_else_mux_9_nl;
  wire[7:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_31_nl;
  wire[7:0] and_1688_nl;
  wire[7:0] mux1h_67_nl;
  wire[0:0] not_374_nl;
  wire[1:0] act_mem_banks_read_read_data_mux_7_nl;
  wire[1:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_27_nl;
  wire[1:0] act_config_ActConfigRead_else_else_mux_8_nl;
  wire[1:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_30_nl;
  wire[5:0] and_1689_nl;
  wire[5:0] mux1h_68_nl;
  wire[0:0] act_mem_banks_read_read_data_and_19_nl;
  wire[0:0] act_mem_banks_read_read_data_and_20_nl;
  wire[0:0] act_mem_banks_read_read_data_and_21_nl;
  wire[0:0] not_378_nl;
  wire[4:0] act_mem_banks_read_read_data_mux_5_nl;
  wire[4:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_25_nl;
  wire[4:0] act_config_ActConfigRead_else_else_mux_7_nl;
  wire[4:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_29_nl;
  wire[2:0] and_1690_nl;
  wire[2:0] mux1h_69_nl;
  wire[0:0] not_382_nl;
  wire[6:0] act_mem_banks_read_read_data_mux_3_nl;
  wire[6:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_23_nl;
  wire[6:0] act_config_ActConfigRead_else_else_mux_6_nl;
  wire[6:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_28_nl;
  wire[0:0] act_mem_banks_read_read_data_mux_2_nl;
  wire[0:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_50_nl;
  wire[0:0] ActUnit_DecodeAxiRead_mux_27_nl;
  wire[0:0] act_config_ActConfigRead_else_mux_18_nl;
  wire[0:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_19_nl;
  wire[6:0] act_mem_banks_read_read_data_mux_1_nl;
  wire[6:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_21_nl;
  wire[6:0] act_config_ActConfigRead_else_else_mux_5_nl;
  wire[6:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_27_nl;
  wire[0:0] act_mem_banks_read_read_data_mux_nl;
  wire[0:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_49_nl;
  wire[0:0] ActUnit_DecodeAxiRead_mux_28_nl;
  wire[0:0] act_config_ActConfigRead_else_mux_20_nl;
  wire[0:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_21_nl;
  wire [127:0] nl_ActUnit_ActUnitRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_ActUnitRun;
  assign act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_40_nl
      = MUX_v_8_2_2(8'b00000000, act_config_inst_regs_31_sva_dfm_6, act_config_ActConfigRead_else_else_not_22);
  assign act_config_ActConfigRead_else_else_mux_18_nl = MUX_v_8_2_2(act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_40_nl,
      act_config_inst_regs_15_sva_dfm_5, and_dcpl_65);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_47_nl = act_config_ActConfigRead_else_else_mux_18_nl
      & ({{7{act_config_ActConfigRead_unequal_tmp_1}}, act_config_ActConfigRead_unequal_tmp_1})
      & (signext_8_1(~ ActUnit_DecodeAxiRead_unequal_tmp_1));
  assign ActUnit_PushAxiRsp_if_mux_10_nl = MUX_v_8_2_2(act_mem_banks_read_for_mux_mx0w0,
      ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_47_nl, or_dcpl_9);
  assign act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_39_nl
      = MUX_v_8_2_2(8'b00000000, act_config_inst_regs_30_sva_dfm_6, act_config_ActConfigRead_else_else_not_22);
  assign act_config_ActConfigRead_else_else_mux_17_nl = MUX_v_8_2_2(act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_39_nl,
      act_config_inst_regs_14_sva_dfm_5, and_dcpl_65);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_45_nl = act_config_ActConfigRead_else_else_mux_17_nl
      & ({{7{act_config_ActConfigRead_unequal_tmp_1}}, act_config_ActConfigRead_unequal_tmp_1})
      & (signext_8_1(~ ActUnit_DecodeAxiRead_unequal_tmp_1));
  assign ActUnit_PushAxiRsp_if_mux_9_nl = MUX_v_8_2_2(act_mem_banks_read_for_mux_1_mx0w0,
      ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_45_nl, or_dcpl_9);
  assign act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_38_nl
      = MUX_v_8_2_2(8'b00000000, act_config_inst_regs_29_sva_dfm_6, act_config_ActConfigRead_else_else_not_22);
  assign act_config_ActConfigRead_else_else_mux_16_nl = MUX_v_8_2_2(act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_38_nl,
      act_config_inst_regs_13_sva_dfm_5, and_dcpl_65);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_43_nl = act_config_ActConfigRead_else_else_mux_16_nl
      & ({{7{act_config_ActConfigRead_unequal_tmp_1}}, act_config_ActConfigRead_unequal_tmp_1})
      & (signext_8_1(~ ActUnit_DecodeAxiRead_unequal_tmp_1));
  assign ActUnit_PushAxiRsp_if_mux_8_nl = MUX_v_8_2_2(act_mem_banks_read_for_mux_2_mx0w0,
      ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_43_nl, or_dcpl_9);
  assign act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_37_nl
      = MUX_v_8_2_2(8'b00000000, act_config_inst_regs_28_sva_dfm_6, act_config_ActConfigRead_else_else_not_22);
  assign act_config_ActConfigRead_else_else_mux_15_nl = MUX_v_8_2_2(act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_37_nl,
      act_config_inst_regs_12_sva_dfm_5, and_dcpl_65);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_41_nl = act_config_ActConfigRead_else_else_mux_15_nl
      & ({{7{act_config_ActConfigRead_unequal_tmp_1}}, act_config_ActConfigRead_unequal_tmp_1})
      & (signext_8_1(~ ActUnit_DecodeAxiRead_unequal_tmp_1));
  assign ActUnit_PushAxiRsp_if_mux_7_nl = MUX_v_8_2_2(act_mem_banks_read_for_mux_3_mx0w0,
      ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_41_nl, or_dcpl_9);
  assign act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_36_nl
      = MUX_v_8_2_2(8'b00000000, act_config_inst_regs_27_sva_dfm_6, act_config_ActConfigRead_else_else_not_22);
  assign act_config_ActConfigRead_else_else_mux_14_nl = MUX_v_8_2_2(act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_36_nl,
      act_config_inst_regs_11_sva_dfm_5, and_dcpl_65);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_39_nl = act_config_ActConfigRead_else_else_mux_14_nl
      & ({{7{act_config_ActConfigRead_unequal_tmp_1}}, act_config_ActConfigRead_unequal_tmp_1})
      & (signext_8_1(~ ActUnit_DecodeAxiRead_unequal_tmp_1));
  assign ActUnit_PushAxiRsp_if_mux_6_nl = MUX_v_8_2_2(act_mem_banks_read_for_mux_4_mx0w0,
      ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_39_nl, or_dcpl_9);
  assign act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_35_nl
      = MUX_v_8_2_2(8'b00000000, act_config_inst_regs_26_sva_dfm_6, act_config_ActConfigRead_else_else_not_22);
  assign act_config_ActConfigRead_else_else_mux_13_nl = MUX_v_8_2_2(act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_35_nl,
      act_config_inst_regs_10_sva_dfm_5, and_dcpl_65);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_37_nl = act_config_ActConfigRead_else_else_mux_13_nl
      & ({{7{act_config_ActConfigRead_unequal_tmp_1}}, act_config_ActConfigRead_unequal_tmp_1})
      & (signext_8_1(~ ActUnit_DecodeAxiRead_unequal_tmp_1));
  assign ActUnit_PushAxiRsp_if_mux_5_nl = MUX_v_8_2_2(act_mem_banks_read_for_mux_5_mx0w0,
      ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_37_nl, or_dcpl_9);
  assign act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_34_nl
      = MUX_v_8_2_2(8'b00000000, act_config_inst_regs_25_sva_dfm_6, act_config_ActConfigRead_else_else_not_22);
  assign act_config_ActConfigRead_else_else_mux_12_nl = MUX_v_8_2_2(act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_34_nl,
      act_config_inst_regs_9_sva_dfm_5, and_dcpl_65);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_35_nl = act_config_ActConfigRead_else_else_mux_12_nl
      & ({{7{act_config_ActConfigRead_unequal_tmp_1}}, act_config_ActConfigRead_unequal_tmp_1})
      & (signext_8_1(~ ActUnit_DecodeAxiRead_unequal_tmp_1));
  assign ActUnit_PushAxiRsp_if_mux_4_nl = MUX_v_8_2_2(act_mem_banks_read_for_mux_6_mx0w0,
      ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_35_nl, or_dcpl_9);
  assign mux1h_65_nl = MUX1HOT_v_8_4_2(act_mem_banks_read_for_mux_7_mx0w0, act_config_output_addr_base_sva,
      act_config_inst_regs_24_sva_dfm_6, act_config_inst_regs_8_sva_dfm_5, {(~ or_dcpl_9)
      , ActUnit_PushAxiRsp_if_and_cse , ActUnit_PushAxiRsp_if_and_1_cse , ActUnit_DecodeAxiRead_and_10_cse});
  assign not_366_nl = ~ and_dcpl_73;
  assign and_1686_nl = MUX_v_8_2_2(8'b00000000, mux1h_65_nl, not_366_nl);
  assign act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_33_nl
      = MUX_v_8_2_2(8'b00000000, act_config_inst_regs_23_sva_dfm_6, act_config_ActConfigRead_else_else_not_22);
  assign act_config_ActConfigRead_else_else_mux_11_nl = MUX_v_8_2_2(act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_33_nl,
      act_config_inst_regs_7_sva_dfm_5, and_dcpl_65);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_33_nl = act_config_ActConfigRead_else_else_mux_11_nl
      & ({{7{act_config_ActConfigRead_unequal_tmp_1}}, act_config_ActConfigRead_unequal_tmp_1})
      & (signext_8_1(~ ActUnit_DecodeAxiRead_unequal_tmp_1));
  assign ActUnit_PushAxiRsp_if_mux_2_nl = MUX_v_8_2_2(act_mem_banks_read_for_mux_8_mx0w0,
      ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_33_nl, or_dcpl_9);
  assign act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_32_nl
      = MUX_v_3_2_2(3'b000, (act_config_inst_regs_22_sva_dfm_6[7:5]), act_config_ActConfigRead_else_else_not_22);
  assign act_config_ActConfigRead_else_else_mux_10_nl = MUX_v_3_2_2(act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_32_nl,
      (act_config_inst_regs_6_sva_dfm_5[7:5]), and_dcpl_65);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_31_nl = act_config_ActConfigRead_else_else_mux_10_nl
      & ({{2{act_config_ActConfigRead_unequal_tmp_1}}, act_config_ActConfigRead_unequal_tmp_1})
      & (signext_3_1(~ ActUnit_DecodeAxiRead_unequal_tmp_1));
  assign act_mem_banks_read_read_data_mux_9_nl = MUX_v_3_2_2((act_mem_banks_read_for_mux_9_mx0w0[7:5]),
      ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_31_nl, or_dcpl_9);
  assign mux1h_66_nl = MUX1HOT_v_5_4_2((act_mem_banks_read_for_mux_9_mx0w0[4:0]),
      act_config_buffer_addr_base_sva, (act_config_inst_regs_22_sva_dfm_6[4:0]),
      (act_config_inst_regs_6_sva_dfm_5[4:0]), {(~ or_dcpl_9) , ActUnit_PushAxiRsp_if_and_cse
      , ActUnit_PushAxiRsp_if_and_1_cse , ActUnit_DecodeAxiRead_and_10_cse});
  assign not_370_nl = ~ and_dcpl_73;
  assign and_1687_nl = MUX_v_5_2_2(5'b00000, mux1h_66_nl, not_370_nl);
  assign act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_31_nl
      = MUX_v_8_2_2(8'b00000000, act_config_inst_regs_21_sva_dfm_6, act_config_ActConfigRead_else_else_not_22);
  assign act_config_ActConfigRead_else_else_mux_9_nl = MUX_v_8_2_2(act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_31_nl,
      act_config_inst_regs_5_sva_dfm_5, and_dcpl_65);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_29_nl = act_config_ActConfigRead_else_else_mux_9_nl
      & ({{7{act_config_ActConfigRead_unequal_tmp_1}}, act_config_ActConfigRead_unequal_tmp_1})
      & (signext_8_1(~ ActUnit_DecodeAxiRead_unequal_tmp_1));
  assign ActUnit_PushAxiRsp_if_mux_1_nl = MUX_v_8_2_2(act_mem_banks_read_for_mux_10_mx0w0,
      ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_29_nl, or_dcpl_9);
  assign mux1h_67_nl = MUX1HOT_v_8_4_2(act_mem_banks_read_for_mux_11_mx0w0, act_config_num_output_sva,
      act_config_inst_regs_20_sva_dfm_6, act_config_inst_regs_4_sva_dfm_5, {(~ or_dcpl_9)
      , ActUnit_PushAxiRsp_if_and_cse , ActUnit_PushAxiRsp_if_and_1_cse , ActUnit_DecodeAxiRead_and_10_cse});
  assign not_374_nl = ~ and_dcpl_73;
  assign and_1688_nl = MUX_v_8_2_2(8'b00000000, mux1h_67_nl, not_374_nl);
  assign act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_30_nl
      = MUX_v_2_2_2(2'b00, (act_config_inst_regs_19_sva_dfm_6[7:6]), act_config_ActConfigRead_else_else_not_22);
  assign act_config_ActConfigRead_else_else_mux_8_nl = MUX_v_2_2_2(act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_30_nl,
      (act_config_inst_regs_3_sva_dfm_5[7:6]), and_dcpl_65);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_27_nl = act_config_ActConfigRead_else_else_mux_8_nl
      & ({{1{act_config_ActConfigRead_unequal_tmp_1}}, act_config_ActConfigRead_unequal_tmp_1})
      & (signext_2_1(~ ActUnit_DecodeAxiRead_unequal_tmp_1));
  assign act_mem_banks_read_read_data_mux_7_nl = MUX_v_2_2_2((act_mem_banks_read_for_mux_12_mx0w0[7:6]),
      ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_27_nl, or_dcpl_9);
  assign act_mem_banks_read_read_data_and_19_nl = (~ ActUnit_DecodeAxiRead_and_cse_1)
      & or_dcpl_9 & (~ and_1551_tmp);
  assign act_mem_banks_read_read_data_and_20_nl = ActUnit_DecodeAxiRead_and_9_cse
      & or_dcpl_9 & (~ and_1551_tmp);
  assign act_mem_banks_read_read_data_and_21_nl = ActUnit_DecodeAxiRead_and_10_cse
      & or_dcpl_9 & (~ and_1551_tmp);
  assign mux1h_68_nl = MUX1HOT_v_6_4_2((act_mem_banks_read_for_mux_12_mx0w0[5:0]),
      act_config_num_inst_sva, (act_config_inst_regs_19_sva_dfm_6[5:0]), (act_config_inst_regs_3_sva_dfm_5[5:0]),
      {(~ or_dcpl_9) , act_mem_banks_read_read_data_and_19_nl , act_mem_banks_read_read_data_and_20_nl
      , act_mem_banks_read_read_data_and_21_nl});
  assign not_378_nl = ~ and_1551_tmp;
  assign and_1689_nl = MUX_v_6_2_2(6'b000000, mux1h_68_nl, not_378_nl);
  assign act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_29_nl
      = MUX_v_5_2_2(5'b00000, (act_config_inst_regs_18_sva_dfm_6[7:3]), act_config_ActConfigRead_else_else_not_22);
  assign act_config_ActConfigRead_else_else_mux_7_nl = MUX_v_5_2_2(act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_29_nl,
      (act_config_inst_regs_2_sva_dfm_5[7:3]), and_dcpl_65);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_25_nl = act_config_ActConfigRead_else_else_mux_7_nl
      & ({{4{act_config_ActConfigRead_unequal_tmp_1}}, act_config_ActConfigRead_unequal_tmp_1})
      & (signext_5_1(~ ActUnit_DecodeAxiRead_unequal_tmp_1));
  assign act_mem_banks_read_read_data_mux_5_nl = MUX_v_5_2_2((act_mem_banks_read_for_mux_13_mx0w0[7:3]),
      ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_25_nl, or_dcpl_9);
  assign mux1h_69_nl = MUX1HOT_v_3_4_2((act_mem_banks_read_for_mux_13_mx0w0[2:0]),
      act_config_adpfloat_bias_sva, (act_config_inst_regs_18_sva_dfm_6[2:0]), (act_config_inst_regs_2_sva_dfm_5[2:0]),
      {(~ or_dcpl_9) , ActUnit_PushAxiRsp_if_and_cse , ActUnit_PushAxiRsp_if_and_1_cse
      , ActUnit_DecodeAxiRead_and_10_cse});
  assign not_382_nl = ~ and_dcpl_73;
  assign and_1690_nl = MUX_v_3_2_2(3'b000, mux1h_69_nl, not_382_nl);
  assign act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_28_nl
      = MUX_v_7_2_2(7'b0000000, (act_config_inst_regs_17_sva_dfm_6[7:1]), act_config_ActConfigRead_else_else_not_22);
  assign act_config_ActConfigRead_else_else_mux_6_nl = MUX_v_7_2_2(act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_28_nl,
      (act_config_inst_regs_1_sva_dfm_5[7:1]), and_dcpl_65);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_23_nl = act_config_ActConfigRead_else_else_mux_6_nl
      & ({{6{act_config_ActConfigRead_unequal_tmp_1}}, act_config_ActConfigRead_unequal_tmp_1})
      & (signext_7_1(~ ActUnit_DecodeAxiRead_unequal_tmp_1));
  assign act_mem_banks_read_read_data_mux_3_nl = MUX_v_7_2_2((act_mem_banks_read_for_mux_14_mx0w0[7:1]),
      ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_23_nl, or_dcpl_9);
  assign act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_19_nl
      = act_config_inst_regs_17_sva_0 & act_config_ActConfigRead_else_else_not_22;
  assign act_config_ActConfigRead_else_mux_18_nl = MUX_s_1_2_2(act_config_inst_regs_1_sva_0,
      act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_19_nl,
      act_config_ActConfigRead_else_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_mux_27_nl = MUX_s_1_2_2(act_config_is_zero_first_sva,
      act_config_ActConfigRead_else_mux_18_nl, act_config_ActConfigRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_50_nl = ActUnit_DecodeAxiRead_mux_27_nl
      & (~ ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign act_mem_banks_read_read_data_mux_2_nl = MUX_s_1_2_2((act_mem_banks_read_for_mux_14_mx0w0[0]),
      ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_50_nl, or_dcpl_9);
  assign act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_27_nl
      = MUX_v_7_2_2(7'b0000000, (act_config_inst_regs_16_sva_dfm_6[7:1]), act_config_ActConfigRead_else_else_not_22);
  assign act_config_ActConfigRead_else_else_mux_5_nl = MUX_v_7_2_2(act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_27_nl,
      (act_config_inst_regs_0_sva_dfm_5[7:1]), and_dcpl_65);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_21_nl = act_config_ActConfigRead_else_else_mux_5_nl
      & ({{6{act_config_ActConfigRead_unequal_tmp_1}}, act_config_ActConfigRead_unequal_tmp_1})
      & (signext_7_1(~ ActUnit_DecodeAxiRead_unequal_tmp_1));
  assign act_mem_banks_read_read_data_mux_1_nl = MUX_v_7_2_2((act_mem_banks_read_for_mux_15_mx0w0[7:1]),
      ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_21_nl, or_dcpl_9);
  assign act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_21_nl
      = act_config_inst_regs_16_sva_0 & act_config_ActConfigRead_else_else_not_22;
  assign act_config_ActConfigRead_else_mux_20_nl = MUX_s_1_2_2(ActUnit_RunInst_switch_lp_nor_7_itm,
      act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_21_nl,
      act_config_ActConfigRead_else_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_mux_28_nl = MUX_s_1_2_2(act_config_is_valid_sva, act_config_ActConfigRead_else_mux_20_nl,
      act_config_ActConfigRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_49_nl = ActUnit_DecodeAxiRead_mux_28_nl
      & (~ ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign act_mem_banks_read_read_data_mux_nl = MUX_s_1_2_2((act_mem_banks_read_for_mux_15_mx0w0[0]),
      ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_49_nl, or_dcpl_9);
  assign nl_ActUnit_ActUnitRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_ActUnitRun
      = {ActUnit_PushAxiRsp_if_mux_10_nl , ActUnit_PushAxiRsp_if_mux_9_nl , ActUnit_PushAxiRsp_if_mux_8_nl
      , ActUnit_PushAxiRsp_if_mux_7_nl , ActUnit_PushAxiRsp_if_mux_6_nl , ActUnit_PushAxiRsp_if_mux_5_nl
      , ActUnit_PushAxiRsp_if_mux_4_nl , and_1686_nl , ActUnit_PushAxiRsp_if_mux_2_nl
      , act_mem_banks_read_read_data_mux_9_nl , and_1687_nl , ActUnit_PushAxiRsp_if_mux_1_nl
      , and_1688_nl , act_mem_banks_read_read_data_mux_7_nl , and_1689_nl , act_mem_banks_read_read_data_mux_5_nl
      , and_1690_nl , act_mem_banks_read_read_data_mux_3_nl , act_mem_banks_read_read_data_mux_2_nl
      , act_mem_banks_read_read_data_mux_1_nl , act_mem_banks_read_read_data_mux_nl};
  wire [127:0] nl_ActUnit_ActUnitRun_output_port_Push_mioi_inst_output_port_Push_mioi_m_data_data_rsc_dat_ActUnitRun;
  assign nl_ActUnit_ActUnitRun_output_port_Push_mioi_inst_output_port_Push_mioi_m_data_data_rsc_dat_ActUnitRun
      = out_data_out;
  wire [7:0] nl_ActUnit_ActUnitRun_output_port_Push_mioi_inst_output_port_Push_mioi_m_logical_addr_rsc_dat_ActUnitRun;
  assign nl_ActUnit_ActUnitRun_output_port_Push_mioi_inst_output_port_Push_mioi_m_logical_addr_rsc_dat_ActUnitRun
      = act_config_output_counter_sva + act_config_output_addr_base_sva;
  ActUnit_EAdd  EAdd_rg (
      .in_1_data(nl_EAdd_rg_in_1_data[319:0]),
      .in_2_data(nl_EAdd_rg_in_2_data[319:0]),
      .out_data(libraries_EAdd_0d1aed8b807329bc366abb192bb53bb66056_1)
    );
  ActUnit_EMul  EMul_rg (
      .in_1_data(nl_EMul_rg_in_1_data[319:0]),
      .in_2_data(nl_EMul_rg_in_2_data[319:0]),
      .out_data(libraries_EMul_50466378fb684d7351699b7bf1bdec8c6525_1)
    );
  ActUnit_Sigmoid  Sigmoid_rg (
      .in_data(nl_Sigmoid_rg_in_data[319:0]),
      .out_data(libraries_Sigmoid_6ea22cc51ee279163d827d3cc5db43491cd81_1)
    );
  ActUnit_Tanh  Tanh_rg (
      .in_data(nl_Tanh_rg_in_data[319:0]),
      .out_data(libraries_Tanh_0c47cc570305d1d8c1a9dd465101e61217b26_1)
    );
  ActUnit_Relu  Relu_rg (
      .in_data(nl_Relu_rg_in_data[319:0]),
      .out_data(libraries_Relu_29d7978308309996bcf6431af85e65007d30_1)
    );
  ActUnit_OneX  OneX_rg (
      .in_data(nl_OneX_rg_in_data[319:0]),
      .out_data(libraries_OneX_6a9c88d8c3af0ca712acdf3bbda5530a55e7_1)
    );
  ActUnit_Adpfloat2Fixed  Adpfloat2Fixed_1_rg (
      .in_data(nl_Adpfloat2Fixed_1_rg_in_data[127:0]),
      .out_data(libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1),
      .adpfloat_bias(act_config_adpfloat_bias_sva)
    );
  ActUnit_Fixed2Adpfloat  Fixed2Adpfloat_rg (
      .in_data(nl_Fixed2Adpfloat_rg_in_data[319:0]),
      .out_data(out_data_out),
      .adpfloat_bias(act_config_adpfloat_bias_sva)
    );
  ActUnit_ActUnit_ActUnitRun_rva_in_PopNB_mioi ActUnit_ActUnitRun_rva_in_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_in_val(rva_in_val),
      .rva_in_rdy(rva_in_rdy),
      .rva_in_msg(rva_in_msg),
      .ActUnitRun_wen(ActUnitRun_wen),
      .rva_in_PopNB_mioi_oswt(reg_rva_in_PopNB_mioi_iswt0_cse),
      .ActUnitRun_wten(ActUnitRun_wten),
      .rva_in_PopNB_mioi_data_data_rsc_z_mxwt(rva_in_PopNB_mioi_data_data_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_addr_rsc_z_mxwt(rva_in_PopNB_mioi_data_addr_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_rw_rsc_z_mxwt(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt),
      .rva_in_PopNB_mioi_return_rsc_z_mxwt(rva_in_PopNB_mioi_return_rsc_z_mxwt),
      .rva_in_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct(and_158_cse)
    );
  ActUnit_ActUnit_ActUnitRun_act_port_PopNB_mioi ActUnit_ActUnitRun_act_port_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .act_port_val(act_port_val),
      .act_port_rdy(act_port_rdy),
      .act_port_msg(act_port_msg),
      .ActUnitRun_wen(ActUnitRun_wen),
      .ActUnitRun_wten(ActUnitRun_wten),
      .act_port_PopNB_mioi_oswt(reg_act_port_PopNB_mioi_iswt0_cse),
      .act_port_PopNB_mioi_data_data_rsc_z_mxwt(act_port_PopNB_mioi_data_data_rsc_z_mxwt),
      .act_port_PopNB_mioi_return_rsc_z_mxwt(act_port_PopNB_mioi_return_rsc_z_mxwt),
      .act_port_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct(act_port_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct_mx0)
    );
  ActUnit_ActUnit_ActUnitRun_rva_out_Push_mioi ActUnit_ActUnitRun_rva_out_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_out_val(rva_out_val),
      .rva_out_rdy(rva_out_rdy),
      .rva_out_msg(rva_out_msg),
      .ActUnitRun_wen(ActUnitRun_wen),
      .rva_out_Push_mioi_oswt(reg_rva_out_Push_mioi_iswt0_cse),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp),
      .rva_out_Push_mioi_m_data_rsc_dat_ActUnitRun(nl_ActUnit_ActUnitRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_ActUnitRun[127:0]),
      .rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct(rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct_mx0)
    );
  ActUnit_ActUnit_ActUnitRun_start_PopNB_mioi ActUnit_ActUnitRun_start_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .start_val(start_val),
      .start_rdy(start_rdy),
      .start_msg(start_msg),
      .ActUnitRun_wen(ActUnitRun_wen),
      .ActUnitRun_wten(ActUnitRun_wten),
      .start_PopNB_mioi_oswt(reg_start_PopNB_mioi_iswt0_cse),
      .start_PopNB_mioi_data_rsc_z_mxwt(start_PopNB_mioi_data_rsc_z_mxwt),
      .start_PopNB_mioi_return_rsc_z_mxwt(start_PopNB_mioi_return_rsc_z_mxwt),
      .start_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct(or_tmp_61)
    );
  ActUnit_ActUnit_ActUnitRun_output_port_Push_mioi ActUnit_ActUnitRun_output_port_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .output_port_val(output_port_val),
      .output_port_rdy(output_port_rdy),
      .output_port_msg(output_port_msg),
      .ActUnitRun_wen(ActUnitRun_wen),
      .output_port_Push_mioi_oswt(reg_output_port_Push_mioi_iswt0_cse),
      .output_port_Push_mioi_wen_comp(output_port_Push_mioi_wen_comp),
      .output_port_Push_mioi_m_data_data_rsc_dat_ActUnitRun(nl_ActUnit_ActUnitRun_output_port_Push_mioi_inst_output_port_Push_mioi_m_data_data_rsc_dat_ActUnitRun[127:0]),
      .output_port_Push_mioi_m_logical_addr_rsc_dat_ActUnitRun(nl_ActUnit_ActUnitRun_output_port_Push_mioi_inst_output_port_Push_mioi_m_logical_addr_rsc_dat_ActUnitRun[7:0]),
      .output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct(output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct_mx0)
    );
  ActUnit_ActUnit_ActUnitRun_done_Push_mioi ActUnit_ActUnitRun_done_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .done_val(done_val),
      .done_rdy(done_rdy),
      .done_msg(done_msg),
      .ActUnitRun_wen(ActUnitRun_wen),
      .done_Push_mioi_oswt(reg_done_Push_mioi_iswt0_cse),
      .done_Push_mioi_wen_comp(done_Push_mioi_wen_comp),
      .done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct(done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct_mx0)
    );
  ActUnit_ActUnit_ActUnitRun_staller ActUnit_ActUnitRun_staller_inst (
      .clk(clk),
      .rst(rst),
      .ActUnitRun_wen(ActUnitRun_wen),
      .ActUnitRun_wten(ActUnitRun_wten),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp),
      .output_port_Push_mioi_wen_comp(output_port_Push_mioi_wen_comp),
      .done_Push_mioi_wen_comp(done_Push_mioi_wen_comp)
    );
  ActUnit_ActUnit_ActUnitRun_ActUnitRun_fsm ActUnit_ActUnitRun_ActUnitRun_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .ActUnitRun_wen(ActUnitRun_wen),
      .fsm_output(fsm_output)
    );
  assign or_55_cse = mux_5_cse & (fsm_output[2]);
  assign act_mem_banks_write_if_for_if_mux_cse = MUX1HOT_s_1_1_2(1'b1, or_55_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb = act_mem_banks_write_if_for_if_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /u/huaixil/workspace/FlexASR/hls/ActUnit/../..//matchlib/cmod/include/mem_array.h: line 146
  // psl default clock = (posedge clk);
  // psl ActUnit_ActUnitRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb );
  assign act_mem_banks_write_if_for_if_mux_1_cse = MUX1HOT_s_1_1_2(ActUnitRun_wen,
      or_55_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb = act_mem_banks_write_if_for_if_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb = act_mem_banks_write_if_for_if_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /u/huaixil/workspace/FlexASR/hls/ActUnit/../..//matchlib/cmod/include/mem_array.h: line 147
  // psl ActUnit_ActUnitRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb = act_mem_banks_write_if_for_if_mux_1_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb
      = act_mem_banks_write_if_for_if_mux_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /u/huaixil/workspace/FlexASR/hls/ActUnit/../..//matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl ActUnit_ActUnitRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb
      = act_mem_banks_write_if_for_if_mux_1_cse;
  assign nor_12_nl = ~((~ rva_in_PopNB_mioi_return_rsc_z_mxwt) | rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:8]!=4'b1001));
  assign mux_10_cse = MUX_s_1_2_2(nor_12_nl, ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_1_tmp,
      is_start_sva);
  assign or_58_cse = mux_10_cse & (fsm_output[2]);
  assign act_mem_banks_read_for_mux_16_cse = MUX1HOT_s_1_1_2(1'b1, or_58_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1 = act_mem_banks_read_for_mux_16_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /u/huaixil/workspace/FlexASR/hls/ActUnit/../..//matchlib/cmod/include/mem_array.h: line 126
  // psl ActUnit_ActUnitRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1 );
  assign act_mem_banks_read_for_mux_17_cse = MUX1HOT_s_1_1_2(ActUnitRun_wen, or_58_cse);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1 = act_mem_banks_read_for_mux_17_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1 = act_mem_banks_read_for_mux_16_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /u/huaixil/workspace/FlexASR/hls/ActUnit/../..//matchlib/cmod/include/mem_array.h: line 127
  // psl ActUnit_ActUnitRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1 = act_mem_banks_read_for_mux_17_cse;
  assign ActUnit_DecodeAxiRead_and_9_cse = (~ and_dcpl_65) & ActUnit_DecodeAxiRead_and_cse_1;
  assign ActUnit_DecodeAxiRead_and_10_cse = and_dcpl_65 & ActUnit_DecodeAxiRead_and_cse_1;
  assign act_regs_data_and_cse = ActUnitRun_wen & (fsm_output[2]);
  assign nor_18_cse = ~(while_asn_1378 | or_dcpl);
  assign nor_19_cse = ~(while_asn_1374 | or_dcpl_122);
  assign nor_20_cse = ~(while_asn_1370 | or_dcpl_123);
  assign nor_21_cse = ~(while_asn_1366 | or_dcpl_124);
  assign act_config_adpfloat_bias_and_cse = ActUnitRun_wen & (~((~ (fsm_output[2]))
      | or_dcpl_22 | or_dcpl_15 | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]) | is_start_sva
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]))));
  assign act_config_inst_regs_and_cse = ActUnitRun_wen & (~((~ (fsm_output[2])) |
      not_tmp_34));
  assign act_config_inst_regs_and_16_cse = ActUnitRun_wen & (~((~ (fsm_output[2]))
      | or_dcpl_27));
  assign or_887_tmp = (act_config_output_counter_sva_mx0c1 & act_config_InstIncr_if_act_config_InstIncr_if_if_act_config_InstIncr_if_if_nor_mdf_sva_1)
      | ((~((~((~ is_start_sva) | (operator_6_false_acc_tmp[5]) | (~ act_config_InstIncr_if_equal_1_tmp)
      | (operator_6_false_acc_tmp[6]) | and_dcpl_45)) | ActUnit_DecodeAxiRead_unequal_tmp_1))
      & (fsm_output[2]));
  assign or_884_itm = or_dcpl_116 | ActUnit_DecodeAxiRead_unequal_tmp_1;
  assign act_mem_banks_bank_array_impl_data0_and_cse = ActUnitRun_wen & (~((~ (fsm_output[2]))
      | (~ mux_5_cse) | or_dcpl_35 | or_dcpl_33));
  assign act_mem_banks_bank_array_impl_data0_and_1_cse = ActUnitRun_wen & (~((~ (fsm_output[2]))
      | (~ mux_5_cse) | or_dcpl_35 | or_dcpl_38));
  assign act_mem_banks_bank_array_impl_data0_and_2_cse = ActUnitRun_wen & (~((~ (fsm_output[2]))
      | (~ mux_5_cse) | or_dcpl_35 | or_dcpl_41));
  assign act_mem_banks_bank_array_impl_data0_and_3_cse = ActUnitRun_wen & (~((~ (fsm_output[2]))
      | (~ mux_5_cse) | or_dcpl_35 | or_dcpl_44));
  assign act_mem_banks_bank_array_impl_data0_and_4_cse = ActUnitRun_wen & (~((~ (fsm_output[2]))
      | (~ mux_5_cse) | or_dcpl_47 | or_dcpl_33));
  assign act_mem_banks_bank_array_impl_data0_and_5_cse = ActUnitRun_wen & (~((~ (fsm_output[2]))
      | (~ mux_5_cse) | or_dcpl_47 | or_dcpl_38));
  assign act_mem_banks_bank_array_impl_data0_and_6_cse = ActUnitRun_wen & (~((~ (fsm_output[2]))
      | (~ mux_5_cse) | or_dcpl_47 | or_dcpl_41));
  assign act_mem_banks_bank_array_impl_data0_and_7_cse = ActUnitRun_wen & (~((~ (fsm_output[2]))
      | (~ mux_5_cse) | or_dcpl_47 | or_dcpl_44));
  assign act_mem_banks_bank_array_impl_data0_and_8_cse = ActUnitRun_wen & (~((~ (fsm_output[2]))
      | (~ mux_5_cse) | or_dcpl_57 | or_dcpl_33));
  assign act_mem_banks_bank_array_impl_data0_and_9_cse = ActUnitRun_wen & (~((~ (fsm_output[2]))
      | (~ mux_5_cse) | or_dcpl_57 | or_dcpl_38));
  assign act_mem_banks_bank_array_impl_data0_and_10_cse = ActUnitRun_wen & (~((~
      (fsm_output[2])) | (~ mux_5_cse) | or_dcpl_57 | or_dcpl_41));
  assign act_mem_banks_bank_array_impl_data0_and_11_cse = ActUnitRun_wen & (~((~
      (fsm_output[2])) | (~ mux_5_cse) | or_dcpl_57 | or_dcpl_44));
  assign act_mem_banks_bank_array_impl_data0_and_12_cse = ActUnitRun_wen & (~((~
      (fsm_output[2])) | (~ mux_5_cse) | or_dcpl_66 | or_dcpl_33));
  assign act_mem_banks_bank_array_impl_data0_and_13_cse = ActUnitRun_wen & (~((~
      (fsm_output[2])) | (~ mux_5_cse) | or_dcpl_66 | or_dcpl_38));
  assign act_mem_banks_bank_array_impl_data0_and_14_cse = ActUnitRun_wen & (~((~
      (fsm_output[2])) | (~ mux_5_cse) | or_dcpl_66 | or_dcpl_41));
  assign act_mem_banks_bank_array_impl_data0_and_15_cse = ActUnitRun_wen & (~((~
      (fsm_output[2])) | (~ mux_5_cse) | or_dcpl_66 | or_dcpl_44));
  assign act_mem_banks_bank_array_impl_data0_and_16_cse = ActUnitRun_wen & (~((~
      (fsm_output[2])) | (~ mux_5_cse) | or_dcpl_76 | or_dcpl_33));
  assign act_mem_banks_bank_array_impl_data0_and_17_cse = ActUnitRun_wen & (~((~
      (fsm_output[2])) | (~ mux_5_cse) | or_dcpl_76 | or_dcpl_38));
  assign act_mem_banks_bank_array_impl_data0_and_18_cse = ActUnitRun_wen & (~((~
      (fsm_output[2])) | (~ mux_5_cse) | or_dcpl_76 | or_dcpl_41));
  assign act_mem_banks_bank_array_impl_data0_and_19_cse = ActUnitRun_wen & (~((~
      (fsm_output[2])) | (~ mux_5_cse) | or_dcpl_76 | or_dcpl_44));
  assign act_mem_banks_bank_array_impl_data0_and_20_cse = ActUnitRun_wen & (~((~
      (fsm_output[2])) | (~ mux_5_cse) | or_dcpl_85 | or_dcpl_33));
  assign act_mem_banks_bank_array_impl_data0_and_21_cse = ActUnitRun_wen & (~((~
      (fsm_output[2])) | (~ mux_5_cse) | or_dcpl_85 | or_dcpl_38));
  assign act_mem_banks_bank_array_impl_data0_and_22_cse = ActUnitRun_wen & (~((~
      (fsm_output[2])) | (~ mux_5_cse) | or_dcpl_85 | or_dcpl_41));
  assign act_mem_banks_bank_array_impl_data0_and_23_cse = ActUnitRun_wen & (~((~
      (fsm_output[2])) | (~ mux_5_cse) | or_dcpl_85 | or_dcpl_44));
  assign act_mem_banks_bank_array_impl_data0_and_24_cse = ActUnitRun_wen & (~((~
      (fsm_output[2])) | (~ mux_5_cse) | or_dcpl_95 | or_dcpl_33));
  assign act_mem_banks_bank_array_impl_data0_and_25_cse = ActUnitRun_wen & (~((~
      (fsm_output[2])) | (~ mux_5_cse) | or_dcpl_95 | or_dcpl_38));
  assign act_mem_banks_bank_array_impl_data0_and_26_cse = ActUnitRun_wen & (~((~
      (fsm_output[2])) | (~ mux_5_cse) | or_dcpl_95 | or_dcpl_41));
  assign act_mem_banks_bank_array_impl_data0_and_27_cse = ActUnitRun_wen & (~((~
      (fsm_output[2])) | (~ mux_5_cse) | or_dcpl_95 | or_dcpl_44));
  assign act_mem_banks_bank_array_impl_data0_and_28_cse = ActUnitRun_wen & (~((~
      (fsm_output[2])) | (~ mux_5_cse) | or_dcpl_104 | or_dcpl_33));
  assign act_mem_banks_bank_array_impl_data0_and_29_cse = ActUnitRun_wen & (~((~
      (fsm_output[2])) | (~ mux_5_cse) | or_dcpl_104 | or_dcpl_38));
  assign act_mem_banks_bank_array_impl_data0_and_30_cse = ActUnitRun_wen & (~((~
      (fsm_output[2])) | (~ mux_5_cse) | or_dcpl_104 | or_dcpl_41));
  assign act_mem_banks_bank_array_impl_data0_and_31_cse = ActUnitRun_wen & (~((~
      (fsm_output[2])) | (~ mux_5_cse) | or_dcpl_104 | or_dcpl_44));
  assign ActUnit_CheckStart_if_ActUnit_CheckStart_if_and_1_cse = start_PopNB_mioi_data_rsc_z_mxwt
      & act_config_is_valid_sva & start_PopNB_mioi_return_rsc_z_mxwt;
  assign act_mem_banks_read_read_data_and_cse = ActUnitRun_wen & (fsm_output[2])
      & mux_10_cse;
  assign or_958_cse = (act_config_inst_regs_0_sva_dfm_5[7:4]!=4'b0010);
  assign or_957_cse = (act_config_inst_regs_1_sva_dfm_5[7:4]!=4'b0010);
  assign or_956_cse = (act_config_inst_regs_2_sva_dfm_5[7:4]!=4'b0010);
  assign or_955_cse = (act_config_inst_regs_3_sva_dfm_5[7:4]!=4'b0010);
  assign or_954_cse = (act_config_inst_regs_4_sva_dfm_5[7:4]!=4'b0010);
  assign or_953_cse = (act_config_inst_regs_5_sva_dfm_5[7:4]!=4'b0010);
  assign or_952_cse = (act_config_inst_regs_6_sva_dfm_5[7:4]!=4'b0010);
  assign or_951_cse = (act_config_inst_regs_7_sva_dfm_5[7:4]!=4'b0010);
  assign or_950_cse = (act_config_inst_regs_8_sva_dfm_5[7:4]!=4'b0010);
  assign or_949_cse = (act_config_inst_regs_9_sva_dfm_5[7:4]!=4'b0010);
  assign or_948_cse = (act_config_inst_regs_10_sva_dfm_5[7:4]!=4'b0010);
  assign or_947_cse = (act_config_inst_regs_11_sva_dfm_5[7:4]!=4'b0010);
  assign or_946_cse = (act_config_inst_regs_12_sva_dfm_5[7:4]!=4'b0010);
  assign or_945_cse = (act_config_inst_regs_13_sva_dfm_5[7:4]!=4'b0010);
  assign or_944_cse = (act_config_inst_regs_14_sva_dfm_5[7:4]!=4'b0010);
  assign or_943_cse = (act_config_inst_regs_15_sva_dfm_5[7:4]!=4'b0010);
  assign or_942_cse = (act_config_inst_regs_16_sva_dfm_6[7:4]!=4'b0010);
  assign or_941_cse = (act_config_inst_regs_17_sva_dfm_6[7:4]!=4'b0010);
  assign or_940_cse = (act_config_inst_regs_18_sva_dfm_6[7:4]!=4'b0010);
  assign or_939_cse = (act_config_inst_regs_19_sva_dfm_6[7:4]!=4'b0010);
  assign or_938_cse = (act_config_inst_regs_20_sva_dfm_6[7:4]!=4'b0010);
  assign or_937_cse = (act_config_inst_regs_21_sva_dfm_6[7:4]!=4'b0010);
  assign or_936_cse = (act_config_inst_regs_22_sva_dfm_6[7:4]!=4'b0010);
  assign or_935_cse = (act_config_inst_regs_23_sva_dfm_6[7:4]!=4'b0010);
  assign or_934_cse = (act_config_inst_regs_24_sva_dfm_6[7:4]!=4'b0010);
  assign or_933_cse = (act_config_inst_regs_25_sva_dfm_6[7:4]!=4'b0010);
  assign or_932_cse = (act_config_inst_regs_26_sva_dfm_6[7:4]!=4'b0010);
  assign or_931_cse = (act_config_inst_regs_27_sva_dfm_6[7:4]!=4'b0010);
  assign or_930_cse = (act_config_inst_regs_28_sva_dfm_6[7:4]!=4'b0010);
  assign or_929_cse = (act_config_inst_regs_29_sva_dfm_6[7:4]!=4'b0010);
  assign or_928_cse = (act_config_inst_regs_30_sva_dfm_6[7:4]!=4'b0010);
  assign or_925_cse = (act_config_inst_regs_31_sva_dfm_6[7:4]!=4'b0010);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_cse = ActUnitRun_wen
      & mux_tmp_1 & and_dcpl_1 & and_dcpl;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_18_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_cse
      & (reg_act_config_inst_regs_19_sva_dfm_6_enexo | reg_act_regs_data_3_15_enexo
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo | reg_act_config_inst_counter_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_19_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_cse
      & (reg_act_config_inst_regs_19_sva_dfm_6_enexo_1 | reg_act_regs_data_1_14_enexo
      | reg_act_config_inst_counter_enexo | reg_act_config_inst_regs_4_sva_dfm_5_enexo_1);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_20_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_2 | reg_act_config_inst_regs_19_sva_dfm_6_enexo_2
      | reg_act_regs_data_1_13_enexo | reg_act_config_inst_counter_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_21_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_cse
      & (reg_act_config_inst_regs_19_sva_dfm_6_enexo_3 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_3
      | reg_act_config_inst_counter_enexo | reg_act_regs_data_0_12_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_22_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_cse
      & (reg_act_config_inst_regs_19_sva_dfm_6_enexo_4 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_4
      | reg_act_regs_data_0_11_enexo | reg_act_config_inst_counter_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_23_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_5 | reg_act_config_inst_regs_19_sva_dfm_6_enexo_5
      | reg_act_regs_data_0_10_enexo | reg_act_config_inst_counter_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_24_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_6 | reg_act_regs_data_3_9_enexo
      | reg_act_config_inst_regs_19_sva_dfm_6_enexo_6 | reg_act_config_inst_counter_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_25_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_cse
      & (reg_act_config_inst_regs_19_sva_dfm_6_enexo_7 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_7
      | reg_act_regs_data_2_8_enexo | reg_act_config_inst_counter_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_26_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_cse
      & (reg_act_regs_data_0_7_enexo | reg_act_config_inst_regs_19_sva_dfm_6_enexo_8
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_8 | reg_act_config_inst_counter_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_27_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_9 | reg_act_config_inst_regs_19_sva_dfm_6_enexo_9
      | reg_act_config_inst_counter_enexo | reg_act_regs_data_1_6_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_28_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_10 | reg_act_config_inst_regs_19_sva_dfm_6_enexo_10
      | reg_act_regs_data_3_5_enexo | reg_act_config_inst_counter_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_29_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_cse
      & (reg_act_config_inst_regs_19_sva_dfm_6_enexo_11 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_11
      | reg_act_regs_data_2_4_enexo | reg_act_config_inst_counter_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_30_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_cse
      & (reg_act_config_inst_regs_19_sva_dfm_6_enexo_12 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_12
      | reg_act_regs_data_3_3_enexo | reg_act_config_inst_counter_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_31_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_13 | reg_act_config_inst_regs_19_sva_dfm_6_enexo_13
      | reg_act_regs_data_1_2_enexo | reg_act_config_inst_counter_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_32_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_14 | reg_act_regs_data_0_1_enexo
      | reg_act_config_inst_regs_19_sva_dfm_6_enexo_14 | reg_act_config_inst_counter_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_33_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_15 | reg_act_config_inst_regs_19_sva_dfm_6_enexo_15
      | reg_act_regs_data_1_0_enexo | reg_act_config_inst_counter_enexo);
  assign act_write_data_data_and_cse = ActUnitRun_wen & mux_tmp_1 & and_dcpl_1 &
      ActUnit_RunInst_switch_lp_nor_13_cse;
  assign done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct_mx0 = or_16_cse &
      and_dcpl_31 & (~ (operator_6_false_acc_tmp[5])) & is_start_sva & (~ (operator_8_false_acc_tmp[8]))
      & (~ act_config_InstIncr_if_if_unequal_tmp) & (fsm_output[2]);
  assign output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct_mx0 = is_start_sva
      & ActUnit_RunInst_switch_lp_equal_tmp_3 & (fsm_output[2]);
  assign rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct_mx0 = rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt) & (~ is_start_sva) & (fsm_output[2]);
  assign act_port_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct_mx0 = mux_tmp_16
      & and_dcpl_1 & (~ (act_config_in_InstFetch_mux_tmp[6])) & (act_config_in_InstFetch_mux_tmp[4])
      & (fsm_output[1]);
  assign ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_23_4_mx1_tmp_7_0
      = MUX_v_8_2_2((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:0]), reg_ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_23_4_ftd_12,
      is_start_sva);
  assign ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0 = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:8]==4'b1001));
  assign act_mem_banks_read_for_mux_mx0w0 = MUX_v_8_32_2(act_mem_banks_bank_array_impl_data0_0_127_120_sva_dfm,
      act_mem_banks_bank_array_impl_data0_1_127_120_sva_dfm, act_mem_banks_bank_array_impl_data0_2_127_120_sva_dfm,
      act_mem_banks_bank_array_impl_data0_3_127_120_sva_dfm, act_mem_banks_bank_array_impl_data0_4_127_120_sva_dfm,
      act_mem_banks_bank_array_impl_data0_5_127_120_sva_dfm, act_mem_banks_bank_array_impl_data0_6_127_120_sva_dfm,
      act_mem_banks_bank_array_impl_data0_7_127_120_sva_dfm, act_mem_banks_bank_array_impl_data0_8_127_120_sva_dfm,
      act_mem_banks_bank_array_impl_data0_9_127_120_sva_dfm, act_mem_banks_bank_array_impl_data0_10_127_120_sva_dfm,
      act_mem_banks_bank_array_impl_data0_11_127_120_sva_dfm, act_mem_banks_bank_array_impl_data0_12_127_120_sva_dfm,
      act_mem_banks_bank_array_impl_data0_13_127_120_sva_dfm, act_mem_banks_bank_array_impl_data0_14_127_120_sva_dfm,
      act_mem_banks_bank_array_impl_data0_15_127_120_sva_dfm, act_mem_banks_bank_array_impl_data0_16_127_120_sva_dfm,
      act_mem_banks_bank_array_impl_data0_17_127_120_sva_dfm, act_mem_banks_bank_array_impl_data0_18_127_120_sva_dfm,
      act_mem_banks_bank_array_impl_data0_19_127_120_sva_dfm, act_mem_banks_bank_array_impl_data0_20_127_120_sva_dfm,
      act_mem_banks_bank_array_impl_data0_21_127_120_sva_dfm, act_mem_banks_bank_array_impl_data0_22_127_120_sva_dfm,
      act_mem_banks_bank_array_impl_data0_23_127_120_sva_dfm, act_mem_banks_bank_array_impl_data0_24_127_120_sva_dfm,
      act_mem_banks_bank_array_impl_data0_25_127_120_sva_dfm, act_mem_banks_bank_array_impl_data0_26_127_120_sva_dfm,
      act_mem_banks_bank_array_impl_data0_27_127_120_sva_dfm, act_mem_banks_bank_array_impl_data0_28_127_120_sva_dfm,
      act_mem_banks_bank_array_impl_data0_29_127_120_sva_dfm, act_mem_banks_bank_array_impl_data0_30_127_120_sva_dfm,
      act_mem_banks_bank_array_impl_data0_31_127_120_sva_dfm, while_mux_124_ssc_mx0);
  assign act_mem_banks_read_for_mux_15_mx0w0 = MUX_v_8_32_2(act_mem_banks_bank_array_impl_data0_0_7_0_sva_dfm,
      act_mem_banks_bank_array_impl_data0_1_7_0_sva_dfm, act_mem_banks_bank_array_impl_data0_2_7_0_sva_dfm,
      act_mem_banks_bank_array_impl_data0_3_7_0_sva_dfm, act_mem_banks_bank_array_impl_data0_4_7_0_sva_dfm,
      act_mem_banks_bank_array_impl_data0_5_7_0_sva_dfm, act_mem_banks_bank_array_impl_data0_6_7_0_sva_dfm,
      act_mem_banks_bank_array_impl_data0_7_7_0_sva_dfm, act_mem_banks_bank_array_impl_data0_8_7_0_sva_dfm,
      act_mem_banks_bank_array_impl_data0_9_7_0_sva_dfm, act_mem_banks_bank_array_impl_data0_10_7_0_sva_dfm,
      act_mem_banks_bank_array_impl_data0_11_7_0_sva_dfm, act_mem_banks_bank_array_impl_data0_12_7_0_sva_dfm,
      act_mem_banks_bank_array_impl_data0_13_7_0_sva_dfm, act_mem_banks_bank_array_impl_data0_14_7_0_sva_dfm,
      act_mem_banks_bank_array_impl_data0_15_7_0_sva_dfm, act_mem_banks_bank_array_impl_data0_16_7_0_sva_dfm,
      act_mem_banks_bank_array_impl_data0_17_7_0_sva_dfm, act_mem_banks_bank_array_impl_data0_18_7_0_sva_dfm,
      act_mem_banks_bank_array_impl_data0_19_7_0_sva_dfm, act_mem_banks_bank_array_impl_data0_20_7_0_sva_dfm,
      act_mem_banks_bank_array_impl_data0_21_7_0_sva_dfm, act_mem_banks_bank_array_impl_data0_22_7_0_sva_dfm,
      act_mem_banks_bank_array_impl_data0_23_7_0_sva_dfm, act_mem_banks_bank_array_impl_data0_24_7_0_sva_dfm,
      act_mem_banks_bank_array_impl_data0_25_7_0_sva_dfm, act_mem_banks_bank_array_impl_data0_26_7_0_sva_dfm,
      act_mem_banks_bank_array_impl_data0_27_7_0_sva_dfm, act_mem_banks_bank_array_impl_data0_28_7_0_sva_dfm,
      act_mem_banks_bank_array_impl_data0_29_7_0_sva_dfm, act_mem_banks_bank_array_impl_data0_30_7_0_sva_dfm,
      act_mem_banks_bank_array_impl_data0_31_7_0_sva_dfm, while_mux_124_ssc_mx0);
  assign act_mem_banks_read_for_mux_1_mx0w0 = MUX_v_8_32_2(act_mem_banks_bank_array_impl_data0_0_119_112_sva_dfm,
      act_mem_banks_bank_array_impl_data0_1_119_112_sva_dfm, act_mem_banks_bank_array_impl_data0_2_119_112_sva_dfm,
      act_mem_banks_bank_array_impl_data0_3_119_112_sva_dfm, act_mem_banks_bank_array_impl_data0_4_119_112_sva_dfm,
      act_mem_banks_bank_array_impl_data0_5_119_112_sva_dfm, act_mem_banks_bank_array_impl_data0_6_119_112_sva_dfm,
      act_mem_banks_bank_array_impl_data0_7_119_112_sva_dfm, act_mem_banks_bank_array_impl_data0_8_119_112_sva_dfm,
      act_mem_banks_bank_array_impl_data0_9_119_112_sva_dfm, act_mem_banks_bank_array_impl_data0_10_119_112_sva_dfm,
      act_mem_banks_bank_array_impl_data0_11_119_112_sva_dfm, act_mem_banks_bank_array_impl_data0_12_119_112_sva_dfm,
      act_mem_banks_bank_array_impl_data0_13_119_112_sva_dfm, act_mem_banks_bank_array_impl_data0_14_119_112_sva_dfm,
      act_mem_banks_bank_array_impl_data0_15_119_112_sva_dfm, act_mem_banks_bank_array_impl_data0_16_119_112_sva_dfm,
      act_mem_banks_bank_array_impl_data0_17_119_112_sva_dfm, act_mem_banks_bank_array_impl_data0_18_119_112_sva_dfm,
      act_mem_banks_bank_array_impl_data0_19_119_112_sva_dfm, act_mem_banks_bank_array_impl_data0_20_119_112_sva_dfm,
      act_mem_banks_bank_array_impl_data0_21_119_112_sva_dfm, act_mem_banks_bank_array_impl_data0_22_119_112_sva_dfm,
      act_mem_banks_bank_array_impl_data0_23_119_112_sva_dfm, act_mem_banks_bank_array_impl_data0_24_119_112_sva_dfm,
      act_mem_banks_bank_array_impl_data0_25_119_112_sva_dfm, act_mem_banks_bank_array_impl_data0_26_119_112_sva_dfm,
      act_mem_banks_bank_array_impl_data0_27_119_112_sva_dfm, act_mem_banks_bank_array_impl_data0_28_119_112_sva_dfm,
      act_mem_banks_bank_array_impl_data0_29_119_112_sva_dfm, act_mem_banks_bank_array_impl_data0_30_119_112_sva_dfm,
      act_mem_banks_bank_array_impl_data0_31_119_112_sva_dfm, while_mux_124_ssc_mx0);
  assign act_mem_banks_read_for_mux_2_mx0w0 = MUX_v_8_32_2(act_mem_banks_bank_array_impl_data0_0_111_104_sva_dfm,
      act_mem_banks_bank_array_impl_data0_1_111_104_sva_dfm, act_mem_banks_bank_array_impl_data0_2_111_104_sva_dfm,
      act_mem_banks_bank_array_impl_data0_3_111_104_sva_dfm, act_mem_banks_bank_array_impl_data0_4_111_104_sva_dfm,
      act_mem_banks_bank_array_impl_data0_5_111_104_sva_dfm, act_mem_banks_bank_array_impl_data0_6_111_104_sva_dfm,
      act_mem_banks_bank_array_impl_data0_7_111_104_sva_dfm, act_mem_banks_bank_array_impl_data0_8_111_104_sva_dfm,
      act_mem_banks_bank_array_impl_data0_9_111_104_sva_dfm, act_mem_banks_bank_array_impl_data0_10_111_104_sva_dfm,
      act_mem_banks_bank_array_impl_data0_11_111_104_sva_dfm, act_mem_banks_bank_array_impl_data0_12_111_104_sva_dfm,
      act_mem_banks_bank_array_impl_data0_13_111_104_sva_dfm, act_mem_banks_bank_array_impl_data0_14_111_104_sva_dfm,
      act_mem_banks_bank_array_impl_data0_15_111_104_sva_dfm, act_mem_banks_bank_array_impl_data0_16_111_104_sva_dfm,
      act_mem_banks_bank_array_impl_data0_17_111_104_sva_dfm, act_mem_banks_bank_array_impl_data0_18_111_104_sva_dfm,
      act_mem_banks_bank_array_impl_data0_19_111_104_sva_dfm, act_mem_banks_bank_array_impl_data0_20_111_104_sva_dfm,
      act_mem_banks_bank_array_impl_data0_21_111_104_sva_dfm, act_mem_banks_bank_array_impl_data0_22_111_104_sva_dfm,
      act_mem_banks_bank_array_impl_data0_23_111_104_sva_dfm, act_mem_banks_bank_array_impl_data0_24_111_104_sva_dfm,
      act_mem_banks_bank_array_impl_data0_25_111_104_sva_dfm, act_mem_banks_bank_array_impl_data0_26_111_104_sva_dfm,
      act_mem_banks_bank_array_impl_data0_27_111_104_sva_dfm, act_mem_banks_bank_array_impl_data0_28_111_104_sva_dfm,
      act_mem_banks_bank_array_impl_data0_29_111_104_sva_dfm, act_mem_banks_bank_array_impl_data0_30_111_104_sva_dfm,
      act_mem_banks_bank_array_impl_data0_31_111_104_sva_dfm, while_mux_124_ssc_mx0);
  assign act_mem_banks_read_for_mux_14_mx0w0 = MUX_v_8_32_2(act_mem_banks_bank_array_impl_data0_0_15_8_sva_dfm,
      act_mem_banks_bank_array_impl_data0_1_15_8_sva_dfm, act_mem_banks_bank_array_impl_data0_2_15_8_sva_dfm,
      act_mem_banks_bank_array_impl_data0_3_15_8_sva_dfm, act_mem_banks_bank_array_impl_data0_4_15_8_sva_dfm,
      act_mem_banks_bank_array_impl_data0_5_15_8_sva_dfm, act_mem_banks_bank_array_impl_data0_6_15_8_sva_dfm,
      act_mem_banks_bank_array_impl_data0_7_15_8_sva_dfm, act_mem_banks_bank_array_impl_data0_8_15_8_sva_dfm,
      act_mem_banks_bank_array_impl_data0_9_15_8_sva_dfm, act_mem_banks_bank_array_impl_data0_10_15_8_sva_dfm,
      act_mem_banks_bank_array_impl_data0_11_15_8_sva_dfm, act_mem_banks_bank_array_impl_data0_12_15_8_sva_dfm,
      act_mem_banks_bank_array_impl_data0_13_15_8_sva_dfm, act_mem_banks_bank_array_impl_data0_14_15_8_sva_dfm,
      act_mem_banks_bank_array_impl_data0_15_15_8_sva_dfm, act_mem_banks_bank_array_impl_data0_16_15_8_sva_dfm,
      act_mem_banks_bank_array_impl_data0_17_15_8_sva_dfm, act_mem_banks_bank_array_impl_data0_18_15_8_sva_dfm,
      act_mem_banks_bank_array_impl_data0_19_15_8_sva_dfm, act_mem_banks_bank_array_impl_data0_20_15_8_sva_dfm,
      act_mem_banks_bank_array_impl_data0_21_15_8_sva_dfm, act_mem_banks_bank_array_impl_data0_22_15_8_sva_dfm,
      act_mem_banks_bank_array_impl_data0_23_15_8_sva_dfm, act_mem_banks_bank_array_impl_data0_24_15_8_sva_dfm,
      act_mem_banks_bank_array_impl_data0_25_15_8_sva_dfm, act_mem_banks_bank_array_impl_data0_26_15_8_sva_dfm,
      act_mem_banks_bank_array_impl_data0_27_15_8_sva_dfm, act_mem_banks_bank_array_impl_data0_28_15_8_sva_dfm,
      act_mem_banks_bank_array_impl_data0_29_15_8_sva_dfm, act_mem_banks_bank_array_impl_data0_30_15_8_sva_dfm,
      act_mem_banks_bank_array_impl_data0_31_15_8_sva_dfm, while_mux_124_ssc_mx0);
  assign act_mem_banks_read_for_mux_3_mx0w0 = MUX_v_8_32_2(act_mem_banks_bank_array_impl_data0_0_103_96_sva_dfm,
      act_mem_banks_bank_array_impl_data0_1_103_96_sva_dfm, act_mem_banks_bank_array_impl_data0_2_103_96_sva_dfm,
      act_mem_banks_bank_array_impl_data0_3_103_96_sva_dfm, act_mem_banks_bank_array_impl_data0_4_103_96_sva_dfm,
      act_mem_banks_bank_array_impl_data0_5_103_96_sva_dfm, act_mem_banks_bank_array_impl_data0_6_103_96_sva_dfm,
      act_mem_banks_bank_array_impl_data0_7_103_96_sva_dfm, act_mem_banks_bank_array_impl_data0_8_103_96_sva_dfm,
      act_mem_banks_bank_array_impl_data0_9_103_96_sva_dfm, act_mem_banks_bank_array_impl_data0_10_103_96_sva_dfm,
      act_mem_banks_bank_array_impl_data0_11_103_96_sva_dfm, act_mem_banks_bank_array_impl_data0_12_103_96_sva_dfm,
      act_mem_banks_bank_array_impl_data0_13_103_96_sva_dfm, act_mem_banks_bank_array_impl_data0_14_103_96_sva_dfm,
      act_mem_banks_bank_array_impl_data0_15_103_96_sva_dfm, act_mem_banks_bank_array_impl_data0_16_103_96_sva_dfm,
      act_mem_banks_bank_array_impl_data0_17_103_96_sva_dfm, act_mem_banks_bank_array_impl_data0_18_103_96_sva_dfm,
      act_mem_banks_bank_array_impl_data0_19_103_96_sva_dfm, act_mem_banks_bank_array_impl_data0_20_103_96_sva_dfm,
      act_mem_banks_bank_array_impl_data0_21_103_96_sva_dfm, act_mem_banks_bank_array_impl_data0_22_103_96_sva_dfm,
      act_mem_banks_bank_array_impl_data0_23_103_96_sva_dfm, act_mem_banks_bank_array_impl_data0_24_103_96_sva_dfm,
      act_mem_banks_bank_array_impl_data0_25_103_96_sva_dfm, act_mem_banks_bank_array_impl_data0_26_103_96_sva_dfm,
      act_mem_banks_bank_array_impl_data0_27_103_96_sva_dfm, act_mem_banks_bank_array_impl_data0_28_103_96_sva_dfm,
      act_mem_banks_bank_array_impl_data0_29_103_96_sva_dfm, act_mem_banks_bank_array_impl_data0_30_103_96_sva_dfm,
      act_mem_banks_bank_array_impl_data0_31_103_96_sva_dfm, while_mux_124_ssc_mx0);
  assign act_mem_banks_read_for_mux_4_mx0w0 = MUX_v_8_32_2(act_mem_banks_bank_array_impl_data0_0_95_88_sva_dfm,
      act_mem_banks_bank_array_impl_data0_1_95_88_sva_dfm, act_mem_banks_bank_array_impl_data0_2_95_88_sva_dfm,
      act_mem_banks_bank_array_impl_data0_3_95_88_sva_dfm, act_mem_banks_bank_array_impl_data0_4_95_88_sva_dfm,
      act_mem_banks_bank_array_impl_data0_5_95_88_sva_dfm, act_mem_banks_bank_array_impl_data0_6_95_88_sva_dfm,
      act_mem_banks_bank_array_impl_data0_7_95_88_sva_dfm, act_mem_banks_bank_array_impl_data0_8_95_88_sva_dfm,
      act_mem_banks_bank_array_impl_data0_9_95_88_sva_dfm, act_mem_banks_bank_array_impl_data0_10_95_88_sva_dfm,
      act_mem_banks_bank_array_impl_data0_11_95_88_sva_dfm, act_mem_banks_bank_array_impl_data0_12_95_88_sva_dfm,
      act_mem_banks_bank_array_impl_data0_13_95_88_sva_dfm, act_mem_banks_bank_array_impl_data0_14_95_88_sva_dfm,
      act_mem_banks_bank_array_impl_data0_15_95_88_sva_dfm, act_mem_banks_bank_array_impl_data0_16_95_88_sva_dfm,
      act_mem_banks_bank_array_impl_data0_17_95_88_sva_dfm, act_mem_banks_bank_array_impl_data0_18_95_88_sva_dfm,
      act_mem_banks_bank_array_impl_data0_19_95_88_sva_dfm, act_mem_banks_bank_array_impl_data0_20_95_88_sva_dfm,
      act_mem_banks_bank_array_impl_data0_21_95_88_sva_dfm, act_mem_banks_bank_array_impl_data0_22_95_88_sva_dfm,
      act_mem_banks_bank_array_impl_data0_23_95_88_sva_dfm, act_mem_banks_bank_array_impl_data0_24_95_88_sva_dfm,
      act_mem_banks_bank_array_impl_data0_25_95_88_sva_dfm, act_mem_banks_bank_array_impl_data0_26_95_88_sva_dfm,
      act_mem_banks_bank_array_impl_data0_27_95_88_sva_dfm, act_mem_banks_bank_array_impl_data0_28_95_88_sva_dfm,
      act_mem_banks_bank_array_impl_data0_29_95_88_sva_dfm, act_mem_banks_bank_array_impl_data0_30_95_88_sva_dfm,
      act_mem_banks_bank_array_impl_data0_31_95_88_sva_dfm, while_mux_124_ssc_mx0);
  assign act_mem_banks_read_for_mux_13_mx0w0 = MUX_v_8_32_2(act_mem_banks_bank_array_impl_data0_0_23_16_sva_dfm,
      act_mem_banks_bank_array_impl_data0_1_23_16_sva_dfm, act_mem_banks_bank_array_impl_data0_2_23_16_sva_dfm,
      act_mem_banks_bank_array_impl_data0_3_23_16_sva_dfm, act_mem_banks_bank_array_impl_data0_4_23_16_sva_dfm,
      act_mem_banks_bank_array_impl_data0_5_23_16_sva_dfm, act_mem_banks_bank_array_impl_data0_6_23_16_sva_dfm,
      act_mem_banks_bank_array_impl_data0_7_23_16_sva_dfm, act_mem_banks_bank_array_impl_data0_8_23_16_sva_dfm,
      act_mem_banks_bank_array_impl_data0_9_23_16_sva_dfm, act_mem_banks_bank_array_impl_data0_10_23_16_sva_dfm,
      act_mem_banks_bank_array_impl_data0_11_23_16_sva_dfm, act_mem_banks_bank_array_impl_data0_12_23_16_sva_dfm,
      act_mem_banks_bank_array_impl_data0_13_23_16_sva_dfm, act_mem_banks_bank_array_impl_data0_14_23_16_sva_dfm,
      act_mem_banks_bank_array_impl_data0_15_23_16_sva_dfm, act_mem_banks_bank_array_impl_data0_16_23_16_sva_dfm,
      act_mem_banks_bank_array_impl_data0_17_23_16_sva_dfm, act_mem_banks_bank_array_impl_data0_18_23_16_sva_dfm,
      act_mem_banks_bank_array_impl_data0_19_23_16_sva_dfm, act_mem_banks_bank_array_impl_data0_20_23_16_sva_dfm,
      act_mem_banks_bank_array_impl_data0_21_23_16_sva_dfm, act_mem_banks_bank_array_impl_data0_22_23_16_sva_dfm,
      act_mem_banks_bank_array_impl_data0_23_23_16_sva_dfm, act_mem_banks_bank_array_impl_data0_24_23_16_sva_dfm,
      act_mem_banks_bank_array_impl_data0_25_23_16_sva_dfm, act_mem_banks_bank_array_impl_data0_26_23_16_sva_dfm,
      act_mem_banks_bank_array_impl_data0_27_23_16_sva_dfm, act_mem_banks_bank_array_impl_data0_28_23_16_sva_dfm,
      act_mem_banks_bank_array_impl_data0_29_23_16_sva_dfm, act_mem_banks_bank_array_impl_data0_30_23_16_sva_dfm,
      act_mem_banks_bank_array_impl_data0_31_23_16_sva_dfm, while_mux_124_ssc_mx0);
  assign act_mem_banks_read_for_mux_5_mx0w0 = MUX_v_8_32_2(act_mem_banks_bank_array_impl_data0_0_87_80_sva_dfm,
      act_mem_banks_bank_array_impl_data0_1_87_80_sva_dfm, act_mem_banks_bank_array_impl_data0_2_87_80_sva_dfm,
      act_mem_banks_bank_array_impl_data0_3_87_80_sva_dfm, act_mem_banks_bank_array_impl_data0_4_87_80_sva_dfm,
      act_mem_banks_bank_array_impl_data0_5_87_80_sva_dfm, act_mem_banks_bank_array_impl_data0_6_87_80_sva_dfm,
      act_mem_banks_bank_array_impl_data0_7_87_80_sva_dfm, act_mem_banks_bank_array_impl_data0_8_87_80_sva_dfm,
      act_mem_banks_bank_array_impl_data0_9_87_80_sva_dfm, act_mem_banks_bank_array_impl_data0_10_87_80_sva_dfm,
      act_mem_banks_bank_array_impl_data0_11_87_80_sva_dfm, act_mem_banks_bank_array_impl_data0_12_87_80_sva_dfm,
      act_mem_banks_bank_array_impl_data0_13_87_80_sva_dfm, act_mem_banks_bank_array_impl_data0_14_87_80_sva_dfm,
      act_mem_banks_bank_array_impl_data0_15_87_80_sva_dfm, act_mem_banks_bank_array_impl_data0_16_87_80_sva_dfm,
      act_mem_banks_bank_array_impl_data0_17_87_80_sva_dfm, act_mem_banks_bank_array_impl_data0_18_87_80_sva_dfm,
      act_mem_banks_bank_array_impl_data0_19_87_80_sva_dfm, act_mem_banks_bank_array_impl_data0_20_87_80_sva_dfm,
      act_mem_banks_bank_array_impl_data0_21_87_80_sva_dfm, act_mem_banks_bank_array_impl_data0_22_87_80_sva_dfm,
      act_mem_banks_bank_array_impl_data0_23_87_80_sva_dfm, act_mem_banks_bank_array_impl_data0_24_87_80_sva_dfm,
      act_mem_banks_bank_array_impl_data0_25_87_80_sva_dfm, act_mem_banks_bank_array_impl_data0_26_87_80_sva_dfm,
      act_mem_banks_bank_array_impl_data0_27_87_80_sva_dfm, act_mem_banks_bank_array_impl_data0_28_87_80_sva_dfm,
      act_mem_banks_bank_array_impl_data0_29_87_80_sva_dfm, act_mem_banks_bank_array_impl_data0_30_87_80_sva_dfm,
      act_mem_banks_bank_array_impl_data0_31_87_80_sva_dfm, while_mux_124_ssc_mx0);
  assign act_mem_banks_read_for_mux_6_mx0w0 = MUX_v_8_32_2(act_mem_banks_bank_array_impl_data0_0_79_72_sva_dfm,
      act_mem_banks_bank_array_impl_data0_1_79_72_sva_dfm, act_mem_banks_bank_array_impl_data0_2_79_72_sva_dfm,
      act_mem_banks_bank_array_impl_data0_3_79_72_sva_dfm, act_mem_banks_bank_array_impl_data0_4_79_72_sva_dfm,
      act_mem_banks_bank_array_impl_data0_5_79_72_sva_dfm, act_mem_banks_bank_array_impl_data0_6_79_72_sva_dfm,
      act_mem_banks_bank_array_impl_data0_7_79_72_sva_dfm, act_mem_banks_bank_array_impl_data0_8_79_72_sva_dfm,
      act_mem_banks_bank_array_impl_data0_9_79_72_sva_dfm, act_mem_banks_bank_array_impl_data0_10_79_72_sva_dfm,
      act_mem_banks_bank_array_impl_data0_11_79_72_sva_dfm, act_mem_banks_bank_array_impl_data0_12_79_72_sva_dfm,
      act_mem_banks_bank_array_impl_data0_13_79_72_sva_dfm, act_mem_banks_bank_array_impl_data0_14_79_72_sva_dfm,
      act_mem_banks_bank_array_impl_data0_15_79_72_sva_dfm, act_mem_banks_bank_array_impl_data0_16_79_72_sva_dfm,
      act_mem_banks_bank_array_impl_data0_17_79_72_sva_dfm, act_mem_banks_bank_array_impl_data0_18_79_72_sva_dfm,
      act_mem_banks_bank_array_impl_data0_19_79_72_sva_dfm, act_mem_banks_bank_array_impl_data0_20_79_72_sva_dfm,
      act_mem_banks_bank_array_impl_data0_21_79_72_sva_dfm, act_mem_banks_bank_array_impl_data0_22_79_72_sva_dfm,
      act_mem_banks_bank_array_impl_data0_23_79_72_sva_dfm, act_mem_banks_bank_array_impl_data0_24_79_72_sva_dfm,
      act_mem_banks_bank_array_impl_data0_25_79_72_sva_dfm, act_mem_banks_bank_array_impl_data0_26_79_72_sva_dfm,
      act_mem_banks_bank_array_impl_data0_27_79_72_sva_dfm, act_mem_banks_bank_array_impl_data0_28_79_72_sva_dfm,
      act_mem_banks_bank_array_impl_data0_29_79_72_sva_dfm, act_mem_banks_bank_array_impl_data0_30_79_72_sva_dfm,
      act_mem_banks_bank_array_impl_data0_31_79_72_sva_dfm, while_mux_124_ssc_mx0);
  assign act_mem_banks_read_for_mux_12_mx0w0 = MUX_v_8_32_2(act_mem_banks_bank_array_impl_data0_0_31_24_sva_dfm,
      act_mem_banks_bank_array_impl_data0_1_31_24_sva_dfm, act_mem_banks_bank_array_impl_data0_2_31_24_sva_dfm,
      act_mem_banks_bank_array_impl_data0_3_31_24_sva_dfm, act_mem_banks_bank_array_impl_data0_4_31_24_sva_dfm,
      act_mem_banks_bank_array_impl_data0_5_31_24_sva_dfm, act_mem_banks_bank_array_impl_data0_6_31_24_sva_dfm,
      act_mem_banks_bank_array_impl_data0_7_31_24_sva_dfm, act_mem_banks_bank_array_impl_data0_8_31_24_sva_dfm,
      act_mem_banks_bank_array_impl_data0_9_31_24_sva_dfm, act_mem_banks_bank_array_impl_data0_10_31_24_sva_dfm,
      act_mem_banks_bank_array_impl_data0_11_31_24_sva_dfm, act_mem_banks_bank_array_impl_data0_12_31_24_sva_dfm,
      act_mem_banks_bank_array_impl_data0_13_31_24_sva_dfm, act_mem_banks_bank_array_impl_data0_14_31_24_sva_dfm,
      act_mem_banks_bank_array_impl_data0_15_31_24_sva_dfm, act_mem_banks_bank_array_impl_data0_16_31_24_sva_dfm,
      act_mem_banks_bank_array_impl_data0_17_31_24_sva_dfm, act_mem_banks_bank_array_impl_data0_18_31_24_sva_dfm,
      act_mem_banks_bank_array_impl_data0_19_31_24_sva_dfm, act_mem_banks_bank_array_impl_data0_20_31_24_sva_dfm,
      act_mem_banks_bank_array_impl_data0_21_31_24_sva_dfm, act_mem_banks_bank_array_impl_data0_22_31_24_sva_dfm,
      act_mem_banks_bank_array_impl_data0_23_31_24_sva_dfm, act_mem_banks_bank_array_impl_data0_24_31_24_sva_dfm,
      act_mem_banks_bank_array_impl_data0_25_31_24_sva_dfm, act_mem_banks_bank_array_impl_data0_26_31_24_sva_dfm,
      act_mem_banks_bank_array_impl_data0_27_31_24_sva_dfm, act_mem_banks_bank_array_impl_data0_28_31_24_sva_dfm,
      act_mem_banks_bank_array_impl_data0_29_31_24_sva_dfm, act_mem_banks_bank_array_impl_data0_30_31_24_sva_dfm,
      act_mem_banks_bank_array_impl_data0_31_31_24_sva_dfm, while_mux_124_ssc_mx0);
  assign act_mem_banks_read_for_mux_7_mx0w0 = MUX_v_8_32_2(act_mem_banks_bank_array_impl_data0_0_71_64_sva_dfm,
      act_mem_banks_bank_array_impl_data0_1_71_64_sva_dfm, act_mem_banks_bank_array_impl_data0_2_71_64_sva_dfm,
      act_mem_banks_bank_array_impl_data0_3_71_64_sva_dfm, act_mem_banks_bank_array_impl_data0_4_71_64_sva_dfm,
      act_mem_banks_bank_array_impl_data0_5_71_64_sva_dfm, act_mem_banks_bank_array_impl_data0_6_71_64_sva_dfm,
      act_mem_banks_bank_array_impl_data0_7_71_64_sva_dfm, act_mem_banks_bank_array_impl_data0_8_71_64_sva_dfm,
      act_mem_banks_bank_array_impl_data0_9_71_64_sva_dfm, act_mem_banks_bank_array_impl_data0_10_71_64_sva_dfm,
      act_mem_banks_bank_array_impl_data0_11_71_64_sva_dfm, act_mem_banks_bank_array_impl_data0_12_71_64_sva_dfm,
      act_mem_banks_bank_array_impl_data0_13_71_64_sva_dfm, act_mem_banks_bank_array_impl_data0_14_71_64_sva_dfm,
      act_mem_banks_bank_array_impl_data0_15_71_64_sva_dfm, act_mem_banks_bank_array_impl_data0_16_71_64_sva_dfm,
      act_mem_banks_bank_array_impl_data0_17_71_64_sva_dfm, act_mem_banks_bank_array_impl_data0_18_71_64_sva_dfm,
      act_mem_banks_bank_array_impl_data0_19_71_64_sva_dfm, act_mem_banks_bank_array_impl_data0_20_71_64_sva_dfm,
      act_mem_banks_bank_array_impl_data0_21_71_64_sva_dfm, act_mem_banks_bank_array_impl_data0_22_71_64_sva_dfm,
      act_mem_banks_bank_array_impl_data0_23_71_64_sva_dfm, act_mem_banks_bank_array_impl_data0_24_71_64_sva_dfm,
      act_mem_banks_bank_array_impl_data0_25_71_64_sva_dfm, act_mem_banks_bank_array_impl_data0_26_71_64_sva_dfm,
      act_mem_banks_bank_array_impl_data0_27_71_64_sva_dfm, act_mem_banks_bank_array_impl_data0_28_71_64_sva_dfm,
      act_mem_banks_bank_array_impl_data0_29_71_64_sva_dfm, act_mem_banks_bank_array_impl_data0_30_71_64_sva_dfm,
      act_mem_banks_bank_array_impl_data0_31_71_64_sva_dfm, while_mux_124_ssc_mx0);
  assign act_mem_banks_read_for_mux_8_mx0w0 = MUX_v_8_32_2(act_mem_banks_bank_array_impl_data0_0_63_56_sva_dfm,
      act_mem_banks_bank_array_impl_data0_1_63_56_sva_dfm, act_mem_banks_bank_array_impl_data0_2_63_56_sva_dfm,
      act_mem_banks_bank_array_impl_data0_3_63_56_sva_dfm, act_mem_banks_bank_array_impl_data0_4_63_56_sva_dfm,
      act_mem_banks_bank_array_impl_data0_5_63_56_sva_dfm, act_mem_banks_bank_array_impl_data0_6_63_56_sva_dfm,
      act_mem_banks_bank_array_impl_data0_7_63_56_sva_dfm, act_mem_banks_bank_array_impl_data0_8_63_56_sva_dfm,
      act_mem_banks_bank_array_impl_data0_9_63_56_sva_dfm, act_mem_banks_bank_array_impl_data0_10_63_56_sva_dfm,
      act_mem_banks_bank_array_impl_data0_11_63_56_sva_dfm, act_mem_banks_bank_array_impl_data0_12_63_56_sva_dfm,
      act_mem_banks_bank_array_impl_data0_13_63_56_sva_dfm, act_mem_banks_bank_array_impl_data0_14_63_56_sva_dfm,
      act_mem_banks_bank_array_impl_data0_15_63_56_sva_dfm, act_mem_banks_bank_array_impl_data0_16_63_56_sva_dfm,
      act_mem_banks_bank_array_impl_data0_17_63_56_sva_dfm, act_mem_banks_bank_array_impl_data0_18_63_56_sva_dfm,
      act_mem_banks_bank_array_impl_data0_19_63_56_sva_dfm, act_mem_banks_bank_array_impl_data0_20_63_56_sva_dfm,
      act_mem_banks_bank_array_impl_data0_21_63_56_sva_dfm, act_mem_banks_bank_array_impl_data0_22_63_56_sva_dfm,
      act_mem_banks_bank_array_impl_data0_23_63_56_sva_dfm, act_mem_banks_bank_array_impl_data0_24_63_56_sva_dfm,
      act_mem_banks_bank_array_impl_data0_25_63_56_sva_dfm, act_mem_banks_bank_array_impl_data0_26_63_56_sva_dfm,
      act_mem_banks_bank_array_impl_data0_27_63_56_sva_dfm, act_mem_banks_bank_array_impl_data0_28_63_56_sva_dfm,
      act_mem_banks_bank_array_impl_data0_29_63_56_sva_dfm, act_mem_banks_bank_array_impl_data0_30_63_56_sva_dfm,
      act_mem_banks_bank_array_impl_data0_31_63_56_sva_dfm, while_mux_124_ssc_mx0);
  assign act_mem_banks_read_for_mux_11_mx0w0 = MUX_v_8_32_2(act_mem_banks_bank_array_impl_data0_0_39_32_sva_dfm,
      act_mem_banks_bank_array_impl_data0_1_39_32_sva_dfm, act_mem_banks_bank_array_impl_data0_2_39_32_sva_dfm,
      act_mem_banks_bank_array_impl_data0_3_39_32_sva_dfm, act_mem_banks_bank_array_impl_data0_4_39_32_sva_dfm,
      act_mem_banks_bank_array_impl_data0_5_39_32_sva_dfm, act_mem_banks_bank_array_impl_data0_6_39_32_sva_dfm,
      act_mem_banks_bank_array_impl_data0_7_39_32_sva_dfm, act_mem_banks_bank_array_impl_data0_8_39_32_sva_dfm,
      act_mem_banks_bank_array_impl_data0_9_39_32_sva_dfm, act_mem_banks_bank_array_impl_data0_10_39_32_sva_dfm,
      act_mem_banks_bank_array_impl_data0_11_39_32_sva_dfm, act_mem_banks_bank_array_impl_data0_12_39_32_sva_dfm,
      act_mem_banks_bank_array_impl_data0_13_39_32_sva_dfm, act_mem_banks_bank_array_impl_data0_14_39_32_sva_dfm,
      act_mem_banks_bank_array_impl_data0_15_39_32_sva_dfm, act_mem_banks_bank_array_impl_data0_16_39_32_sva_dfm,
      act_mem_banks_bank_array_impl_data0_17_39_32_sva_dfm, act_mem_banks_bank_array_impl_data0_18_39_32_sva_dfm,
      act_mem_banks_bank_array_impl_data0_19_39_32_sva_dfm, act_mem_banks_bank_array_impl_data0_20_39_32_sva_dfm,
      act_mem_banks_bank_array_impl_data0_21_39_32_sva_dfm, act_mem_banks_bank_array_impl_data0_22_39_32_sva_dfm,
      act_mem_banks_bank_array_impl_data0_23_39_32_sva_dfm, act_mem_banks_bank_array_impl_data0_24_39_32_sva_dfm,
      act_mem_banks_bank_array_impl_data0_25_39_32_sva_dfm, act_mem_banks_bank_array_impl_data0_26_39_32_sva_dfm,
      act_mem_banks_bank_array_impl_data0_27_39_32_sva_dfm, act_mem_banks_bank_array_impl_data0_28_39_32_sva_dfm,
      act_mem_banks_bank_array_impl_data0_29_39_32_sva_dfm, act_mem_banks_bank_array_impl_data0_30_39_32_sva_dfm,
      act_mem_banks_bank_array_impl_data0_31_39_32_sva_dfm, while_mux_124_ssc_mx0);
  assign act_mem_banks_read_for_mux_9_mx0w0 = MUX_v_8_32_2(act_mem_banks_bank_array_impl_data0_0_55_48_sva_dfm,
      act_mem_banks_bank_array_impl_data0_1_55_48_sva_dfm, act_mem_banks_bank_array_impl_data0_2_55_48_sva_dfm,
      act_mem_banks_bank_array_impl_data0_3_55_48_sva_dfm, act_mem_banks_bank_array_impl_data0_4_55_48_sva_dfm,
      act_mem_banks_bank_array_impl_data0_5_55_48_sva_dfm, act_mem_banks_bank_array_impl_data0_6_55_48_sva_dfm,
      act_mem_banks_bank_array_impl_data0_7_55_48_sva_dfm, act_mem_banks_bank_array_impl_data0_8_55_48_sva_dfm,
      act_mem_banks_bank_array_impl_data0_9_55_48_sva_dfm, act_mem_banks_bank_array_impl_data0_10_55_48_sva_dfm,
      act_mem_banks_bank_array_impl_data0_11_55_48_sva_dfm, act_mem_banks_bank_array_impl_data0_12_55_48_sva_dfm,
      act_mem_banks_bank_array_impl_data0_13_55_48_sva_dfm, act_mem_banks_bank_array_impl_data0_14_55_48_sva_dfm,
      act_mem_banks_bank_array_impl_data0_15_55_48_sva_dfm, act_mem_banks_bank_array_impl_data0_16_55_48_sva_dfm,
      act_mem_banks_bank_array_impl_data0_17_55_48_sva_dfm, act_mem_banks_bank_array_impl_data0_18_55_48_sva_dfm,
      act_mem_banks_bank_array_impl_data0_19_55_48_sva_dfm, act_mem_banks_bank_array_impl_data0_20_55_48_sva_dfm,
      act_mem_banks_bank_array_impl_data0_21_55_48_sva_dfm, act_mem_banks_bank_array_impl_data0_22_55_48_sva_dfm,
      act_mem_banks_bank_array_impl_data0_23_55_48_sva_dfm, act_mem_banks_bank_array_impl_data0_24_55_48_sva_dfm,
      act_mem_banks_bank_array_impl_data0_25_55_48_sva_dfm, act_mem_banks_bank_array_impl_data0_26_55_48_sva_dfm,
      act_mem_banks_bank_array_impl_data0_27_55_48_sva_dfm, act_mem_banks_bank_array_impl_data0_28_55_48_sva_dfm,
      act_mem_banks_bank_array_impl_data0_29_55_48_sva_dfm, act_mem_banks_bank_array_impl_data0_30_55_48_sva_dfm,
      act_mem_banks_bank_array_impl_data0_31_55_48_sva_dfm, while_mux_124_ssc_mx0);
  assign act_mem_banks_read_for_mux_10_mx0w0 = MUX_v_8_32_2(act_mem_banks_bank_array_impl_data0_0_47_40_sva_dfm,
      act_mem_banks_bank_array_impl_data0_1_47_40_sva_dfm, act_mem_banks_bank_array_impl_data0_2_47_40_sva_dfm,
      act_mem_banks_bank_array_impl_data0_3_47_40_sva_dfm, act_mem_banks_bank_array_impl_data0_4_47_40_sva_dfm,
      act_mem_banks_bank_array_impl_data0_5_47_40_sva_dfm, act_mem_banks_bank_array_impl_data0_6_47_40_sva_dfm,
      act_mem_banks_bank_array_impl_data0_7_47_40_sva_dfm, act_mem_banks_bank_array_impl_data0_8_47_40_sva_dfm,
      act_mem_banks_bank_array_impl_data0_9_47_40_sva_dfm, act_mem_banks_bank_array_impl_data0_10_47_40_sva_dfm,
      act_mem_banks_bank_array_impl_data0_11_47_40_sva_dfm, act_mem_banks_bank_array_impl_data0_12_47_40_sva_dfm,
      act_mem_banks_bank_array_impl_data0_13_47_40_sva_dfm, act_mem_banks_bank_array_impl_data0_14_47_40_sva_dfm,
      act_mem_banks_bank_array_impl_data0_15_47_40_sva_dfm, act_mem_banks_bank_array_impl_data0_16_47_40_sva_dfm,
      act_mem_banks_bank_array_impl_data0_17_47_40_sva_dfm, act_mem_banks_bank_array_impl_data0_18_47_40_sva_dfm,
      act_mem_banks_bank_array_impl_data0_19_47_40_sva_dfm, act_mem_banks_bank_array_impl_data0_20_47_40_sva_dfm,
      act_mem_banks_bank_array_impl_data0_21_47_40_sva_dfm, act_mem_banks_bank_array_impl_data0_22_47_40_sva_dfm,
      act_mem_banks_bank_array_impl_data0_23_47_40_sva_dfm, act_mem_banks_bank_array_impl_data0_24_47_40_sva_dfm,
      act_mem_banks_bank_array_impl_data0_25_47_40_sva_dfm, act_mem_banks_bank_array_impl_data0_26_47_40_sva_dfm,
      act_mem_banks_bank_array_impl_data0_27_47_40_sva_dfm, act_mem_banks_bank_array_impl_data0_28_47_40_sva_dfm,
      act_mem_banks_bank_array_impl_data0_29_47_40_sva_dfm, act_mem_banks_bank_array_impl_data0_30_47_40_sva_dfm,
      act_mem_banks_bank_array_impl_data0_31_47_40_sva_dfm, while_mux_124_ssc_mx0);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_3_mx0w2 = act_read_addrs_lpi_1_dfm_9
      & ({{4{ActUnit_DecodeAxiRead_unequal_tmp_1}}, ActUnit_DecodeAxiRead_unequal_tmp_1})
      & ({{4{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt})
      & ({{4{rva_in_PopNB_mioi_return_rsc_z_mxwt}}, rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_cse_1 = ~(ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0
      | ActUnit_RunInst_switch_lp_equal_tmp_11 | ActUnit_RunInst_switch_lp_equal_tmp_12
      | ActUnit_RunInst_switch_lp_equal_tmp_13 | ActUnit_RunInst_switch_lp_equal_tmp_14
      | ActUnit_RunInst_switch_lp_equal_tmp_15 | ActUnit_RunInst_switch_lp_equal_tmp_16
      | ActUnit_RunInst_switch_lp_equal_tmp_17 | ActUnit_RunInst_switch_lp_equal_tmp_18
      | ActUnit_RunInst_switch_lp_equal_tmp_19 | ActUnit_RunInst_switch_lp_nor_tmp_1);
  assign ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0 = (act_config_in_InstFetch_mux_tmp[7:4]==4'b0010);
  assign ActUnit_RunInst_switch_lp_nor_7_itm_mx0w0 = ~((act_config_in_InstFetch_mux_tmp[7:5]!=3'b000));
  assign act_config_in_InstFetch_mux_tmp = MUX_v_8_32_2(act_config_inst_regs_0_sva_dfm_5,
      act_config_inst_regs_1_sva_dfm_5, act_config_inst_regs_2_sva_dfm_5, act_config_inst_regs_3_sva_dfm_5,
      act_config_inst_regs_4_sva_dfm_5, act_config_inst_regs_5_sva_dfm_5, act_config_inst_regs_6_sva_dfm_5,
      act_config_inst_regs_7_sva_dfm_5, act_config_inst_regs_8_sva_dfm_5, act_config_inst_regs_9_sva_dfm_5,
      act_config_inst_regs_10_sva_dfm_5, act_config_inst_regs_11_sva_dfm_5, act_config_inst_regs_12_sva_dfm_5,
      act_config_inst_regs_13_sva_dfm_5, act_config_inst_regs_14_sva_dfm_5, act_config_inst_regs_15_sva_dfm_5,
      act_config_inst_regs_16_sva_dfm_6, act_config_inst_regs_17_sva_dfm_6, act_config_inst_regs_18_sva_dfm_6,
      act_config_inst_regs_19_sva_dfm_6, act_config_inst_regs_20_sva_dfm_6, act_config_inst_regs_21_sva_dfm_6,
      act_config_inst_regs_22_sva_dfm_6, act_config_inst_regs_23_sva_dfm_6, act_config_inst_regs_24_sva_dfm_6,
      act_config_inst_regs_25_sva_dfm_6, act_config_inst_regs_26_sva_dfm_6, act_config_inst_regs_27_sva_dfm_6,
      act_config_inst_regs_28_sva_dfm_6, act_config_inst_regs_29_sva_dfm_6, act_config_inst_regs_30_sva_dfm_6,
      act_config_inst_regs_31_sva_dfm_6, act_config_inst_counter_sva);
  assign ActUnit_RunInst_switch_lp_equal_tmp_11 = (act_config_in_InstFetch_mux_tmp[7:4]==4'b0011);
  assign ActUnit_RunInst_switch_lp_equal_tmp_12 = (act_config_in_InstFetch_mux_tmp[7:4]==4'b0100);
  assign ActUnit_RunInst_switch_lp_equal_tmp_13 = (act_config_in_InstFetch_mux_tmp[7:4]==4'b0111);
  assign ActUnit_RunInst_switch_lp_equal_tmp_14 = (act_config_in_InstFetch_mux_tmp[7:4]==4'b1000);
  assign ActUnit_RunInst_switch_lp_equal_tmp_15 = (act_config_in_InstFetch_mux_tmp[7:4]==4'b1001);
  assign ActUnit_RunInst_switch_lp_nor_13_cse = ~((act_config_in_InstFetch_mux_tmp[6])
      | (act_config_in_InstFetch_mux_tmp[4]));
  assign ActUnit_RunInst_switch_lp_equal_tmp_16 = (act_config_in_InstFetch_mux_tmp[7])
      & (act_config_in_InstFetch_mux_tmp[5]) & ActUnit_RunInst_switch_lp_nor_13_cse;
  assign ActUnit_RunInst_switch_lp_equal_tmp_17 = (act_config_in_InstFetch_mux_tmp[7:4]==4'b1011);
  assign ActUnit_RunInst_switch_lp_equal_tmp_18 = (act_config_in_InstFetch_mux_tmp[7:4]==4'b1100);
  assign ActUnit_RunInst_switch_lp_equal_tmp_19 = (act_config_in_InstFetch_mux_tmp[7:4]==4'b1101);
  assign ActUnit_RunInst_switch_lp_nor_tmp_1 = ~(((act_config_in_InstFetch_mux_tmp[4])
      & ActUnit_RunInst_switch_lp_nor_7_itm_mx0w0) | ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0
      | ActUnit_RunInst_switch_lp_equal_tmp_11 | ActUnit_RunInst_switch_lp_equal_tmp_12
      | ActUnit_RunInst_switch_lp_equal_tmp_13 | ActUnit_RunInst_switch_lp_equal_tmp_14
      | ActUnit_RunInst_switch_lp_equal_tmp_15 | ActUnit_RunInst_switch_lp_equal_tmp_16
      | ActUnit_RunInst_switch_lp_equal_tmp_17 | ActUnit_RunInst_switch_lp_equal_tmp_18
      | ActUnit_RunInst_switch_lp_equal_tmp_19);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      = MUX_v_20_4_2(act_regs_data_0_15_sva, act_regs_data_1_15_sva, act_regs_data_2_15_sva,
      act_regs_data_3_15_sva, act_config_in_InstFetch_mux_tmp[1:0]);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      = MUX_v_20_4_2(act_regs_data_0_14_sva, act_regs_data_1_14_sva, act_regs_data_2_14_sva,
      act_regs_data_3_14_sva, act_config_in_InstFetch_mux_tmp[1:0]);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      = MUX_v_20_4_2(act_regs_data_0_13_sva, act_regs_data_1_13_sva, act_regs_data_2_13_sva,
      act_regs_data_3_13_sva, act_config_in_InstFetch_mux_tmp[1:0]);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      = MUX_v_20_4_2(act_regs_data_0_12_sva, act_regs_data_1_12_sva, act_regs_data_2_12_sva,
      act_regs_data_3_12_sva, act_config_in_InstFetch_mux_tmp[1:0]);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      = MUX_v_20_4_2(act_regs_data_0_11_sva, act_regs_data_1_11_sva, act_regs_data_2_11_sva,
      act_regs_data_3_11_sva, act_config_in_InstFetch_mux_tmp[1:0]);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      = MUX_v_20_4_2(act_regs_data_0_10_sva, act_regs_data_1_10_sva, act_regs_data_2_10_sva,
      act_regs_data_3_10_sva, act_config_in_InstFetch_mux_tmp[1:0]);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      = MUX_v_20_4_2(act_regs_data_0_9_sva, act_regs_data_1_9_sva, act_regs_data_2_9_sva,
      act_regs_data_3_9_sva, act_config_in_InstFetch_mux_tmp[1:0]);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      = MUX_v_20_4_2(act_regs_data_0_8_sva, act_regs_data_1_8_sva, act_regs_data_2_8_sva,
      act_regs_data_3_8_sva, act_config_in_InstFetch_mux_tmp[1:0]);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      = MUX_v_20_4_2(act_regs_data_0_7_sva, act_regs_data_1_7_sva, act_regs_data_2_7_sva,
      act_regs_data_3_7_sva, act_config_in_InstFetch_mux_tmp[1:0]);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      = MUX_v_20_4_2(act_regs_data_0_6_sva, act_regs_data_1_6_sva, act_regs_data_2_6_sva,
      act_regs_data_3_6_sva, act_config_in_InstFetch_mux_tmp[1:0]);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      = MUX_v_20_4_2(act_regs_data_0_5_sva, act_regs_data_1_5_sva, act_regs_data_2_5_sva,
      act_regs_data_3_5_sva, act_config_in_InstFetch_mux_tmp[1:0]);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      = MUX_v_20_4_2(act_regs_data_0_4_sva, act_regs_data_1_4_sva, act_regs_data_2_4_sva,
      act_regs_data_3_4_sva, act_config_in_InstFetch_mux_tmp[1:0]);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      = MUX_v_20_4_2(act_regs_data_0_3_sva, act_regs_data_1_3_sva, act_regs_data_2_3_sva,
      act_regs_data_3_3_sva, act_config_in_InstFetch_mux_tmp[1:0]);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      = MUX_v_20_4_2(act_regs_data_0_2_sva, act_regs_data_1_2_sva, act_regs_data_2_2_sva,
      act_regs_data_3_2_sva, act_config_in_InstFetch_mux_tmp[1:0]);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      = MUX_v_20_4_2(act_regs_data_0_1_sva, act_regs_data_1_1_sva, act_regs_data_2_1_sva,
      act_regs_data_3_1_sva, act_config_in_InstFetch_mux_tmp[1:0]);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1
      = MUX_v_20_4_2(act_regs_data_0_0_sva, act_regs_data_1_0_sva, act_regs_data_2_0_sva,
      act_regs_data_3_0_sva, act_config_in_InstFetch_mux_tmp[1:0]);
  assign nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm
      = MUX_v_20_4_2(act_regs_data_0_15_sva, act_regs_data_1_15_sva, act_regs_data_2_15_sva,
      act_regs_data_3_15_sva, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm
      = MUX_v_20_4_2(act_regs_data_0_14_sva, act_regs_data_1_14_sva, act_regs_data_2_14_sva,
      act_regs_data_3_14_sva, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm
      = MUX_v_20_4_2(act_regs_data_0_13_sva, act_regs_data_1_13_sva, act_regs_data_2_13_sva,
      act_regs_data_3_13_sva, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_nv_scvector_cctor_nv_scvector_5_for_mux_1_itm
      = MUX_v_20_4_2(act_regs_data_0_12_sva, act_regs_data_1_12_sva, act_regs_data_2_12_sva,
      act_regs_data_3_12_sva, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      = MUX_v_20_4_2(act_regs_data_0_11_sva, act_regs_data_1_11_sva, act_regs_data_2_11_sva,
      act_regs_data_3_11_sva, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      = MUX_v_20_4_2(act_regs_data_0_10_sva, act_regs_data_1_10_sva, act_regs_data_2_10_sva,
      act_regs_data_3_10_sva, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      = MUX_v_20_4_2(act_regs_data_0_9_sva, act_regs_data_1_9_sva, act_regs_data_2_9_sva,
      act_regs_data_3_9_sva, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      = MUX_v_20_4_2(act_regs_data_0_8_sva, act_regs_data_1_8_sva, act_regs_data_2_8_sva,
      act_regs_data_3_8_sva, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      = MUX_v_20_4_2(act_regs_data_0_7_sva, act_regs_data_1_7_sva, act_regs_data_2_7_sva,
      act_regs_data_3_7_sva, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      = MUX_v_20_4_2(act_regs_data_0_6_sva, act_regs_data_1_6_sva, act_regs_data_2_6_sva,
      act_regs_data_3_6_sva, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      = MUX_v_20_4_2(act_regs_data_0_5_sva, act_regs_data_1_5_sva, act_regs_data_2_5_sva,
      act_regs_data_3_5_sva, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      = MUX_v_20_4_2(act_regs_data_0_4_sva, act_regs_data_1_4_sva, act_regs_data_2_4_sva,
      act_regs_data_3_4_sva, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      = MUX_v_20_4_2(act_regs_data_0_3_sva, act_regs_data_1_3_sva, act_regs_data_2_3_sva,
      act_regs_data_3_3_sva, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      = MUX_v_20_4_2(act_regs_data_0_2_sva, act_regs_data_1_2_sva, act_regs_data_2_2_sva,
      act_regs_data_3_2_sva, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      = MUX_v_20_4_2(act_regs_data_0_1_sva, act_regs_data_1_1_sva, act_regs_data_2_1_sva,
      act_regs_data_3_1_sva, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      = MUX_v_20_4_2(act_regs_data_0_0_sva, act_regs_data_1_0_sva, act_regs_data_2_0_sva,
      act_regs_data_3_0_sva, act_config_in_InstFetch_mux_tmp[3:2]);
  assign act_config_ActConfigRead_else_unequal_tmp_1 = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:0]==8'b00000010));
  assign act_config_ActConfigRead_unequal_tmp_1 = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:0]==8'b00000001));
  assign ActUnit_DecodeAxiRead_unequal_tmp_1 = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:8]==4'b1000));
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_21_nl = act_read_addrs_lpi_1_dfm_9
      & ({{4{ActUnit_DecodeAxiRead_unequal_tmp_1}}, ActUnit_DecodeAxiRead_unequal_tmp_1})
      & (signext_5_1(~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)) & ({{4{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign while_mux_124_ssc_mx0 = MUX_v_5_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_21_nl,
      act_read_addrs_lpi_1_dfm_5, is_start_sva);
  assign ActUnit_DecodeAxiWrite_else_not_17_nl = ~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0;
  assign act_read_addrs_lpi_1_dfm_9 = MUX_v_5_2_2(5'b00000, (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4:0]),
      ActUnit_DecodeAxiWrite_else_not_17_nl);
  assign ActUnit_DecodeAxiRead_and_cse_1 = act_config_ActConfigRead_unequal_tmp_1
      & (~ ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign act_config_InstIncr_if_if_unequal_tmp = act_config_output_counter_sva !=
      (operator_8_false_acc_tmp[7:0]);
  assign act_config_InstIncr_if_act_config_InstIncr_if_if_act_config_InstIncr_if_if_nor_mdf_sva_1
      = ~(act_config_InstIncr_if_if_unequal_tmp | (operator_8_false_acc_tmp[8]));
  assign nl_operator_8_false_acc_tmp = conv_u2s_8_9(act_config_num_output_sva) +
      9'b111111111;
  assign operator_8_false_acc_tmp = nl_operator_8_false_acc_tmp[8:0];
  assign act_config_InstIncr_if_equal_1_tmp = act_config_inst_counter_sva == (operator_6_false_acc_tmp[4:0]);
  assign act_config_InstIncr_act_config_InstIncr_if_and_svs_1 = act_config_InstIncr_if_equal_1_tmp
      & (operator_6_false_acc_tmp[6:5]==2'b00);
  assign nl_operator_6_false_acc_tmp = conv_u2s_6_7(act_config_num_inst_sva) + 7'b1111111;
  assign operator_6_false_acc_tmp = nl_operator_6_false_acc_tmp[6:0];
  assign ActUnit_RunInst_switch_lp_nor_ssc_sva_1 = ~((act_config_in_InstFetch_return_sva_4_2[1:0]!=2'b00));
  assign ActUnit_RunInst_switch_lp_and_ssc_sva_1 = (act_config_in_InstFetch_return_sva_4_2[1:0]==2'b11);
  assign ActUnit_RunInst_switch_lp_and_ssc_2_sva_1 = (act_config_in_InstFetch_return_sva_4_2[1:0]==2'b01);
  assign ActUnit_RunInst_switch_lp_and_ssc_1_sva_1 = (act_config_in_InstFetch_return_sva_4_2[1:0]==2'b10);
  assign ActUnit_RunInst_switch_lp_and_66_tmp_1 = (act_config_in_InstFetch_return_sva_4_2[1:0]==2'b11)
      & act_port_PopNB_mioi_return_rsc_z_mxwt;
  assign ActUnit_RunInst_switch_lp_and_50_tmp_1 = (act_config_in_InstFetch_return_sva_4_2[1:0]==2'b10)
      & act_port_PopNB_mioi_return_rsc_z_mxwt;
  assign ActUnit_RunInst_switch_lp_and_34_tmp_1 = (act_config_in_InstFetch_return_sva_4_2[1:0]==2'b01)
      & act_port_PopNB_mioi_return_rsc_z_mxwt;
  assign ActUnit_RunInst_switch_lp_and_18_tmp_1 = ActUnit_RunInst_switch_lp_nor_ssc_sva_1
      & act_port_PopNB_mioi_return_rsc_z_mxwt;
  assign ActUnit_RunInst_switch_lp_equal_tmp_20 = (act_config_in_InstFetch_return_sva_4_2[2])
      & ActUnit_RunInst_switch_lp_nor_7_itm;
  assign act_regs_data_0_15_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_0_15_sva,
      (act_port_PopNB_mioi_data_data_rsc_z_mxwt[319:300]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[319:300]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[319:300]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[319:300]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[319:300]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[319:300]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[319:300]),
      {while_asn_1344 , while_asn_1346 , while_asn_1348 , while_asn_1350 , while_asn_1352
      , while_asn_1354 , while_asn_1356 , while_asn_1358 , while_asn_1360});
  assign act_regs_data_1_15_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_1_15_sva,
      (act_port_PopNB_mioi_data_data_rsc_z_mxwt[319:300]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[319:300]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[319:300]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[319:300]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[319:300]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[319:300]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[319:300]),
      {while_asn_1326 , while_asn_1328 , while_asn_1330 , while_asn_1332 , while_asn_1334
      , while_asn_1336 , while_asn_1338 , while_asn_1340 , while_asn_1342});
  assign act_regs_data_2_15_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_2_15_sva,
      (act_port_PopNB_mioi_data_data_rsc_z_mxwt[319:300]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[319:300]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[319:300]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[319:300]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[319:300]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[319:300]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[319:300]),
      {while_asn_1308 , while_asn_1310 , while_asn_1312 , while_asn_1314 , while_asn_1316
      , while_asn_1318 , while_asn_1320 , while_asn_1322 , while_asn_1324});
  assign act_regs_data_3_15_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_3_15_sva,
      (act_port_PopNB_mioi_data_data_rsc_z_mxwt[319:300]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[319:300]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[319:300]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[319:300]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[319:300]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[319:300]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[319:300]),
      {while_asn_1290 , while_asn_1292 , while_asn_1294 , while_asn_1296 , while_asn_1298
      , while_asn_1300 , while_asn_1302 , while_asn_1304 , while_asn_1306});
  assign nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_1_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[3:2]),
      (act_config_inst_regs_16_sva_dfm_6[3:2]), not_tmp_34);
  assign nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_4_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[11:10]),
      (act_config_inst_regs_17_sva_dfm_6[3:2]), not_tmp_34);
  assign nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_7_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[19:18]),
      (act_config_inst_regs_18_sva_dfm_6[3:2]), not_tmp_34);
  assign nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_9_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[27:26]),
      (act_config_inst_regs_19_sva_dfm_6[3:2]), not_tmp_34);
  assign act_config_ActConfigWrite_if_mux_3_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[35:34]),
      (act_config_inst_regs_20_sva_dfm_6[3:2]), not_tmp_34);
  assign nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_11_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[43:42]),
      (act_config_inst_regs_21_sva_dfm_6[3:2]), not_tmp_34);
  assign nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_13_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[51:50]),
      (act_config_inst_regs_22_sva_dfm_6[3:2]), not_tmp_34);
  assign nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_15_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[59:58]),
      (act_config_inst_regs_23_sva_dfm_6[3:2]), not_tmp_34);
  assign act_config_ActConfigWrite_if_mux_5_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[67:66]),
      (act_config_inst_regs_24_sva_dfm_6[3:2]), not_tmp_34);
  assign nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_17_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[75:74]),
      (act_config_inst_regs_25_sva_dfm_6[3:2]), not_tmp_34);
  assign nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_19_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[83:82]),
      (act_config_inst_regs_26_sva_dfm_6[3:2]), not_tmp_34);
  assign nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_21_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[91:90]),
      (act_config_inst_regs_27_sva_dfm_6[3:2]), not_tmp_34);
  assign nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_23_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[99:98]),
      (act_config_inst_regs_28_sva_dfm_6[3:2]), not_tmp_34);
  assign nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_25_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[107:106]),
      (act_config_inst_regs_29_sva_dfm_6[3:2]), not_tmp_34);
  assign nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_27_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[115:114]),
      (act_config_inst_regs_30_sva_dfm_6[3:2]), not_tmp_34);
  assign nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_29_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[123:122]),
      (act_config_inst_regs_31_sva_dfm_6[3:2]), not_tmp_34);
  assign nvhls_get_slc_2U_NVUINT8_return_3_sva_1 = MUX_v_2_32_2((act_config_inst_regs_0_sva_dfm_5[3:2]),
      (act_config_inst_regs_1_sva_dfm_5[3:2]), (act_config_inst_regs_2_sva_dfm_5[3:2]),
      (act_config_inst_regs_3_sva_dfm_5[3:2]), (act_config_inst_regs_4_sva_dfm_5[3:2]),
      (act_config_inst_regs_5_sva_dfm_5[3:2]), (act_config_inst_regs_6_sva_dfm_5[3:2]),
      (act_config_inst_regs_7_sva_dfm_5[3:2]), (act_config_inst_regs_8_sva_dfm_5[3:2]),
      (act_config_inst_regs_9_sva_dfm_5[3:2]), (act_config_inst_regs_10_sva_dfm_5[3:2]),
      (act_config_inst_regs_11_sva_dfm_5[3:2]), (act_config_inst_regs_12_sva_dfm_5[3:2]),
      (act_config_inst_regs_13_sva_dfm_5[3:2]), (act_config_inst_regs_14_sva_dfm_5[3:2]),
      (act_config_inst_regs_15_sva_dfm_5[3:2]), nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_1_nl,
      nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_4_nl, nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_7_nl,
      nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_9_nl, act_config_ActConfigWrite_if_mux_3_nl,
      nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_11_nl, nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_13_nl,
      nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_15_nl, act_config_ActConfigWrite_if_mux_5_nl,
      nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_17_nl, nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_19_nl,
      nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_21_nl, nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_23_nl,
      nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_25_nl, nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_27_nl,
      nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_29_nl, act_config_inst_counter_sva);
  assign act_regs_data_0_14_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_0_14_sva,
      (act_port_PopNB_mioi_data_data_rsc_z_mxwt[299:280]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[299:280]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[299:280]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[299:280]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[299:280]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[299:280]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[299:280]),
      {while_asn_1344 , while_asn_1346 , while_asn_1348 , while_asn_1350 , while_asn_1352
      , while_asn_1354 , while_asn_1356 , while_asn_1358 , while_asn_1360});
  assign act_regs_data_1_14_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_1_14_sva,
      (act_port_PopNB_mioi_data_data_rsc_z_mxwt[299:280]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[299:280]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[299:280]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[299:280]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[299:280]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[299:280]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[299:280]),
      {while_asn_1326 , while_asn_1328 , while_asn_1330 , while_asn_1332 , while_asn_1334
      , while_asn_1336 , while_asn_1338 , while_asn_1340 , while_asn_1342});
  assign act_regs_data_2_14_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_2_14_sva,
      (act_port_PopNB_mioi_data_data_rsc_z_mxwt[299:280]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[299:280]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[299:280]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[299:280]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[299:280]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[299:280]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[299:280]),
      {while_asn_1308 , while_asn_1310 , while_asn_1312 , while_asn_1314 , while_asn_1316
      , while_asn_1318 , while_asn_1320 , while_asn_1322 , while_asn_1324});
  assign act_regs_data_3_14_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_3_14_sva,
      (act_port_PopNB_mioi_data_data_rsc_z_mxwt[299:280]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[299:280]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[299:280]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[299:280]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[299:280]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[299:280]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[299:280]),
      {while_asn_1290 , while_asn_1292 , while_asn_1294 , while_asn_1296 , while_asn_1298
      , while_asn_1300 , while_asn_1302 , while_asn_1304 , while_asn_1306});
  assign act_regs_data_0_13_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_0_13_sva,
      (act_port_PopNB_mioi_data_data_rsc_z_mxwt[279:260]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[279:260]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[279:260]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[279:260]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[279:260]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[279:260]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[279:260]),
      {while_asn_1344 , while_asn_1346 , while_asn_1348 , while_asn_1350 , while_asn_1352
      , while_asn_1354 , while_asn_1356 , while_asn_1358 , while_asn_1360});
  assign act_regs_data_1_13_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_1_13_sva,
      (act_port_PopNB_mioi_data_data_rsc_z_mxwt[279:260]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[279:260]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[279:260]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[279:260]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[279:260]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[279:260]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[279:260]),
      {while_asn_1326 , while_asn_1328 , while_asn_1330 , while_asn_1332 , while_asn_1334
      , while_asn_1336 , while_asn_1338 , while_asn_1340 , while_asn_1342});
  assign act_regs_data_2_13_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_2_13_sva,
      (act_port_PopNB_mioi_data_data_rsc_z_mxwt[279:260]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[279:260]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[279:260]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[279:260]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[279:260]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[279:260]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[279:260]),
      {while_asn_1308 , while_asn_1310 , while_asn_1312 , while_asn_1314 , while_asn_1316
      , while_asn_1318 , while_asn_1320 , while_asn_1322 , while_asn_1324});
  assign act_regs_data_3_13_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_3_13_sva,
      (act_port_PopNB_mioi_data_data_rsc_z_mxwt[279:260]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[279:260]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[279:260]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[279:260]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[279:260]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[279:260]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[279:260]),
      {while_asn_1290 , while_asn_1292 , while_asn_1294 , while_asn_1296 , while_asn_1298
      , while_asn_1300 , while_asn_1302 , while_asn_1304 , while_asn_1306});
  assign act_regs_data_0_12_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_0_12_sva,
      (act_port_PopNB_mioi_data_data_rsc_z_mxwt[259:240]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[259:240]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[259:240]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[259:240]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[259:240]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[259:240]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[259:240]),
      {while_asn_1344 , while_asn_1346 , while_asn_1348 , while_asn_1350 , while_asn_1352
      , while_asn_1354 , while_asn_1356 , while_asn_1358 , while_asn_1360});
  assign act_regs_data_1_12_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_1_12_sva,
      (act_port_PopNB_mioi_data_data_rsc_z_mxwt[259:240]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[259:240]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[259:240]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[259:240]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[259:240]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[259:240]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[259:240]),
      {while_asn_1326 , while_asn_1328 , while_asn_1330 , while_asn_1332 , while_asn_1334
      , while_asn_1336 , while_asn_1338 , while_asn_1340 , while_asn_1342});
  assign act_regs_data_2_12_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_2_12_sva,
      (act_port_PopNB_mioi_data_data_rsc_z_mxwt[259:240]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[259:240]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[259:240]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[259:240]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[259:240]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[259:240]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[259:240]),
      {while_asn_1308 , while_asn_1310 , while_asn_1312 , while_asn_1314 , while_asn_1316
      , while_asn_1318 , while_asn_1320 , while_asn_1322 , while_asn_1324});
  assign act_regs_data_3_12_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_3_12_sva,
      (act_port_PopNB_mioi_data_data_rsc_z_mxwt[259:240]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[259:240]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[259:240]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[259:240]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[259:240]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[259:240]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[259:240]),
      {while_asn_1290 , while_asn_1292 , while_asn_1294 , while_asn_1296 , while_asn_1298
      , while_asn_1300 , while_asn_1302 , while_asn_1304 , while_asn_1306});
  assign act_regs_data_0_11_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_0_11_sva,
      (act_port_PopNB_mioi_data_data_rsc_z_mxwt[239:220]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[239:220]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[239:220]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[239:220]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[239:220]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[239:220]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[239:220]),
      {while_asn_1344 , while_asn_1346 , while_asn_1348 , while_asn_1350 , while_asn_1352
      , while_asn_1354 , while_asn_1356 , while_asn_1358 , while_asn_1360});
  assign act_regs_data_1_11_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_1_11_sva,
      (act_port_PopNB_mioi_data_data_rsc_z_mxwt[239:220]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[239:220]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[239:220]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[239:220]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[239:220]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[239:220]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[239:220]),
      {while_asn_1326 , while_asn_1328 , while_asn_1330 , while_asn_1332 , while_asn_1334
      , while_asn_1336 , while_asn_1338 , while_asn_1340 , while_asn_1342});
  assign act_regs_data_2_11_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_2_11_sva,
      (act_port_PopNB_mioi_data_data_rsc_z_mxwt[239:220]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[239:220]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[239:220]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[239:220]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[239:220]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[239:220]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[239:220]),
      {while_asn_1308 , while_asn_1310 , while_asn_1312 , while_asn_1314 , while_asn_1316
      , while_asn_1318 , while_asn_1320 , while_asn_1322 , while_asn_1324});
  assign act_regs_data_3_11_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_3_11_sva,
      (act_port_PopNB_mioi_data_data_rsc_z_mxwt[239:220]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[239:220]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[239:220]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[239:220]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[239:220]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[239:220]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[239:220]),
      {while_asn_1290 , while_asn_1292 , while_asn_1294 , while_asn_1296 , while_asn_1298
      , while_asn_1300 , while_asn_1302 , while_asn_1304 , while_asn_1306});
  assign act_regs_data_0_10_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_0_10_sva,
      (act_port_PopNB_mioi_data_data_rsc_z_mxwt[219:200]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[219:200]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[219:200]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[219:200]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[219:200]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[219:200]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[219:200]),
      {while_asn_1344 , while_asn_1346 , while_asn_1348 , while_asn_1350 , while_asn_1352
      , while_asn_1354 , while_asn_1356 , while_asn_1358 , while_asn_1360});
  assign act_regs_data_1_10_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_1_10_sva,
      (act_port_PopNB_mioi_data_data_rsc_z_mxwt[219:200]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[219:200]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[219:200]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[219:200]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[219:200]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[219:200]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[219:200]),
      {while_asn_1326 , while_asn_1328 , while_asn_1330 , while_asn_1332 , while_asn_1334
      , while_asn_1336 , while_asn_1338 , while_asn_1340 , while_asn_1342});
  assign act_regs_data_2_10_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_2_10_sva,
      (act_port_PopNB_mioi_data_data_rsc_z_mxwt[219:200]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[219:200]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[219:200]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[219:200]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[219:200]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[219:200]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[219:200]),
      {while_asn_1308 , while_asn_1310 , while_asn_1312 , while_asn_1314 , while_asn_1316
      , while_asn_1318 , while_asn_1320 , while_asn_1322 , while_asn_1324});
  assign act_regs_data_3_10_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_3_10_sva,
      (act_port_PopNB_mioi_data_data_rsc_z_mxwt[219:200]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[219:200]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[219:200]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[219:200]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[219:200]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[219:200]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[219:200]),
      {while_asn_1290 , while_asn_1292 , while_asn_1294 , while_asn_1296 , while_asn_1298
      , while_asn_1300 , while_asn_1302 , while_asn_1304 , while_asn_1306});
  assign act_regs_data_0_9_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_0_9_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[199:180]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[199:180]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[199:180]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[199:180]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[199:180]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[199:180]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[199:180]),
      {while_asn_1344 , while_asn_1346 , while_asn_1348 , while_asn_1350 , while_asn_1352
      , while_asn_1354 , while_asn_1356 , while_asn_1358 , while_asn_1360});
  assign act_regs_data_1_9_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_1_9_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[199:180]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[199:180]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[199:180]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[199:180]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[199:180]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[199:180]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[199:180]),
      {while_asn_1326 , while_asn_1328 , while_asn_1330 , while_asn_1332 , while_asn_1334
      , while_asn_1336 , while_asn_1338 , while_asn_1340 , while_asn_1342});
  assign act_regs_data_2_9_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_2_9_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[199:180]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[199:180]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[199:180]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[199:180]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[199:180]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[199:180]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[199:180]),
      {while_asn_1308 , while_asn_1310 , while_asn_1312 , while_asn_1314 , while_asn_1316
      , while_asn_1318 , while_asn_1320 , while_asn_1322 , while_asn_1324});
  assign act_regs_data_3_9_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_3_9_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[199:180]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[199:180]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[199:180]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[199:180]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[199:180]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[199:180]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[199:180]),
      {while_asn_1290 , while_asn_1292 , while_asn_1294 , while_asn_1296 , while_asn_1298
      , while_asn_1300 , while_asn_1302 , while_asn_1304 , while_asn_1306});
  assign act_regs_data_0_8_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_0_8_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[179:160]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[179:160]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[179:160]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[179:160]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[179:160]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[179:160]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[179:160]),
      {while_asn_1344 , while_asn_1346 , while_asn_1348 , while_asn_1350 , while_asn_1352
      , while_asn_1354 , while_asn_1356 , while_asn_1358 , while_asn_1360});
  assign act_regs_data_1_8_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_1_8_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[179:160]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[179:160]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[179:160]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[179:160]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[179:160]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[179:160]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[179:160]),
      {while_asn_1326 , while_asn_1328 , while_asn_1330 , while_asn_1332 , while_asn_1334
      , while_asn_1336 , while_asn_1338 , while_asn_1340 , while_asn_1342});
  assign act_regs_data_2_8_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_2_8_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[179:160]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[179:160]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[179:160]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[179:160]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[179:160]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[179:160]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[179:160]),
      {while_asn_1308 , while_asn_1310 , while_asn_1312 , while_asn_1314 , while_asn_1316
      , while_asn_1318 , while_asn_1320 , while_asn_1322 , while_asn_1324});
  assign act_regs_data_3_8_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_3_8_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[179:160]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[179:160]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[179:160]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[179:160]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[179:160]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[179:160]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[179:160]),
      {while_asn_1290 , while_asn_1292 , while_asn_1294 , while_asn_1296 , while_asn_1298
      , while_asn_1300 , while_asn_1302 , while_asn_1304 , while_asn_1306});
  assign act_regs_data_0_7_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_0_7_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[159:140]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[159:140]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[159:140]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[159:140]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[159:140]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[159:140]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[159:140]),
      {while_asn_1344 , while_asn_1346 , while_asn_1348 , while_asn_1350 , while_asn_1352
      , while_asn_1354 , while_asn_1356 , while_asn_1358 , while_asn_1360});
  assign act_regs_data_1_7_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_1_7_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[159:140]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[159:140]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[159:140]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[159:140]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[159:140]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[159:140]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[159:140]),
      {while_asn_1326 , while_asn_1328 , while_asn_1330 , while_asn_1332 , while_asn_1334
      , while_asn_1336 , while_asn_1338 , while_asn_1340 , while_asn_1342});
  assign act_regs_data_2_7_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_2_7_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[159:140]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[159:140]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[159:140]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[159:140]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[159:140]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[159:140]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[159:140]),
      {while_asn_1308 , while_asn_1310 , while_asn_1312 , while_asn_1314 , while_asn_1316
      , while_asn_1318 , while_asn_1320 , while_asn_1322 , while_asn_1324});
  assign act_regs_data_3_7_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_3_7_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[159:140]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[159:140]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[159:140]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[159:140]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[159:140]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[159:140]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[159:140]),
      {while_asn_1290 , while_asn_1292 , while_asn_1294 , while_asn_1296 , while_asn_1298
      , while_asn_1300 , while_asn_1302 , while_asn_1304 , while_asn_1306});
  assign act_regs_data_0_6_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_0_6_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[139:120]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[139:120]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[139:120]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[139:120]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[139:120]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[139:120]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[139:120]),
      {while_asn_1344 , while_asn_1346 , while_asn_1348 , while_asn_1350 , while_asn_1352
      , while_asn_1354 , while_asn_1356 , while_asn_1358 , while_asn_1360});
  assign act_regs_data_1_6_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_1_6_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[139:120]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[139:120]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[139:120]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[139:120]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[139:120]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[139:120]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[139:120]),
      {while_asn_1326 , while_asn_1328 , while_asn_1330 , while_asn_1332 , while_asn_1334
      , while_asn_1336 , while_asn_1338 , while_asn_1340 , while_asn_1342});
  assign act_regs_data_2_6_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_2_6_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[139:120]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[139:120]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[139:120]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[139:120]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[139:120]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[139:120]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[139:120]),
      {while_asn_1308 , while_asn_1310 , while_asn_1312 , while_asn_1314 , while_asn_1316
      , while_asn_1318 , while_asn_1320 , while_asn_1322 , while_asn_1324});
  assign act_regs_data_3_6_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_3_6_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[139:120]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[139:120]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[139:120]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[139:120]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[139:120]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[139:120]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[139:120]),
      {while_asn_1290 , while_asn_1292 , while_asn_1294 , while_asn_1296 , while_asn_1298
      , while_asn_1300 , while_asn_1302 , while_asn_1304 , while_asn_1306});
  assign act_regs_data_0_5_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_0_5_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[119:100]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[119:100]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[119:100]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[119:100]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[119:100]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[119:100]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[119:100]),
      {while_asn_1344 , while_asn_1346 , while_asn_1348 , while_asn_1350 , while_asn_1352
      , while_asn_1354 , while_asn_1356 , while_asn_1358 , while_asn_1360});
  assign act_regs_data_1_5_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_1_5_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[119:100]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[119:100]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[119:100]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[119:100]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[119:100]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[119:100]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[119:100]),
      {while_asn_1326 , while_asn_1328 , while_asn_1330 , while_asn_1332 , while_asn_1334
      , while_asn_1336 , while_asn_1338 , while_asn_1340 , while_asn_1342});
  assign act_regs_data_2_5_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_2_5_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[119:100]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[119:100]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[119:100]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[119:100]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[119:100]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[119:100]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[119:100]),
      {while_asn_1308 , while_asn_1310 , while_asn_1312 , while_asn_1314 , while_asn_1316
      , while_asn_1318 , while_asn_1320 , while_asn_1322 , while_asn_1324});
  assign act_regs_data_3_5_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_3_5_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[119:100]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[119:100]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[119:100]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[119:100]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[119:100]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[119:100]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[119:100]),
      {while_asn_1290 , while_asn_1292 , while_asn_1294 , while_asn_1296 , while_asn_1298
      , while_asn_1300 , while_asn_1302 , while_asn_1304 , while_asn_1306});
  assign act_regs_data_0_4_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_0_4_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[99:80]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[99:80]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[99:80]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[99:80]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[99:80]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[99:80]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[99:80]),
      {while_asn_1344 , while_asn_1346 , while_asn_1348 , while_asn_1350 , while_asn_1352
      , while_asn_1354 , while_asn_1356 , while_asn_1358 , while_asn_1360});
  assign act_regs_data_1_4_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_1_4_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[99:80]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[99:80]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[99:80]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[99:80]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[99:80]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[99:80]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[99:80]),
      {while_asn_1326 , while_asn_1328 , while_asn_1330 , while_asn_1332 , while_asn_1334
      , while_asn_1336 , while_asn_1338 , while_asn_1340 , while_asn_1342});
  assign act_regs_data_2_4_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_2_4_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[99:80]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[99:80]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[99:80]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[99:80]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[99:80]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[99:80]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[99:80]),
      {while_asn_1308 , while_asn_1310 , while_asn_1312 , while_asn_1314 , while_asn_1316
      , while_asn_1318 , while_asn_1320 , while_asn_1322 , while_asn_1324});
  assign act_regs_data_3_4_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_3_4_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[99:80]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[99:80]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[99:80]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[99:80]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[99:80]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[99:80]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[99:80]),
      {while_asn_1290 , while_asn_1292 , while_asn_1294 , while_asn_1296 , while_asn_1298
      , while_asn_1300 , while_asn_1302 , while_asn_1304 , while_asn_1306});
  assign act_regs_data_0_3_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_0_3_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[79:60]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[79:60]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[79:60]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[79:60]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[79:60]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[79:60]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[79:60]),
      {while_asn_1344 , while_asn_1346 , while_asn_1348 , while_asn_1350 , while_asn_1352
      , while_asn_1354 , while_asn_1356 , while_asn_1358 , while_asn_1360});
  assign act_regs_data_1_3_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_1_3_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[79:60]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[79:60]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[79:60]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[79:60]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[79:60]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[79:60]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[79:60]),
      {while_asn_1326 , while_asn_1328 , while_asn_1330 , while_asn_1332 , while_asn_1334
      , while_asn_1336 , while_asn_1338 , while_asn_1340 , while_asn_1342});
  assign act_regs_data_2_3_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_2_3_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[79:60]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[79:60]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[79:60]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[79:60]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[79:60]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[79:60]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[79:60]),
      {while_asn_1308 , while_asn_1310 , while_asn_1312 , while_asn_1314 , while_asn_1316
      , while_asn_1318 , while_asn_1320 , while_asn_1322 , while_asn_1324});
  assign act_regs_data_3_3_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_3_3_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[79:60]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[79:60]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[79:60]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[79:60]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[79:60]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[79:60]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[79:60]),
      {while_asn_1290 , while_asn_1292 , while_asn_1294 , while_asn_1296 , while_asn_1298
      , while_asn_1300 , while_asn_1302 , while_asn_1304 , while_asn_1306});
  assign act_regs_data_0_2_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_0_2_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[59:40]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[59:40]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[59:40]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[59:40]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[59:40]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[59:40]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[59:40]),
      {while_asn_1344 , while_asn_1346 , while_asn_1348 , while_asn_1350 , while_asn_1352
      , while_asn_1354 , while_asn_1356 , while_asn_1358 , while_asn_1360});
  assign act_regs_data_1_2_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_1_2_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[59:40]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[59:40]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[59:40]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[59:40]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[59:40]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[59:40]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[59:40]),
      {while_asn_1326 , while_asn_1328 , while_asn_1330 , while_asn_1332 , while_asn_1334
      , while_asn_1336 , while_asn_1338 , while_asn_1340 , while_asn_1342});
  assign act_regs_data_2_2_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_2_2_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[59:40]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[59:40]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[59:40]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[59:40]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[59:40]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[59:40]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[59:40]),
      {while_asn_1308 , while_asn_1310 , while_asn_1312 , while_asn_1314 , while_asn_1316
      , while_asn_1318 , while_asn_1320 , while_asn_1322 , while_asn_1324});
  assign act_regs_data_3_2_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_3_2_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[59:40]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[59:40]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[59:40]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[59:40]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[59:40]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[59:40]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[59:40]),
      {while_asn_1290 , while_asn_1292 , while_asn_1294 , while_asn_1296 , while_asn_1298
      , while_asn_1300 , while_asn_1302 , while_asn_1304 , while_asn_1306});
  assign act_regs_data_0_1_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_0_1_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[39:20]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[39:20]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[39:20]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[39:20]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[39:20]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[39:20]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[39:20]),
      {while_asn_1344 , while_asn_1346 , while_asn_1348 , while_asn_1350 , while_asn_1352
      , while_asn_1354 , while_asn_1356 , while_asn_1358 , while_asn_1360});
  assign act_regs_data_1_1_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_1_1_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[39:20]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[39:20]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[39:20]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[39:20]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[39:20]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[39:20]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[39:20]),
      {while_asn_1326 , while_asn_1328 , while_asn_1330 , while_asn_1332 , while_asn_1334
      , while_asn_1336 , while_asn_1338 , while_asn_1340 , while_asn_1342});
  assign act_regs_data_2_1_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_2_1_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[39:20]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[39:20]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[39:20]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[39:20]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[39:20]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[39:20]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[39:20]),
      {while_asn_1308 , while_asn_1310 , while_asn_1312 , while_asn_1314 , while_asn_1316
      , while_asn_1318 , while_asn_1320 , while_asn_1322 , while_asn_1324});
  assign act_regs_data_3_1_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_3_1_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[39:20]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[39:20]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[39:20]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[39:20]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[39:20]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[39:20]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[39:20]),
      {while_asn_1290 , while_asn_1292 , while_asn_1294 , while_asn_1296 , while_asn_1298
      , while_asn_1300 , while_asn_1302 , while_asn_1304 , while_asn_1306});
  assign act_regs_data_0_0_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_0_0_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[19:0]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[19:0]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[19:0]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[19:0]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[19:0]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[19:0]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[19:0]),
      {while_asn_1344 , while_asn_1346 , while_asn_1348 , while_asn_1350 , while_asn_1352
      , while_asn_1354 , while_asn_1356 , while_asn_1358 , while_asn_1360});
  assign act_regs_data_1_0_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_1_0_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[19:0]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[19:0]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[19:0]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[19:0]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[19:0]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[19:0]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[19:0]),
      {while_asn_1326 , while_asn_1328 , while_asn_1330 , while_asn_1332 , while_asn_1334
      , while_asn_1336 , while_asn_1338 , while_asn_1340 , while_asn_1342});
  assign act_regs_data_2_0_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_2_0_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[19:0]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[19:0]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[19:0]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[19:0]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[19:0]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[19:0]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[19:0]),
      {while_asn_1308 , while_asn_1310 , while_asn_1312 , while_asn_1314 , while_asn_1316
      , while_asn_1318 , while_asn_1320 , while_asn_1322 , while_asn_1324});
  assign act_regs_data_3_0_sva_dfm_3 = MUX1HOT_v_20_9_2(act_regs_data_3_0_sva, (act_port_PopNB_mioi_data_data_rsc_z_mxwt[19:0]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva,
      (ActUnit_RunInst_case_8_EAdd_act_regs_data_sva[19:0]), (ActUnit_RunInst_case_9_EMul_act_regs_data_sva[19:0]),
      (ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva[19:0]), (ActUnit_RunInst_case_11_Tanh_act_regs_data_sva[19:0]),
      (ActUnit_RunInst_case_12_Relu_act_regs_data_sva[19:0]), (ActUnit_RunInst_case_13_OneX_act_regs_data_sva[19:0]),
      {while_asn_1290 , while_asn_1292 , while_asn_1294 , while_asn_1296 , while_asn_1298
      , while_asn_1300 , while_asn_1302 , while_asn_1304 , while_asn_1306});
  assign act_config_ActConfigWrite_mux_34_nl = MUX_s_1_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[8]),
      act_config_is_zero_first_sva, act_config_ActConfigRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiWrite_mux_37_nl = MUX_s_1_2_2(act_config_ActConfigWrite_mux_34_nl,
      act_config_is_zero_first_sva, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxi_if_mux_83_nl = MUX_s_1_2_2(act_config_is_zero_first_sva,
      ActUnit_DecodeAxiWrite_mux_37_nl, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign ActUnit_DecodeAxi_mux_89_nl = MUX_s_1_2_2(act_config_is_zero_first_sva,
      ActUnit_DecodeAxi_if_mux_83_nl, rva_in_PopNB_mioi_return_rsc_z_mxwt);
  assign act_config_is_zero_first_sva_dfm_4_mx0 = MUX_s_1_2_2(ActUnit_DecodeAxi_mux_89_nl,
      act_config_is_zero_first_sva, is_start_sva);
  assign is_incr_lpi_1_dfm_2 = act_port_PopNB_mioi_return_rsc_z_mxwt | (~ ActUnit_RunInst_switch_lp_equal_tmp_2)
      | (~ is_start_sva);
  assign ActUnit_RunLoad_if_else_nor_ssc_sva_1 = ~((nvhls_get_slc_2U_NVUINT8_return_3_sva_1!=2'b00));
  assign ActUnit_RunLoad_if_else_and_ssc_2_sva_1 = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b01);
  assign ActUnit_RunLoad_if_else_and_ssc_1_sva_1 = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b10);
  assign ActUnit_RunLoad_if_else_and_ssc_sva_1 = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b11);
  assign ActUnit_PushOutput_and_tmp_1 = ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_cse
      & (~ ActUnit_RunInst_switch_lp_equal_tmp_3);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_22_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[7:0])
      & (signext_8_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{7{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{7{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_0_lpi_1_dfm_5_mx0 = MUX_v_8_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_22_nl,
      act_write_data_data_0_0_lpi_1_dfm_4, is_start_sva);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_23_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[15:8])
      & (signext_8_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{7{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{7{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_1_lpi_1_dfm_5_mx0 = MUX_v_8_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_23_nl,
      act_write_data_data_0_1_lpi_1_dfm_4, is_start_sva);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_24_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[23:16])
      & (signext_8_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{7{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{7{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_2_lpi_1_dfm_5_mx0 = MUX_v_8_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_24_nl,
      act_write_data_data_0_2_lpi_1_dfm_4, is_start_sva);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_25_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[31:24])
      & (signext_8_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{7{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{7{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_3_lpi_1_dfm_5_mx0 = MUX_v_8_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_25_nl,
      act_write_data_data_0_3_lpi_1_dfm_4, is_start_sva);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_26_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[39:32])
      & (signext_8_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{7{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{7{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_4_lpi_1_dfm_5_mx0 = MUX_v_8_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_26_nl,
      act_write_data_data_0_4_lpi_1_dfm_4, is_start_sva);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_27_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[47:40])
      & (signext_8_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{7{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{7{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_5_lpi_1_dfm_5_mx0 = MUX_v_8_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_27_nl,
      act_write_data_data_0_5_lpi_1_dfm_4, is_start_sva);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_28_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[55:48])
      & (signext_8_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{7{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{7{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_6_lpi_1_dfm_5_mx0 = MUX_v_8_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_28_nl,
      act_write_data_data_0_6_lpi_1_dfm_4, is_start_sva);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_29_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[63:56])
      & (signext_8_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{7{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{7{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_7_lpi_1_dfm_5_mx0 = MUX_v_8_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_29_nl,
      act_write_data_data_0_7_lpi_1_dfm_4, is_start_sva);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_30_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[71:64])
      & (signext_8_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{7{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{7{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_8_lpi_1_dfm_5_mx0 = MUX_v_8_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_30_nl,
      act_write_data_data_0_8_lpi_1_dfm_4, is_start_sva);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_31_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[79:72])
      & (signext_8_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{7{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{7{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_9_lpi_1_dfm_5_mx0 = MUX_v_8_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_31_nl,
      act_write_data_data_0_9_lpi_1_dfm_4, is_start_sva);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_32_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[87:80])
      & (signext_8_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{7{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{7{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_10_lpi_1_dfm_5_mx0 = MUX_v_8_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_32_nl,
      act_write_data_data_0_10_lpi_1_dfm_4, is_start_sva);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_33_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[95:88])
      & (signext_8_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{7{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{7{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_11_lpi_1_dfm_5_mx0 = MUX_v_8_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_33_nl,
      act_write_data_data_0_11_lpi_1_dfm_4, is_start_sva);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_34_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[103:96])
      & (signext_8_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{7{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{7{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_12_lpi_1_dfm_5_mx0 = MUX_v_8_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_34_nl,
      act_write_data_data_0_12_lpi_1_dfm_4, is_start_sva);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_35_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[111:104])
      & (signext_8_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{7{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{7{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_13_lpi_1_dfm_5_mx0 = MUX_v_8_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_35_nl,
      act_write_data_data_0_13_lpi_1_dfm_4, is_start_sva);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_36_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[119:112])
      & (signext_8_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{7{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{7{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_14_lpi_1_dfm_5_mx0 = MUX_v_8_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_36_nl,
      act_write_data_data_0_14_lpi_1_dfm_4, is_start_sva);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_37_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[127:120])
      & (signext_8_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{7{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{7{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_15_lpi_1_dfm_5_mx0 = MUX_v_8_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_37_nl,
      act_write_data_data_0_15_lpi_1_dfm_4, is_start_sva);
  assign act_config_ActConfigRead_else_else_not_22 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:0]==8'b00000011);
  assign while_asn_1290 = ~(is_start_sva & (~(ActUnit_RunInst_switch_lp_equal_tmp_20
      | ActUnit_RunInst_switch_lp_equal_tmp_1 | ActUnit_RunInst_switch_lp_equal_tmp_3
      | ActUnit_RunInst_switch_lp_nor_tmp | ((~ ActUnit_RunInst_switch_lp_and_ssc_sva_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_4) | ((~ ActUnit_RunInst_switch_lp_and_ssc_sva_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_5) | ((~ ActUnit_RunInst_switch_lp_and_ssc_sva_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_6) | ((~ ActUnit_RunInst_switch_lp_and_ssc_sva_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_7) | ((~ ActUnit_RunInst_switch_lp_and_ssc_sva_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_8) | ((~ ActUnit_RunInst_switch_lp_and_ssc_sva_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_9) | ((~ ActUnit_RunInst_switch_lp_and_ssc_sva_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_10) | ((~ ActUnit_RunInst_switch_lp_and_66_tmp_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_2))));
  assign while_asn_1292 = ActUnit_RunInst_switch_lp_and_66_tmp_1 & ActUnit_RunInst_switch_lp_equal_tmp_2
      & is_start_sva;
  assign while_asn_1294 = ActUnit_RunInst_switch_lp_and_ssc_sva_1 & ActUnit_RunInst_switch_lp_equal_tmp_4
      & is_start_sva;
  assign while_asn_1296 = ActUnit_RunInst_switch_lp_and_ssc_sva_1 & ActUnit_RunInst_switch_lp_equal_tmp_5
      & is_start_sva;
  assign while_asn_1298 = ActUnit_RunInst_switch_lp_and_ssc_sva_1 & ActUnit_RunInst_switch_lp_equal_tmp_6
      & is_start_sva;
  assign while_asn_1300 = ActUnit_RunInst_switch_lp_and_ssc_sva_1 & ActUnit_RunInst_switch_lp_equal_tmp_7
      & is_start_sva;
  assign while_asn_1302 = ActUnit_RunInst_switch_lp_and_ssc_sva_1 & ActUnit_RunInst_switch_lp_equal_tmp_8
      & is_start_sva;
  assign while_asn_1304 = ActUnit_RunInst_switch_lp_and_ssc_sva_1 & ActUnit_RunInst_switch_lp_equal_tmp_9
      & is_start_sva;
  assign while_asn_1306 = ActUnit_RunInst_switch_lp_and_ssc_sva_1 & ActUnit_RunInst_switch_lp_equal_tmp_10
      & is_start_sva;
  assign while_asn_1308 = ~(is_start_sva & (~(ActUnit_RunInst_switch_lp_equal_tmp_20
      | ActUnit_RunInst_switch_lp_equal_tmp_1 | ActUnit_RunInst_switch_lp_equal_tmp_3
      | ActUnit_RunInst_switch_lp_nor_tmp | ((~ ActUnit_RunInst_switch_lp_and_ssc_1_sva_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_4) | ((~ ActUnit_RunInst_switch_lp_and_ssc_1_sva_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_5) | ((~ ActUnit_RunInst_switch_lp_and_ssc_1_sva_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_6) | ((~ ActUnit_RunInst_switch_lp_and_ssc_1_sva_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_7) | ((~ ActUnit_RunInst_switch_lp_and_ssc_1_sva_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_8) | ((~ ActUnit_RunInst_switch_lp_and_ssc_1_sva_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_9) | ((~ ActUnit_RunInst_switch_lp_and_ssc_1_sva_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_10) | ((~ ActUnit_RunInst_switch_lp_and_50_tmp_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_2))));
  assign while_asn_1310 = ActUnit_RunInst_switch_lp_and_50_tmp_1 & ActUnit_RunInst_switch_lp_equal_tmp_2
      & is_start_sva;
  assign while_asn_1312 = ActUnit_RunInst_switch_lp_and_ssc_1_sva_1 & ActUnit_RunInst_switch_lp_equal_tmp_4
      & is_start_sva;
  assign while_asn_1314 = ActUnit_RunInst_switch_lp_and_ssc_1_sva_1 & ActUnit_RunInst_switch_lp_equal_tmp_5
      & is_start_sva;
  assign while_asn_1316 = ActUnit_RunInst_switch_lp_and_ssc_1_sva_1 & ActUnit_RunInst_switch_lp_equal_tmp_6
      & is_start_sva;
  assign while_asn_1318 = ActUnit_RunInst_switch_lp_and_ssc_1_sva_1 & ActUnit_RunInst_switch_lp_equal_tmp_7
      & is_start_sva;
  assign while_asn_1320 = ActUnit_RunInst_switch_lp_and_ssc_1_sva_1 & ActUnit_RunInst_switch_lp_equal_tmp_8
      & is_start_sva;
  assign while_asn_1322 = ActUnit_RunInst_switch_lp_and_ssc_1_sva_1 & ActUnit_RunInst_switch_lp_equal_tmp_9
      & is_start_sva;
  assign while_asn_1324 = ActUnit_RunInst_switch_lp_and_ssc_1_sva_1 & ActUnit_RunInst_switch_lp_equal_tmp_10
      & is_start_sva;
  assign while_asn_1326 = ~(is_start_sva & (~(ActUnit_RunInst_switch_lp_equal_tmp_20
      | ActUnit_RunInst_switch_lp_equal_tmp_1 | ActUnit_RunInst_switch_lp_equal_tmp_3
      | ActUnit_RunInst_switch_lp_nor_tmp | ((~ ActUnit_RunInst_switch_lp_and_ssc_2_sva_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_4) | ((~ ActUnit_RunInst_switch_lp_and_ssc_2_sva_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_5) | ((~ ActUnit_RunInst_switch_lp_and_ssc_2_sva_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_6) | ((~ ActUnit_RunInst_switch_lp_and_ssc_2_sva_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_7) | ((~ ActUnit_RunInst_switch_lp_and_ssc_2_sva_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_8) | ((~ ActUnit_RunInst_switch_lp_and_ssc_2_sva_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_9) | ((~ ActUnit_RunInst_switch_lp_and_ssc_2_sva_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_10) | ((~ ActUnit_RunInst_switch_lp_and_34_tmp_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_2))));
  assign while_asn_1328 = ActUnit_RunInst_switch_lp_and_34_tmp_1 & ActUnit_RunInst_switch_lp_equal_tmp_2
      & is_start_sva;
  assign while_asn_1330 = ActUnit_RunInst_switch_lp_and_ssc_2_sva_1 & ActUnit_RunInst_switch_lp_equal_tmp_4
      & is_start_sva;
  assign while_asn_1332 = ActUnit_RunInst_switch_lp_and_ssc_2_sva_1 & ActUnit_RunInst_switch_lp_equal_tmp_5
      & is_start_sva;
  assign while_asn_1334 = ActUnit_RunInst_switch_lp_and_ssc_2_sva_1 & ActUnit_RunInst_switch_lp_equal_tmp_6
      & is_start_sva;
  assign while_asn_1336 = ActUnit_RunInst_switch_lp_and_ssc_2_sva_1 & ActUnit_RunInst_switch_lp_equal_tmp_7
      & is_start_sva;
  assign while_asn_1338 = ActUnit_RunInst_switch_lp_and_ssc_2_sva_1 & ActUnit_RunInst_switch_lp_equal_tmp_8
      & is_start_sva;
  assign while_asn_1340 = ActUnit_RunInst_switch_lp_and_ssc_2_sva_1 & ActUnit_RunInst_switch_lp_equal_tmp_9
      & is_start_sva;
  assign while_asn_1342 = ActUnit_RunInst_switch_lp_and_ssc_2_sva_1 & ActUnit_RunInst_switch_lp_equal_tmp_10
      & is_start_sva;
  assign while_asn_1344 = ~(is_start_sva & (~(ActUnit_RunInst_switch_lp_equal_tmp_20
      | ActUnit_RunInst_switch_lp_equal_tmp_1 | ActUnit_RunInst_switch_lp_equal_tmp_3
      | ActUnit_RunInst_switch_lp_nor_tmp | ((~ ActUnit_RunInst_switch_lp_nor_ssc_sva_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_4) | ((~ ActUnit_RunInst_switch_lp_nor_ssc_sva_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_5) | ((~ ActUnit_RunInst_switch_lp_nor_ssc_sva_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_6) | ((~ ActUnit_RunInst_switch_lp_nor_ssc_sva_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_7) | ((~ ActUnit_RunInst_switch_lp_nor_ssc_sva_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_8) | ((~ ActUnit_RunInst_switch_lp_nor_ssc_sva_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_9) | ((~ ActUnit_RunInst_switch_lp_nor_ssc_sva_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_10) | ((~ ActUnit_RunInst_switch_lp_and_18_tmp_1)
      & ActUnit_RunInst_switch_lp_equal_tmp_2))));
  assign while_asn_1346 = ActUnit_RunInst_switch_lp_and_18_tmp_1 & ActUnit_RunInst_switch_lp_equal_tmp_2
      & is_start_sva;
  assign while_asn_1348 = ActUnit_RunInst_switch_lp_nor_ssc_sva_1 & ActUnit_RunInst_switch_lp_equal_tmp_4
      & is_start_sva;
  assign while_asn_1350 = ActUnit_RunInst_switch_lp_nor_ssc_sva_1 & ActUnit_RunInst_switch_lp_equal_tmp_5
      & is_start_sva;
  assign while_asn_1352 = ActUnit_RunInst_switch_lp_nor_ssc_sva_1 & ActUnit_RunInst_switch_lp_equal_tmp_6
      & is_start_sva;
  assign while_asn_1354 = ActUnit_RunInst_switch_lp_nor_ssc_sva_1 & ActUnit_RunInst_switch_lp_equal_tmp_7
      & is_start_sva;
  assign while_asn_1356 = ActUnit_RunInst_switch_lp_nor_ssc_sva_1 & ActUnit_RunInst_switch_lp_equal_tmp_8
      & is_start_sva;
  assign while_asn_1358 = ActUnit_RunInst_switch_lp_nor_ssc_sva_1 & ActUnit_RunInst_switch_lp_equal_tmp_9
      & is_start_sva;
  assign while_asn_1360 = ActUnit_RunInst_switch_lp_nor_ssc_sva_1 & ActUnit_RunInst_switch_lp_equal_tmp_10
      & is_start_sva;
  assign while_asn_1364 = act_config_is_zero_first_sva_dfm_4_mx0 & ActUnit_PushOutput_and_tmp_1
      & is_start_sva;
  assign while_asn_1366 = ActUnit_RunLoad_if_else_and_ssc_sva_1 & (~ act_config_is_zero_first_sva_dfm_4_mx0)
      & ActUnit_PushOutput_and_tmp_1 & is_start_sva;
  assign while_asn_1370 = ActUnit_RunLoad_if_else_and_ssc_1_sva_1 & (~ act_config_is_zero_first_sva_dfm_4_mx0)
      & ActUnit_PushOutput_and_tmp_1 & is_start_sva;
  assign while_asn_1374 = ActUnit_RunLoad_if_else_and_ssc_2_sva_1 & (~ act_config_is_zero_first_sva_dfm_4_mx0)
      & ActUnit_PushOutput_and_tmp_1 & is_start_sva;
  assign while_asn_1378 = ActUnit_RunLoad_if_else_nor_ssc_sva_1 & (~ act_config_is_zero_first_sva_dfm_4_mx0)
      & ActUnit_PushOutput_and_tmp_1 & is_start_sva;
  assign ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_1_tmp
      = ~(act_config_is_zero_first_sva | ActUnit_RunInst_switch_lp_equal_tmp_1 |
      ActUnit_RunInst_switch_lp_equal_tmp_2 | ActUnit_RunInst_switch_lp_equal_tmp_3
      | ActUnit_RunInst_switch_lp_equal_tmp_4 | ActUnit_RunInst_switch_lp_equal_tmp_5
      | ActUnit_RunInst_switch_lp_equal_tmp_6 | ActUnit_RunInst_switch_lp_equal_tmp_7
      | ActUnit_RunInst_switch_lp_equal_tmp_8 | ActUnit_RunInst_switch_lp_equal_tmp_9
      | ActUnit_RunInst_switch_lp_equal_tmp_10 | ActUnit_RunInst_switch_lp_nor_tmp);
  assign ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_and_1_nl
      = MUX_v_5_2_2(5'b00000, act_write_addrs_lpi_1_dfm_5, ActUnit_RunInst_switch_lp_equal_tmp_1);
  assign while_mux_125_tmp = MUX_v_5_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_3_mx0w2,
      ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_and_1_nl,
      is_start_sva);
  assign mux_nl = MUX_s_1_2_2(ActUnit_CheckStart_if_ActUnit_CheckStart_if_and_1_cse,
      ActUnit_RunInst_switch_lp_equal_tmp_1, is_start_sva);
  assign mux_tmp_1 = MUX_s_1_2_2(is_start_sva, mux_nl, ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_cse);
  assign and_dcpl = (act_config_in_InstFetch_mux_tmp[6]) & (act_config_in_InstFetch_mux_tmp[4]);
  assign and_dcpl_1 = (act_config_in_InstFetch_mux_tmp[5]) & (~ (act_config_in_InstFetch_mux_tmp[7]));
  assign and_dcpl_5 = (~ (act_config_in_InstFetch_mux_tmp[5])) & (act_config_in_InstFetch_mux_tmp[7]);
  assign and_dcpl_8 = (~ (act_config_in_InstFetch_mux_tmp[6])) & (act_config_in_InstFetch_mux_tmp[4]);
  assign and_dcpl_11 = (act_config_in_InstFetch_mux_tmp[5]) & (act_config_in_InstFetch_mux_tmp[7]);
  assign or_16_cse = act_port_PopNB_mioi_return_rsc_z_mxwt | (~ ActUnit_RunInst_switch_lp_equal_tmp_2);
  assign nor_14_nl = ~((~ rva_in_PopNB_mioi_return_rsc_z_mxwt) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:8]!=4'b1001));
  assign mux_5_cse = MUX_s_1_2_2(nor_14_nl, ActUnit_RunInst_switch_lp_equal_tmp_1,
      is_start_sva);
  assign or_dcpl_8 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:10]!=2'b10);
  assign or_dcpl_9 = or_dcpl_8 | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9:8]!=2'b01);
  assign and_dcpl_31 = (~ (operator_6_false_acc_tmp[6])) & act_config_InstIncr_if_equal_1_tmp;
  assign nor_tmp_6 = is_start_sva & ActUnit_RunInst_switch_lp_equal_tmp_1;
  assign or_64_nl = (~ is_start_sva) | ActUnit_RunInst_switch_lp_equal_tmp_1;
  assign mux_15_nl = MUX_s_1_2_2(nor_tmp_6, or_64_nl, ActUnit_CheckStart_if_ActUnit_CheckStart_if_and_1_cse);
  assign mux_tmp_16 = MUX_s_1_2_2(is_start_sva, mux_15_nl, ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_cse);
  assign or_dcpl_13 = ~(rva_in_PopNB_mioi_return_rsc_z_mxwt & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign or_dcpl_15 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9:8]!=2'b00) | or_dcpl_13;
  assign or_dcpl_22 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:2]!=6'b000000) |
      or_dcpl_8;
  assign not_tmp_34 = ~((ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_23_4_mx1_tmp_7_0==8'b00000011)
      & act_config_ActConfigRead_else_unequal_tmp_1 & act_config_ActConfigRead_unequal_tmp_1
      & (~ ActUnit_DecodeAxiRead_unequal_tmp_1) & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & rva_in_PopNB_mioi_return_rsc_z_mxwt & (~ is_start_sva));
  assign or_dcpl_27 = or_dcpl_22 | or_dcpl_15 | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | is_start_sva | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]);
  assign and_dcpl_45 = (~ act_port_PopNB_mioi_return_rsc_z_mxwt) & ActUnit_RunInst_switch_lp_equal_tmp_2;
  assign or_dcpl_33 = (while_mux_125_tmp[1:0]!=2'b00);
  assign or_dcpl_34 = (while_mux_125_tmp[4:3]!=2'b00);
  assign or_dcpl_35 = or_dcpl_34 | (while_mux_125_tmp[2]);
  assign or_dcpl_38 = (while_mux_125_tmp[1:0]!=2'b01);
  assign or_dcpl_41 = (while_mux_125_tmp[1:0]!=2'b10);
  assign or_dcpl_44 = ~((while_mux_125_tmp[1:0]==2'b11));
  assign or_dcpl_47 = or_dcpl_34 | (~ (while_mux_125_tmp[2]));
  assign or_dcpl_56 = (while_mux_125_tmp[4:3]!=2'b01);
  assign or_dcpl_57 = or_dcpl_56 | (while_mux_125_tmp[2]);
  assign or_dcpl_66 = or_dcpl_56 | (~ (while_mux_125_tmp[2]));
  assign or_dcpl_75 = (while_mux_125_tmp[4:3]!=2'b10);
  assign or_dcpl_76 = or_dcpl_75 | (while_mux_125_tmp[2]);
  assign or_dcpl_85 = or_dcpl_75 | (~ (while_mux_125_tmp[2]));
  assign or_dcpl_94 = ~((while_mux_125_tmp[4:3]==2'b11));
  assign or_dcpl_95 = or_dcpl_94 | (while_mux_125_tmp[2]);
  assign or_dcpl_104 = or_dcpl_94 | (~ (while_mux_125_tmp[2]));
  assign or_dcpl_116 = or_dcpl_13 | is_start_sva;
  assign and_dcpl_65 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:0]==8'b00000010);
  assign or_tmp_61 = (~ is_start_sva) & (fsm_output[2]);
  assign and_158_cse = (~ mux_tmp_16) & (fsm_output[1]);
  assign act_config_is_valid_sva_mx0c0 = (~ ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_cse)
      & (fsm_output[1]);
  assign act_config_output_counter_sva_mx0c1 = or_16_cse & and_dcpl_31 & (~ (operator_6_false_acc_tmp[5]))
      & is_start_sva & (fsm_output[2]);
  assign is_start_sva_mx0c1 = (~ is_start_sva) & ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_cse
      & (fsm_output[1]);
  assign act_write_addrs_lpi_1_dfm_5_mx0c2 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:8]==4'b1001)
      & rva_in_PopNB_mioi_return_rsc_z_mxwt & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (~ is_start_sva) & (fsm_output[2]);
  assign or_dcpl = (while_asn_1364 & (~ ActUnit_RunLoad_if_else_nor_ssc_sva_1)) |
      (~(is_start_sva & ActUnit_PushOutput_and_tmp_1 & (ActUnit_RunLoad_if_else_nor_ssc_sva_1
      | act_config_is_zero_first_sva_dfm_4_mx0)));
  assign or_dcpl_122 = (while_asn_1364 & (~ ActUnit_RunLoad_if_else_and_ssc_2_sva_1))
      | (~(is_start_sva & ActUnit_PushOutput_and_tmp_1 & (ActUnit_RunLoad_if_else_and_ssc_2_sva_1
      | act_config_is_zero_first_sva_dfm_4_mx0)));
  assign or_dcpl_123 = (while_asn_1364 & (~ ActUnit_RunLoad_if_else_and_ssc_1_sva_1))
      | (~(is_start_sva & ActUnit_PushOutput_and_tmp_1 & (ActUnit_RunLoad_if_else_and_ssc_1_sva_1
      | act_config_is_zero_first_sva_dfm_4_mx0)));
  assign or_dcpl_124 = (while_asn_1364 & (~ ActUnit_RunLoad_if_else_and_ssc_sva_1))
      | (~(is_start_sva & ActUnit_PushOutput_and_tmp_1 & (ActUnit_RunLoad_if_else_and_ssc_sva_1
      | act_config_is_zero_first_sva_dfm_4_mx0)));
  assign and_tmp = (and_dcpl_45 | (~ is_start_sva)) & or_884_itm;
  assign and_dcpl_73 = (((~ act_config_ActConfigRead_else_else_not_22) & ActUnit_DecodeAxiRead_and_9_cse)
      | ActUnit_DecodeAxiRead_unequal_tmp_1) & or_dcpl_9;
  assign and_1551_tmp = (((~ act_config_ActConfigRead_else_else_not_22) & ActUnit_DecodeAxiRead_and_cse_1
      & (~ and_dcpl_65)) | ActUnit_DecodeAxiRead_unequal_tmp_1) & or_dcpl_9;
  assign ActUnit_PushAxiRsp_if_and_cse = (~ ActUnit_DecodeAxiRead_and_cse_1) & or_dcpl_9
      & (~ and_dcpl_73);
  assign ActUnit_PushAxiRsp_if_and_1_cse = ActUnit_DecodeAxiRead_and_9_cse & (~ and_dcpl_73);
  assign or_tmp_756 = ((operator_6_false_acc_tmp[6]) | (~ act_config_InstIncr_if_equal_1_tmp)
      | (operator_6_false_acc_tmp[5])) & (fsm_output[2]);
  assign mux_118_nl = MUX_s_1_2_2(or_958_cse, or_957_cse, act_config_inst_counter_sva[0]);
  assign mux_117_nl = MUX_s_1_2_2(or_956_cse, or_955_cse, act_config_inst_counter_sva[0]);
  assign mux_119_nl = MUX_s_1_2_2(mux_118_nl, mux_117_nl, act_config_inst_counter_sva[1]);
  assign mux_115_nl = MUX_s_1_2_2(or_954_cse, or_953_cse, act_config_inst_counter_sva[0]);
  assign mux_114_nl = MUX_s_1_2_2(or_952_cse, or_951_cse, act_config_inst_counter_sva[0]);
  assign mux_116_nl = MUX_s_1_2_2(mux_115_nl, mux_114_nl, act_config_inst_counter_sva[1]);
  assign mux_120_nl = MUX_s_1_2_2(mux_119_nl, mux_116_nl, act_config_inst_counter_sva[2]);
  assign mux_111_nl = MUX_s_1_2_2(or_950_cse, or_949_cse, act_config_inst_counter_sva[0]);
  assign mux_110_nl = MUX_s_1_2_2(or_948_cse, or_947_cse, act_config_inst_counter_sva[0]);
  assign mux_112_nl = MUX_s_1_2_2(mux_111_nl, mux_110_nl, act_config_inst_counter_sva[1]);
  assign mux_108_nl = MUX_s_1_2_2(or_946_cse, or_945_cse, act_config_inst_counter_sva[0]);
  assign mux_107_nl = MUX_s_1_2_2(or_944_cse, or_943_cse, act_config_inst_counter_sva[0]);
  assign mux_109_nl = MUX_s_1_2_2(mux_108_nl, mux_107_nl, act_config_inst_counter_sva[1]);
  assign mux_113_nl = MUX_s_1_2_2(mux_112_nl, mux_109_nl, act_config_inst_counter_sva[2]);
  assign mux_121_nl = MUX_s_1_2_2(mux_120_nl, mux_113_nl, act_config_inst_counter_sva[3]);
  assign mux_103_nl = MUX_s_1_2_2(or_942_cse, or_941_cse, act_config_inst_counter_sva[0]);
  assign mux_102_nl = MUX_s_1_2_2(or_940_cse, or_939_cse, act_config_inst_counter_sva[0]);
  assign mux_104_nl = MUX_s_1_2_2(mux_103_nl, mux_102_nl, act_config_inst_counter_sva[1]);
  assign mux_100_nl = MUX_s_1_2_2(or_938_cse, or_937_cse, act_config_inst_counter_sva[0]);
  assign mux_99_nl = MUX_s_1_2_2(or_936_cse, or_935_cse, act_config_inst_counter_sva[0]);
  assign mux_101_nl = MUX_s_1_2_2(mux_100_nl, mux_99_nl, act_config_inst_counter_sva[1]);
  assign mux_105_nl = MUX_s_1_2_2(mux_104_nl, mux_101_nl, act_config_inst_counter_sva[2]);
  assign mux_96_nl = MUX_s_1_2_2(or_934_cse, or_933_cse, act_config_inst_counter_sva[0]);
  assign mux_95_nl = MUX_s_1_2_2(or_932_cse, or_931_cse, act_config_inst_counter_sva[0]);
  assign mux_97_nl = MUX_s_1_2_2(mux_96_nl, mux_95_nl, act_config_inst_counter_sva[1]);
  assign mux_93_nl = MUX_s_1_2_2(or_930_cse, or_929_cse, act_config_inst_counter_sva[0]);
  assign mux_92_nl = MUX_s_1_2_2(or_928_cse, or_925_cse, act_config_inst_counter_sva[0]);
  assign mux_94_nl = MUX_s_1_2_2(mux_93_nl, mux_92_nl, act_config_inst_counter_sva[1]);
  assign mux_98_nl = MUX_s_1_2_2(mux_97_nl, mux_94_nl, act_config_inst_counter_sva[2]);
  assign mux_106_nl = MUX_s_1_2_2(mux_105_nl, mux_98_nl, act_config_inst_counter_sva[3]);
  assign mux_tmp_118 = MUX_s_1_2_2(mux_121_nl, mux_106_nl, act_config_inst_counter_sva[4]);
  assign not_tmp_67 = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11]) & (fsm_output[2]));
  assign or_tmp_791 = (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10:8]!=3'b001) | not_tmp_67;
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_done_Push_mioi_iswt0_cse <= 1'b0;
      reg_output_port_Push_mioi_iswt0_cse <= 1'b0;
      reg_start_PopNB_mioi_iswt0_cse <= 1'b0;
      reg_rva_out_Push_mioi_iswt0_cse <= 1'b0;
      reg_act_port_PopNB_mioi_iswt0_cse <= 1'b0;
      reg_rva_in_PopNB_mioi_iswt0_cse <= 1'b0;
      act_config_inst_counter_sva <= 5'b00000;
      act_config_inst_regs_16_sva_0 <= 1'b0;
      act_config_inst_regs_1_sva_0 <= 1'b0;
      act_config_inst_regs_17_sva_0 <= 1'b0;
      ActUnit_RunInst_switch_lp_equal_tmp_1 <= 1'b0;
      act_config_in_InstFetch_return_sva_4_2 <= 3'b000;
      ActUnit_RunInst_switch_lp_equal_tmp_2 <= 1'b0;
      ActUnit_RunInst_switch_lp_equal_tmp_3 <= 1'b0;
      ActUnit_RunInst_switch_lp_equal_tmp_4 <= 1'b0;
      ActUnit_RunInst_switch_lp_equal_tmp_5 <= 1'b0;
      ActUnit_RunInst_switch_lp_equal_tmp_6 <= 1'b0;
      ActUnit_RunInst_switch_lp_equal_tmp_7 <= 1'b0;
      ActUnit_RunInst_switch_lp_equal_tmp_8 <= 1'b0;
      ActUnit_RunInst_switch_lp_equal_tmp_9 <= 1'b0;
      ActUnit_RunInst_switch_lp_equal_tmp_10 <= 1'b0;
      ActUnit_RunInst_switch_lp_nor_tmp <= 1'b0;
      reg_ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_23_4_ftd_12
          <= 8'b00000000;
    end
    else if ( ActUnitRun_wen ) begin
      reg_done_Push_mioi_iswt0_cse <= done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct_mx0;
      reg_output_port_Push_mioi_iswt0_cse <= output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct_mx0;
      reg_start_PopNB_mioi_iswt0_cse <= or_tmp_61;
      reg_rva_out_Push_mioi_iswt0_cse <= rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct_mx0;
      reg_act_port_PopNB_mioi_iswt0_cse <= act_port_PopNB_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_psct_mx0;
      reg_rva_in_PopNB_mioi_iswt0_cse <= and_158_cse;
      act_config_inst_counter_sva <= MUX_v_5_2_2(and_1554_nl, act_config_inst_counter_sva,
          nand_6_nl);
      act_config_inst_regs_16_sva_0 <= MUX_s_1_2_2(act_config_inst_regs_16_sva_0,
          nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_2_nl, fsm_output[2]);
      act_config_inst_regs_1_sva_0 <= MUX_s_1_2_2(act_config_inst_regs_1_sva_0, nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_33_nl,
          fsm_output[2]);
      act_config_inst_regs_17_sva_0 <= MUX_s_1_2_2(act_config_inst_regs_17_sva_0,
          nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_5_nl, fsm_output[2]);
      ActUnit_RunInst_switch_lp_equal_tmp_1 <= MUX_s_1_2_2(ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0,
          while_else_1_while_else_1_nand_nl, fsm_output[2]);
      act_config_in_InstFetch_return_sva_4_2 <= act_config_in_InstFetch_mux_tmp[4:2];
      ActUnit_RunInst_switch_lp_equal_tmp_2 <= ActUnit_RunInst_switch_lp_equal_tmp_11;
      ActUnit_RunInst_switch_lp_equal_tmp_3 <= ActUnit_RunInst_switch_lp_equal_tmp_12;
      ActUnit_RunInst_switch_lp_equal_tmp_4 <= ActUnit_RunInst_switch_lp_equal_tmp_13;
      ActUnit_RunInst_switch_lp_equal_tmp_5 <= ActUnit_RunInst_switch_lp_equal_tmp_14;
      ActUnit_RunInst_switch_lp_equal_tmp_6 <= ActUnit_RunInst_switch_lp_equal_tmp_15;
      ActUnit_RunInst_switch_lp_equal_tmp_7 <= ActUnit_RunInst_switch_lp_equal_tmp_16;
      ActUnit_RunInst_switch_lp_equal_tmp_8 <= ActUnit_RunInst_switch_lp_equal_tmp_17;
      ActUnit_RunInst_switch_lp_equal_tmp_9 <= ActUnit_RunInst_switch_lp_equal_tmp_18;
      ActUnit_RunInst_switch_lp_equal_tmp_10 <= ActUnit_RunInst_switch_lp_equal_tmp_19;
      ActUnit_RunInst_switch_lp_nor_tmp <= ActUnit_RunInst_switch_lp_nor_tmp_1;
      reg_ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_23_4_ftd_12
          <= MUX_v_8_2_2(reg_ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_23_4_ftd_12,
          (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:0]), or_tmp_61);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_config_is_valid_sva <= 1'b0;
    end
    else if ( ActUnitRun_wen & (((~(act_config_ActConfigRead_unequal_tmp_1 | ActUnit_DecodeAxiRead_unequal_tmp_1))
        & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt & rva_in_PopNB_mioi_return_rsc_z_mxwt
        & (~((ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_cse & (fsm_output[1]))
        | (is_start_sva & (fsm_output[2])) | (fsm_output[0])))) | act_config_is_valid_sva_mx0c0)
        ) begin
      act_config_is_valid_sva <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[0]) & (~
          act_config_is_valid_sva_mx0c0);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_config_is_zero_first_sva <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((act_config_InstIncr_act_config_InstIncr_if_and_svs_1
        & is_incr_lpi_1_dfm_2 & (fsm_output[2])) | or_tmp_61) ) begin
      act_config_is_zero_first_sva <= MUX_s_1_2_2(act_config_InstIncr_if_act_config_InstIncr_if_and_1_nl,
          ActUnit_DecodeAxi_mux_88_nl, or_tmp_61);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_regs_data_0_15_sva <= 20'b00000000000000000000;
      act_regs_data_1_15_sva <= 20'b00000000000000000000;
      act_regs_data_2_15_sva <= 20'b00000000000000000000;
      act_regs_data_3_15_sva <= 20'b00000000000000000000;
      act_regs_data_0_14_sva <= 20'b00000000000000000000;
      act_regs_data_1_14_sva <= 20'b00000000000000000000;
      act_regs_data_2_14_sva <= 20'b00000000000000000000;
      act_regs_data_3_14_sva <= 20'b00000000000000000000;
      act_regs_data_0_13_sva <= 20'b00000000000000000000;
      act_regs_data_1_13_sva <= 20'b00000000000000000000;
      act_regs_data_2_13_sva <= 20'b00000000000000000000;
      act_regs_data_3_13_sva <= 20'b00000000000000000000;
      act_regs_data_0_12_sva <= 20'b00000000000000000000;
      act_regs_data_1_12_sva <= 20'b00000000000000000000;
      act_regs_data_2_12_sva <= 20'b00000000000000000000;
      act_regs_data_3_12_sva <= 20'b00000000000000000000;
      act_regs_data_0_11_sva <= 20'b00000000000000000000;
      act_regs_data_1_11_sva <= 20'b00000000000000000000;
      act_regs_data_2_11_sva <= 20'b00000000000000000000;
      act_regs_data_3_11_sva <= 20'b00000000000000000000;
      act_regs_data_0_10_sva <= 20'b00000000000000000000;
      act_regs_data_1_10_sva <= 20'b00000000000000000000;
      act_regs_data_2_10_sva <= 20'b00000000000000000000;
      act_regs_data_3_10_sva <= 20'b00000000000000000000;
      act_regs_data_0_9_sva <= 20'b00000000000000000000;
      act_regs_data_1_9_sva <= 20'b00000000000000000000;
      act_regs_data_2_9_sva <= 20'b00000000000000000000;
      act_regs_data_3_9_sva <= 20'b00000000000000000000;
      act_regs_data_0_8_sva <= 20'b00000000000000000000;
      act_regs_data_1_8_sva <= 20'b00000000000000000000;
      act_regs_data_2_8_sva <= 20'b00000000000000000000;
      act_regs_data_3_8_sva <= 20'b00000000000000000000;
      act_regs_data_0_7_sva <= 20'b00000000000000000000;
      act_regs_data_1_7_sva <= 20'b00000000000000000000;
      act_regs_data_2_7_sva <= 20'b00000000000000000000;
      act_regs_data_3_7_sva <= 20'b00000000000000000000;
      act_regs_data_0_6_sva <= 20'b00000000000000000000;
      act_regs_data_1_6_sva <= 20'b00000000000000000000;
      act_regs_data_2_6_sva <= 20'b00000000000000000000;
      act_regs_data_3_6_sva <= 20'b00000000000000000000;
      act_regs_data_0_5_sva <= 20'b00000000000000000000;
      act_regs_data_1_5_sva <= 20'b00000000000000000000;
      act_regs_data_2_5_sva <= 20'b00000000000000000000;
      act_regs_data_3_5_sva <= 20'b00000000000000000000;
      act_regs_data_0_4_sva <= 20'b00000000000000000000;
      act_regs_data_1_4_sva <= 20'b00000000000000000000;
      act_regs_data_2_4_sva <= 20'b00000000000000000000;
      act_regs_data_3_4_sva <= 20'b00000000000000000000;
      act_regs_data_0_3_sva <= 20'b00000000000000000000;
      act_regs_data_1_3_sva <= 20'b00000000000000000000;
      act_regs_data_2_3_sva <= 20'b00000000000000000000;
      act_regs_data_3_3_sva <= 20'b00000000000000000000;
      act_regs_data_0_2_sva <= 20'b00000000000000000000;
      act_regs_data_1_2_sva <= 20'b00000000000000000000;
      act_regs_data_2_2_sva <= 20'b00000000000000000000;
      act_regs_data_3_2_sva <= 20'b00000000000000000000;
      act_regs_data_0_1_sva <= 20'b00000000000000000000;
      act_regs_data_1_1_sva <= 20'b00000000000000000000;
      act_regs_data_2_1_sva <= 20'b00000000000000000000;
      act_regs_data_3_1_sva <= 20'b00000000000000000000;
      act_regs_data_0_0_sva <= 20'b00000000000000000000;
      act_regs_data_1_0_sva <= 20'b00000000000000000000;
      act_regs_data_2_0_sva <= 20'b00000000000000000000;
      act_regs_data_3_0_sva <= 20'b00000000000000000000;
    end
    else if ( act_regs_data_and_cse ) begin
      act_regs_data_0_15_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_nor_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[319:300]),
          act_regs_data_0_15_sva_dfm_3, {nor_18_cse , while_asn_1378 , or_dcpl});
      act_regs_data_1_15_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_2_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[319:300]),
          act_regs_data_1_15_sva_dfm_3, {nor_19_cse , while_asn_1374 , or_dcpl_122});
      act_regs_data_2_15_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_1_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[319:300]),
          act_regs_data_2_15_sva_dfm_3, {nor_20_cse , while_asn_1370 , or_dcpl_123});
      act_regs_data_3_15_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[319:300]),
          act_regs_data_3_15_sva_dfm_3, {nor_21_cse , while_asn_1366 , or_dcpl_124});
      act_regs_data_0_14_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_nor_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[299:280]),
          act_regs_data_0_14_sva_dfm_3, {nor_18_cse , while_asn_1378 , or_dcpl});
      act_regs_data_1_14_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_2_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[299:280]),
          act_regs_data_1_14_sva_dfm_3, {nor_19_cse , while_asn_1374 , or_dcpl_122});
      act_regs_data_2_14_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_1_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[299:280]),
          act_regs_data_2_14_sva_dfm_3, {nor_20_cse , while_asn_1370 , or_dcpl_123});
      act_regs_data_3_14_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[299:280]),
          act_regs_data_3_14_sva_dfm_3, {nor_21_cse , while_asn_1366 , or_dcpl_124});
      act_regs_data_0_13_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_nor_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[279:260]),
          act_regs_data_0_13_sva_dfm_3, {nor_18_cse , while_asn_1378 , or_dcpl});
      act_regs_data_1_13_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_2_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[279:260]),
          act_regs_data_1_13_sva_dfm_3, {nor_19_cse , while_asn_1374 , or_dcpl_122});
      act_regs_data_2_13_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_1_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[279:260]),
          act_regs_data_2_13_sva_dfm_3, {nor_20_cse , while_asn_1370 , or_dcpl_123});
      act_regs_data_3_13_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[279:260]),
          act_regs_data_3_13_sva_dfm_3, {nor_21_cse , while_asn_1366 , or_dcpl_124});
      act_regs_data_0_12_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_nor_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[259:240]),
          act_regs_data_0_12_sva_dfm_3, {nor_18_cse , while_asn_1378 , or_dcpl});
      act_regs_data_1_12_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_2_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[259:240]),
          act_regs_data_1_12_sva_dfm_3, {nor_19_cse , while_asn_1374 , or_dcpl_122});
      act_regs_data_2_12_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_1_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[259:240]),
          act_regs_data_2_12_sva_dfm_3, {nor_20_cse , while_asn_1370 , or_dcpl_123});
      act_regs_data_3_12_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[259:240]),
          act_regs_data_3_12_sva_dfm_3, {nor_21_cse , while_asn_1366 , or_dcpl_124});
      act_regs_data_0_11_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_nor_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[239:220]),
          act_regs_data_0_11_sva_dfm_3, {nor_18_cse , while_asn_1378 , or_dcpl});
      act_regs_data_1_11_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_2_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[239:220]),
          act_regs_data_1_11_sva_dfm_3, {nor_19_cse , while_asn_1374 , or_dcpl_122});
      act_regs_data_2_11_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_1_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[239:220]),
          act_regs_data_2_11_sva_dfm_3, {nor_20_cse , while_asn_1370 , or_dcpl_123});
      act_regs_data_3_11_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[239:220]),
          act_regs_data_3_11_sva_dfm_3, {nor_21_cse , while_asn_1366 , or_dcpl_124});
      act_regs_data_0_10_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_nor_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[219:200]),
          act_regs_data_0_10_sva_dfm_3, {nor_18_cse , while_asn_1378 , or_dcpl});
      act_regs_data_1_10_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_2_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[219:200]),
          act_regs_data_1_10_sva_dfm_3, {nor_19_cse , while_asn_1374 , or_dcpl_122});
      act_regs_data_2_10_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_1_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[219:200]),
          act_regs_data_2_10_sva_dfm_3, {nor_20_cse , while_asn_1370 , or_dcpl_123});
      act_regs_data_3_10_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[219:200]),
          act_regs_data_3_10_sva_dfm_3, {nor_21_cse , while_asn_1366 , or_dcpl_124});
      act_regs_data_0_9_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_nor_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[199:180]),
          act_regs_data_0_9_sva_dfm_3, {nor_18_cse , while_asn_1378 , or_dcpl});
      act_regs_data_1_9_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_2_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[199:180]),
          act_regs_data_1_9_sva_dfm_3, {nor_19_cse , while_asn_1374 , or_dcpl_122});
      act_regs_data_2_9_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_1_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[199:180]),
          act_regs_data_2_9_sva_dfm_3, {nor_20_cse , while_asn_1370 , or_dcpl_123});
      act_regs_data_3_9_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[199:180]),
          act_regs_data_3_9_sva_dfm_3, {nor_21_cse , while_asn_1366 , or_dcpl_124});
      act_regs_data_0_8_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_nor_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[179:160]),
          act_regs_data_0_8_sva_dfm_3, {nor_18_cse , while_asn_1378 , or_dcpl});
      act_regs_data_1_8_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_2_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[179:160]),
          act_regs_data_1_8_sva_dfm_3, {nor_19_cse , while_asn_1374 , or_dcpl_122});
      act_regs_data_2_8_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_1_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[179:160]),
          act_regs_data_2_8_sva_dfm_3, {nor_20_cse , while_asn_1370 , or_dcpl_123});
      act_regs_data_3_8_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[179:160]),
          act_regs_data_3_8_sva_dfm_3, {nor_21_cse , while_asn_1366 , or_dcpl_124});
      act_regs_data_0_7_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_nor_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[159:140]),
          act_regs_data_0_7_sva_dfm_3, {nor_18_cse , while_asn_1378 , or_dcpl});
      act_regs_data_1_7_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_2_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[159:140]),
          act_regs_data_1_7_sva_dfm_3, {nor_19_cse , while_asn_1374 , or_dcpl_122});
      act_regs_data_2_7_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_1_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[159:140]),
          act_regs_data_2_7_sva_dfm_3, {nor_20_cse , while_asn_1370 , or_dcpl_123});
      act_regs_data_3_7_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[159:140]),
          act_regs_data_3_7_sva_dfm_3, {nor_21_cse , while_asn_1366 , or_dcpl_124});
      act_regs_data_0_6_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_nor_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[139:120]),
          act_regs_data_0_6_sva_dfm_3, {nor_18_cse , while_asn_1378 , or_dcpl});
      act_regs_data_1_6_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_2_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[139:120]),
          act_regs_data_1_6_sva_dfm_3, {nor_19_cse , while_asn_1374 , or_dcpl_122});
      act_regs_data_2_6_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_1_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[139:120]),
          act_regs_data_2_6_sva_dfm_3, {nor_20_cse , while_asn_1370 , or_dcpl_123});
      act_regs_data_3_6_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[139:120]),
          act_regs_data_3_6_sva_dfm_3, {nor_21_cse , while_asn_1366 , or_dcpl_124});
      act_regs_data_0_5_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_nor_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[119:100]),
          act_regs_data_0_5_sva_dfm_3, {nor_18_cse , while_asn_1378 , or_dcpl});
      act_regs_data_1_5_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_2_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[119:100]),
          act_regs_data_1_5_sva_dfm_3, {nor_19_cse , while_asn_1374 , or_dcpl_122});
      act_regs_data_2_5_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_1_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[119:100]),
          act_regs_data_2_5_sva_dfm_3, {nor_20_cse , while_asn_1370 , or_dcpl_123});
      act_regs_data_3_5_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[119:100]),
          act_regs_data_3_5_sva_dfm_3, {nor_21_cse , while_asn_1366 , or_dcpl_124});
      act_regs_data_0_4_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_nor_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[99:80]),
          act_regs_data_0_4_sva_dfm_3, {nor_18_cse , while_asn_1378 , or_dcpl});
      act_regs_data_1_4_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_2_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[99:80]),
          act_regs_data_1_4_sva_dfm_3, {nor_19_cse , while_asn_1374 , or_dcpl_122});
      act_regs_data_2_4_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_1_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[99:80]),
          act_regs_data_2_4_sva_dfm_3, {nor_20_cse , while_asn_1370 , or_dcpl_123});
      act_regs_data_3_4_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[99:80]),
          act_regs_data_3_4_sva_dfm_3, {nor_21_cse , while_asn_1366 , or_dcpl_124});
      act_regs_data_0_3_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_nor_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[79:60]),
          act_regs_data_0_3_sva_dfm_3, {nor_18_cse , while_asn_1378 , or_dcpl});
      act_regs_data_1_3_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_2_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[79:60]),
          act_regs_data_1_3_sva_dfm_3, {nor_19_cse , while_asn_1374 , or_dcpl_122});
      act_regs_data_2_3_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_1_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[79:60]),
          act_regs_data_2_3_sva_dfm_3, {nor_20_cse , while_asn_1370 , or_dcpl_123});
      act_regs_data_3_3_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[79:60]),
          act_regs_data_3_3_sva_dfm_3, {nor_21_cse , while_asn_1366 , or_dcpl_124});
      act_regs_data_0_2_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_nor_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[59:40]),
          act_regs_data_0_2_sva_dfm_3, {nor_18_cse , while_asn_1378 , or_dcpl});
      act_regs_data_1_2_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_2_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[59:40]),
          act_regs_data_1_2_sva_dfm_3, {nor_19_cse , while_asn_1374 , or_dcpl_122});
      act_regs_data_2_2_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_1_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[59:40]),
          act_regs_data_2_2_sva_dfm_3, {nor_20_cse , while_asn_1370 , or_dcpl_123});
      act_regs_data_3_2_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[59:40]),
          act_regs_data_3_2_sva_dfm_3, {nor_21_cse , while_asn_1366 , or_dcpl_124});
      act_regs_data_0_1_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_nor_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[39:20]),
          act_regs_data_0_1_sva_dfm_3, {nor_18_cse , while_asn_1378 , or_dcpl});
      act_regs_data_1_1_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_2_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[39:20]),
          act_regs_data_1_1_sva_dfm_3, {nor_19_cse , while_asn_1374 , or_dcpl_122});
      act_regs_data_2_1_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_1_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[39:20]),
          act_regs_data_2_1_sva_dfm_3, {nor_20_cse , while_asn_1370 , or_dcpl_123});
      act_regs_data_3_1_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[39:20]),
          act_regs_data_3_1_sva_dfm_3, {nor_21_cse , while_asn_1366 , or_dcpl_124});
      act_regs_data_0_0_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_nor_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[19:0]),
          act_regs_data_0_0_sva_dfm_3, {nor_18_cse , while_asn_1378 , or_dcpl});
      act_regs_data_1_0_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_2_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[19:0]),
          act_regs_data_1_0_sva_dfm_3, {nor_19_cse , while_asn_1374 , or_dcpl_122});
      act_regs_data_2_0_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_1_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[19:0]),
          act_regs_data_2_0_sva_dfm_3, {nor_20_cse , while_asn_1370 , or_dcpl_123});
      act_regs_data_3_0_sva <= MUX1HOT_v_20_3_2((signext_20_1(~ ActUnit_RunLoad_if_else_and_ssc_sva_1)),
          (libraries_Adpfloat2Fixed_7fa345e634188c2e895631ad5a7aad3d14627_1[19:0]),
          act_regs_data_3_0_sva_dfm_3, {nor_21_cse , while_asn_1366 , or_dcpl_124});
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_config_adpfloat_bias_sva <= 3'b000;
      act_config_output_addr_base_sva <= 8'b00000000;
      act_config_buffer_addr_base_sva <= 5'b00000;
      act_config_num_inst_sva <= 6'b000001;
      act_config_num_output_sva <= 8'b00000001;
    end
    else if ( act_config_adpfloat_bias_and_cse ) begin
      act_config_adpfloat_bias_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[18:16];
      act_config_output_addr_base_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[71:64];
      act_config_buffer_addr_base_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[52:48];
      act_config_num_inst_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[29:24];
      act_config_num_output_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[39:32];
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_config_inst_regs_16_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_17_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_18_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_19_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_20_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_21_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_22_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_23_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_24_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_25_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_26_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_27_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_28_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_29_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_30_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_31_sva_dfm_6 <= 8'b00000000;
    end
    else if ( act_config_inst_regs_and_cse ) begin
      act_config_inst_regs_16_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[7:0];
      act_config_inst_regs_17_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[15:8];
      act_config_inst_regs_18_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[23:16];
      act_config_inst_regs_19_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[31:24];
      act_config_inst_regs_20_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[39:32];
      act_config_inst_regs_21_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[47:40];
      act_config_inst_regs_22_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[55:48];
      act_config_inst_regs_23_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[63:56];
      act_config_inst_regs_24_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[71:64];
      act_config_inst_regs_25_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[79:72];
      act_config_inst_regs_26_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[87:80];
      act_config_inst_regs_27_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[95:88];
      act_config_inst_regs_28_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[103:96];
      act_config_inst_regs_29_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[111:104];
      act_config_inst_regs_30_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[119:112];
      act_config_inst_regs_31_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[127:120];
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_config_inst_regs_0_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_1_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_2_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_3_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_4_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_5_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_6_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_7_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_8_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_9_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_10_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_11_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_12_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_13_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_14_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_15_sva_dfm_5 <= 8'b00000000;
    end
    else if ( act_config_inst_regs_and_16_cse ) begin
      act_config_inst_regs_0_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[7:0];
      act_config_inst_regs_1_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[15:8];
      act_config_inst_regs_2_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[23:16];
      act_config_inst_regs_3_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[31:24];
      act_config_inst_regs_4_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[39:32];
      act_config_inst_regs_5_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[47:40];
      act_config_inst_regs_6_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[55:48];
      act_config_inst_regs_7_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[63:56];
      act_config_inst_regs_8_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[71:64];
      act_config_inst_regs_9_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[79:72];
      act_config_inst_regs_10_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[87:80];
      act_config_inst_regs_11_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[95:88];
      act_config_inst_regs_12_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[103:96];
      act_config_inst_regs_13_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[111:104];
      act_config_inst_regs_14_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[119:112];
      act_config_inst_regs_15_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[127:120];
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_config_output_counter_sva <= 8'b00000000;
    end
    else if ( ActUnitRun_wen & ((~ or_dcpl_116) | (fsm_output[1]) | act_config_output_counter_sva_mx0c1)
        ) begin
      act_config_output_counter_sva <= MUX_v_8_2_2(8'b00000000, mux_91_nl, not_235_nl);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_0_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_0_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_0_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_0_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_0_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_0_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_0_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_0_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_0_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_0_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_0_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_0_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_0_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_0_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_0_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_0_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_cse ) begin
      act_mem_banks_bank_array_impl_data0_0_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_0_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_0_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_0_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_0_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_0_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_0_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_0_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_0_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_0_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_0_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_0_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_0_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_0_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_0_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_0_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_1_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_1_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_1_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_1_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_1_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_1_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_1_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_1_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_1_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_1_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_1_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_1_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_1_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_1_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_1_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_1_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_1_cse ) begin
      act_mem_banks_bank_array_impl_data0_1_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_1_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_1_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_1_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_1_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_1_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_1_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_1_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_1_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_1_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_1_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_1_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_1_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_1_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_1_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_1_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_2_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_2_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_2_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_2_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_2_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_2_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_2_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_2_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_2_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_2_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_2_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_2_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_2_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_2_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_2_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_2_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_2_cse ) begin
      act_mem_banks_bank_array_impl_data0_2_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_2_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_2_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_2_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_2_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_2_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_2_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_2_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_2_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_2_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_2_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_2_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_2_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_2_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_2_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_2_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_3_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_3_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_3_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_3_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_3_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_3_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_3_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_3_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_3_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_3_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_3_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_3_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_3_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_3_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_3_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_3_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_3_cse ) begin
      act_mem_banks_bank_array_impl_data0_3_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_3_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_3_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_3_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_3_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_3_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_3_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_3_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_3_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_3_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_3_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_3_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_3_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_3_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_3_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_3_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_4_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_4_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_4_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_4_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_4_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_4_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_4_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_4_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_4_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_4_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_4_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_4_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_4_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_4_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_4_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_4_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_4_cse ) begin
      act_mem_banks_bank_array_impl_data0_4_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_4_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_4_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_4_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_4_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_4_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_4_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_4_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_4_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_4_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_4_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_4_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_4_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_4_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_4_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_4_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_5_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_5_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_5_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_5_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_5_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_5_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_5_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_5_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_5_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_5_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_5_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_5_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_5_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_5_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_5_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_5_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_5_cse ) begin
      act_mem_banks_bank_array_impl_data0_5_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_5_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_5_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_5_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_5_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_5_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_5_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_5_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_5_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_5_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_5_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_5_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_5_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_5_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_5_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_5_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_6_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_6_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_6_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_6_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_6_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_6_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_6_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_6_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_6_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_6_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_6_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_6_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_6_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_6_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_6_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_6_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_6_cse ) begin
      act_mem_banks_bank_array_impl_data0_6_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_6_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_6_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_6_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_6_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_6_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_6_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_6_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_6_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_6_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_6_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_6_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_6_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_6_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_6_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_6_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_7_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_7_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_7_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_7_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_7_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_7_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_7_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_7_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_7_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_7_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_7_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_7_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_7_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_7_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_7_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_7_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_7_cse ) begin
      act_mem_banks_bank_array_impl_data0_7_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_7_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_7_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_7_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_7_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_7_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_7_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_7_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_7_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_7_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_7_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_7_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_7_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_7_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_7_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_7_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_8_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_8_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_8_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_8_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_8_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_8_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_8_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_8_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_8_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_8_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_8_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_8_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_8_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_8_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_8_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_8_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_8_cse ) begin
      act_mem_banks_bank_array_impl_data0_8_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_8_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_8_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_8_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_8_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_8_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_8_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_8_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_8_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_8_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_8_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_8_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_8_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_8_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_8_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_8_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_9_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_9_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_9_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_9_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_9_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_9_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_9_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_9_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_9_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_9_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_9_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_9_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_9_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_9_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_9_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_9_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_9_cse ) begin
      act_mem_banks_bank_array_impl_data0_9_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_9_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_9_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_9_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_9_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_9_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_9_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_9_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_9_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_9_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_9_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_9_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_9_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_9_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_9_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_9_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_10_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_10_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_10_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_10_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_10_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_10_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_10_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_10_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_10_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_10_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_10_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_10_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_10_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_10_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_10_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_10_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_10_cse ) begin
      act_mem_banks_bank_array_impl_data0_10_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_10_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_10_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_10_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_10_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_10_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_10_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_10_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_10_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_10_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_10_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_10_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_10_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_10_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_10_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_10_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_11_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_11_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_11_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_11_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_11_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_11_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_11_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_11_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_11_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_11_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_11_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_11_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_11_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_11_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_11_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_11_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_11_cse ) begin
      act_mem_banks_bank_array_impl_data0_11_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_11_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_11_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_11_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_11_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_11_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_11_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_11_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_11_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_11_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_11_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_11_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_11_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_11_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_11_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_11_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_12_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_12_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_12_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_12_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_12_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_12_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_12_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_12_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_12_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_12_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_12_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_12_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_12_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_12_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_12_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_12_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_12_cse ) begin
      act_mem_banks_bank_array_impl_data0_12_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_12_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_12_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_12_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_12_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_12_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_12_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_12_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_12_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_12_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_12_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_12_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_12_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_12_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_12_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_12_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_13_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_13_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_13_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_13_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_13_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_13_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_13_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_13_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_13_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_13_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_13_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_13_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_13_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_13_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_13_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_13_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_13_cse ) begin
      act_mem_banks_bank_array_impl_data0_13_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_13_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_13_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_13_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_13_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_13_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_13_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_13_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_13_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_13_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_13_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_13_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_13_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_13_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_13_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_13_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_14_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_14_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_14_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_14_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_14_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_14_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_14_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_14_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_14_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_14_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_14_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_14_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_14_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_14_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_14_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_14_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_14_cse ) begin
      act_mem_banks_bank_array_impl_data0_14_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_14_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_14_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_14_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_14_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_14_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_14_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_14_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_14_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_14_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_14_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_14_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_14_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_14_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_14_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_14_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_15_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_15_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_15_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_15_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_15_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_15_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_15_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_15_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_15_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_15_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_15_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_15_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_15_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_15_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_15_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_15_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_15_cse ) begin
      act_mem_banks_bank_array_impl_data0_15_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_15_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_15_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_15_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_15_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_15_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_15_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_15_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_15_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_15_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_15_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_15_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_15_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_15_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_15_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_15_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_16_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_16_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_16_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_16_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_16_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_16_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_16_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_16_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_16_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_16_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_16_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_16_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_16_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_16_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_16_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_16_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_16_cse ) begin
      act_mem_banks_bank_array_impl_data0_16_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_16_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_16_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_16_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_16_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_16_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_16_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_16_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_16_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_16_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_16_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_16_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_16_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_16_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_16_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_16_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_17_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_17_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_17_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_17_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_17_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_17_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_17_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_17_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_17_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_17_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_17_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_17_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_17_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_17_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_17_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_17_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_17_cse ) begin
      act_mem_banks_bank_array_impl_data0_17_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_17_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_17_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_17_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_17_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_17_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_17_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_17_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_17_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_17_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_17_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_17_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_17_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_17_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_17_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_17_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_18_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_18_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_18_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_18_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_18_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_18_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_18_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_18_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_18_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_18_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_18_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_18_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_18_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_18_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_18_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_18_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_18_cse ) begin
      act_mem_banks_bank_array_impl_data0_18_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_18_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_18_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_18_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_18_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_18_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_18_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_18_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_18_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_18_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_18_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_18_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_18_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_18_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_18_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_18_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_19_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_19_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_19_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_19_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_19_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_19_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_19_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_19_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_19_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_19_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_19_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_19_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_19_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_19_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_19_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_19_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_19_cse ) begin
      act_mem_banks_bank_array_impl_data0_19_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_19_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_19_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_19_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_19_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_19_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_19_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_19_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_19_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_19_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_19_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_19_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_19_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_19_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_19_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_19_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_20_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_20_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_20_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_20_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_20_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_20_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_20_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_20_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_20_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_20_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_20_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_20_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_20_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_20_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_20_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_20_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_20_cse ) begin
      act_mem_banks_bank_array_impl_data0_20_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_20_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_20_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_20_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_20_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_20_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_20_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_20_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_20_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_20_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_20_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_20_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_20_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_20_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_20_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_20_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_21_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_21_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_21_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_21_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_21_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_21_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_21_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_21_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_21_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_21_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_21_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_21_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_21_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_21_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_21_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_21_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_21_cse ) begin
      act_mem_banks_bank_array_impl_data0_21_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_21_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_21_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_21_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_21_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_21_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_21_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_21_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_21_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_21_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_21_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_21_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_21_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_21_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_21_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_21_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_22_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_22_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_22_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_22_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_22_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_22_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_22_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_22_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_22_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_22_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_22_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_22_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_22_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_22_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_22_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_22_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_22_cse ) begin
      act_mem_banks_bank_array_impl_data0_22_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_22_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_22_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_22_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_22_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_22_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_22_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_22_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_22_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_22_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_22_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_22_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_22_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_22_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_22_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_22_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_23_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_23_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_23_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_23_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_23_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_23_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_23_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_23_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_23_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_23_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_23_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_23_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_23_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_23_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_23_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_23_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_23_cse ) begin
      act_mem_banks_bank_array_impl_data0_23_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_23_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_23_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_23_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_23_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_23_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_23_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_23_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_23_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_23_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_23_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_23_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_23_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_23_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_23_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_23_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_24_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_24_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_24_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_24_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_24_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_24_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_24_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_24_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_24_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_24_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_24_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_24_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_24_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_24_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_24_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_24_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_24_cse ) begin
      act_mem_banks_bank_array_impl_data0_24_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_24_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_24_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_24_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_24_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_24_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_24_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_24_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_24_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_24_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_24_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_24_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_24_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_24_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_24_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_24_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_25_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_25_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_25_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_25_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_25_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_25_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_25_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_25_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_25_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_25_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_25_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_25_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_25_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_25_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_25_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_25_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_25_cse ) begin
      act_mem_banks_bank_array_impl_data0_25_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_25_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_25_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_25_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_25_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_25_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_25_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_25_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_25_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_25_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_25_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_25_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_25_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_25_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_25_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_25_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_26_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_26_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_26_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_26_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_26_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_26_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_26_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_26_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_26_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_26_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_26_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_26_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_26_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_26_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_26_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_26_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_26_cse ) begin
      act_mem_banks_bank_array_impl_data0_26_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_26_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_26_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_26_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_26_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_26_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_26_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_26_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_26_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_26_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_26_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_26_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_26_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_26_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_26_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_26_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_27_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_27_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_27_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_27_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_27_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_27_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_27_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_27_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_27_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_27_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_27_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_27_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_27_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_27_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_27_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_27_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_27_cse ) begin
      act_mem_banks_bank_array_impl_data0_27_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_27_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_27_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_27_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_27_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_27_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_27_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_27_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_27_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_27_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_27_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_27_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_27_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_27_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_27_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_27_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_28_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_28_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_28_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_28_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_28_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_28_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_28_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_28_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_28_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_28_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_28_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_28_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_28_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_28_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_28_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_28_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_28_cse ) begin
      act_mem_banks_bank_array_impl_data0_28_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_28_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_28_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_28_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_28_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_28_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_28_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_28_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_28_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_28_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_28_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_28_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_28_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_28_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_28_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_28_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_29_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_29_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_29_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_29_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_29_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_29_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_29_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_29_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_29_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_29_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_29_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_29_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_29_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_29_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_29_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_29_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_29_cse ) begin
      act_mem_banks_bank_array_impl_data0_29_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_29_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_29_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_29_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_29_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_29_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_29_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_29_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_29_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_29_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_29_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_29_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_29_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_29_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_29_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_29_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_30_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_30_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_30_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_30_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_30_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_30_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_30_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_30_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_30_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_30_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_30_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_30_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_30_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_30_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_30_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_30_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_30_cse ) begin
      act_mem_banks_bank_array_impl_data0_30_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_30_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_30_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_30_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_30_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_30_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_30_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_30_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_30_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_30_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_30_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_30_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_30_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_30_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_30_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_30_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_array_impl_data0_31_127_120_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_31_7_0_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_31_119_112_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_31_15_8_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_31_111_104_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_31_23_16_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_31_103_96_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_31_31_24_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_31_95_88_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_31_39_32_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_31_87_80_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_31_47_40_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_31_79_72_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_31_55_48_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_31_71_64_sva_dfm <= 8'b00000000;
      act_mem_banks_bank_array_impl_data0_31_63_56_sva_dfm <= 8'b00000000;
    end
    else if ( act_mem_banks_bank_array_impl_data0_and_31_cse ) begin
      act_mem_banks_bank_array_impl_data0_31_127_120_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_31_7_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_31_119_112_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_31_15_8_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_31_111_104_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_31_23_16_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_31_103_96_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_31_31_24_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_31_95_88_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_31_39_32_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_31_87_80_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_31_47_40_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_31_79_72_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_31_55_48_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_31_71_64_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_5_mx0;
      act_mem_banks_bank_array_impl_data0_31_63_56_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_5_mx0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      is_start_sva <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((is_start_sva & ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_cse
        & (fsm_output[1])) | is_start_sva_mx0c1) ) begin
      is_start_sva <= MUX_s_1_2_2(ActUnit_RunInst_switch_lp_equal_tmp_1, ActUnit_CheckStart_if_ActUnit_CheckStart_if_and_1_cse,
          is_start_sva_mx0c1);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_127_120 <= 8'b00000000;
      act_mem_banks_read_read_data_lpi_1_dfm_1_7_0 <= 8'b00000000;
      act_mem_banks_read_read_data_lpi_1_dfm_1_119_112 <= 8'b00000000;
      act_mem_banks_read_read_data_lpi_1_dfm_1_111_104 <= 8'b00000000;
      act_mem_banks_read_read_data_lpi_1_dfm_1_15_8 <= 8'b00000000;
      act_mem_banks_read_read_data_lpi_1_dfm_1_103_96 <= 8'b00000000;
      act_mem_banks_read_read_data_lpi_1_dfm_1_95_88 <= 8'b00000000;
      act_mem_banks_read_read_data_lpi_1_dfm_1_23_16 <= 8'b00000000;
      act_mem_banks_read_read_data_lpi_1_dfm_1_87_80 <= 8'b00000000;
      act_mem_banks_read_read_data_lpi_1_dfm_1_79_72 <= 8'b00000000;
      act_mem_banks_read_read_data_lpi_1_dfm_1_31_24 <= 8'b00000000;
      act_mem_banks_read_read_data_lpi_1_dfm_1_71_64 <= 8'b00000000;
      act_mem_banks_read_read_data_lpi_1_dfm_1_63_56 <= 8'b00000000;
      act_mem_banks_read_read_data_lpi_1_dfm_1_39_32 <= 8'b00000000;
      act_mem_banks_read_read_data_lpi_1_dfm_1_55_48 <= 8'b00000000;
      act_mem_banks_read_read_data_lpi_1_dfm_1_47_40 <= 8'b00000000;
    end
    else if ( act_mem_banks_read_read_data_and_cse ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_127_120 <= act_mem_banks_read_for_mux_mx0w0;
      act_mem_banks_read_read_data_lpi_1_dfm_1_7_0 <= act_mem_banks_read_for_mux_15_mx0w0;
      act_mem_banks_read_read_data_lpi_1_dfm_1_119_112 <= act_mem_banks_read_for_mux_1_mx0w0;
      act_mem_banks_read_read_data_lpi_1_dfm_1_111_104 <= act_mem_banks_read_for_mux_2_mx0w0;
      act_mem_banks_read_read_data_lpi_1_dfm_1_15_8 <= act_mem_banks_read_for_mux_14_mx0w0;
      act_mem_banks_read_read_data_lpi_1_dfm_1_103_96 <= act_mem_banks_read_for_mux_3_mx0w0;
      act_mem_banks_read_read_data_lpi_1_dfm_1_95_88 <= act_mem_banks_read_for_mux_4_mx0w0;
      act_mem_banks_read_read_data_lpi_1_dfm_1_23_16 <= act_mem_banks_read_for_mux_13_mx0w0;
      act_mem_banks_read_read_data_lpi_1_dfm_1_87_80 <= act_mem_banks_read_for_mux_5_mx0w0;
      act_mem_banks_read_read_data_lpi_1_dfm_1_79_72 <= act_mem_banks_read_for_mux_6_mx0w0;
      act_mem_banks_read_read_data_lpi_1_dfm_1_31_24 <= act_mem_banks_read_for_mux_12_mx0w0;
      act_mem_banks_read_read_data_lpi_1_dfm_1_71_64 <= act_mem_banks_read_for_mux_7_mx0w0;
      act_mem_banks_read_read_data_lpi_1_dfm_1_63_56 <= act_mem_banks_read_for_mux_8_mx0w0;
      act_mem_banks_read_read_data_lpi_1_dfm_1_39_32 <= act_mem_banks_read_for_mux_11_mx0w0;
      act_mem_banks_read_read_data_lpi_1_dfm_1_55_48 <= act_mem_banks_read_for_mux_9_mx0w0;
      act_mem_banks_read_read_data_lpi_1_dfm_1_47_40 <= act_mem_banks_read_for_mux_10_mx0w0;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_write_addrs_lpi_1_dfm_5 <= 5'b00000;
    end
    else if ( (~ mux_158_nl) & ActUnitRun_wen & ((mux_tmp_16 & and_dcpl_1 & (~ (act_config_in_InstFetch_mux_tmp[6]))
        & (~ (act_config_in_InstFetch_mux_tmp[4])) & (fsm_output[1])) | (nor_tmp_6
        & (fsm_output[2])) | act_write_addrs_lpi_1_dfm_5_mx0c2) ) begin
      act_write_addrs_lpi_1_dfm_5 <= MUX_v_5_2_2((z_out_7_0[4:0]), ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_3_mx0w2,
          act_write_addrs_lpi_1_dfm_5_mx0c2);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_cse <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((fsm_output[2:1]!=2'b00)) ) begin
      ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_cse <= ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_cse_1
          | (fsm_output[2]);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      ActUnit_RunInst_switch_lp_nor_7_itm <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((mux_tmp_16 & (fsm_output[1])) | (fsm_output[2]))
        ) begin
      ActUnit_RunInst_switch_lp_nor_7_itm <= MUX_s_1_2_2(ActUnit_RunInst_switch_lp_nor_7_itm_mx0w0,
          nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_31_nl, fsm_output[2]);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= 20'b00000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_18_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= 20'b00000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_19_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= 20'b00000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_20_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= 20'b00000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_21_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= 20'b00000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_22_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= 20'b00000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_23_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= 20'b00000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_24_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= 20'b00000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_25_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= 20'b00000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_26_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= 20'b00000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_27_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= 20'b00000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_28_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= 20'b00000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_29_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= 20'b00000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_30_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= 20'b00000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_31_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= 20'b00000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_32_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= 20'b00000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_33_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva
          <= nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_slc_act_regs_data_20_19_0_1_ctmp_sva_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      ActUnit_RunInst_case_8_EAdd_act_regs_data_sva <= 320'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ActUnitRun_wen & mux_tmp_1 & and_dcpl_5 & ActUnit_RunInst_switch_lp_nor_13_cse
        ) begin
      ActUnit_RunInst_case_8_EAdd_act_regs_data_sva <= libraries_EAdd_0d1aed8b807329bc366abb192bb53bb66056_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      ActUnit_RunInst_case_9_EMul_act_regs_data_sva <= 320'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ActUnitRun_wen & mux_tmp_1 & and_dcpl_5 & and_dcpl_8 ) begin
      ActUnit_RunInst_case_9_EMul_act_regs_data_sva <= libraries_EMul_50466378fb684d7351699b7bf1bdec8c6525_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva <= 320'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ActUnitRun_wen & mux_tmp_1 & and_dcpl_11 & ActUnit_RunInst_switch_lp_nor_13_cse
        ) begin
      ActUnit_RunInst_case_10_Sigmoid_act_regs_data_sva <= libraries_Sigmoid_6ea22cc51ee279163d827d3cc5db43491cd81_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      ActUnit_RunInst_case_11_Tanh_act_regs_data_sva <= 320'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ActUnitRun_wen & mux_tmp_1 & and_dcpl_11 & and_dcpl_8 ) begin
      ActUnit_RunInst_case_11_Tanh_act_regs_data_sva <= libraries_Tanh_0c47cc570305d1d8c1a9dd465101e61217b26_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      ActUnit_RunInst_case_12_Relu_act_regs_data_sva <= 320'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ActUnitRun_wen & mux_tmp_1 & and_dcpl_5 & (act_config_in_InstFetch_mux_tmp[6])
        & (~ (act_config_in_InstFetch_mux_tmp[4])) ) begin
      ActUnit_RunInst_case_12_Relu_act_regs_data_sva <= libraries_Relu_29d7978308309996bcf6431af85e65007d30_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      ActUnit_RunInst_case_13_OneX_act_regs_data_sva <= 320'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ActUnitRun_wen & mux_tmp_1 & and_dcpl_5 & and_dcpl ) begin
      ActUnit_RunInst_case_13_OneX_act_regs_data_sva <= libraries_OneX_6a9c88d8c3af0ca712acdf3bbda5530a55e7_1;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_write_data_data_0_15_lpi_1_dfm_4 <= 8'b00000000;
      act_write_data_data_0_14_lpi_1_dfm_4 <= 8'b00000000;
      act_write_data_data_0_13_lpi_1_dfm_4 <= 8'b00000000;
      act_write_data_data_0_12_lpi_1_dfm_4 <= 8'b00000000;
      act_write_data_data_0_11_lpi_1_dfm_4 <= 8'b00000000;
      act_write_data_data_0_10_lpi_1_dfm_4 <= 8'b00000000;
      act_write_data_data_0_9_lpi_1_dfm_4 <= 8'b00000000;
      act_write_data_data_0_8_lpi_1_dfm_4 <= 8'b00000000;
      act_write_data_data_0_7_lpi_1_dfm_4 <= 8'b00000000;
      act_write_data_data_0_6_lpi_1_dfm_4 <= 8'b00000000;
      act_write_data_data_0_5_lpi_1_dfm_4 <= 8'b00000000;
      act_write_data_data_0_4_lpi_1_dfm_4 <= 8'b00000000;
      act_write_data_data_0_3_lpi_1_dfm_4 <= 8'b00000000;
      act_write_data_data_0_2_lpi_1_dfm_4 <= 8'b00000000;
      act_write_data_data_0_1_lpi_1_dfm_4 <= 8'b00000000;
      act_write_data_data_0_0_lpi_1_dfm_4 <= 8'b00000000;
    end
    else if ( act_write_data_data_and_cse ) begin
      act_write_data_data_0_15_lpi_1_dfm_4 <= MUX_v_8_2_2(8'b00000000, (out_data_out[127:120]),
          ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0);
      act_write_data_data_0_14_lpi_1_dfm_4 <= MUX_v_8_2_2(8'b00000000, (out_data_out[119:112]),
          ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0);
      act_write_data_data_0_13_lpi_1_dfm_4 <= MUX_v_8_2_2(8'b00000000, (out_data_out[111:104]),
          ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0);
      act_write_data_data_0_12_lpi_1_dfm_4 <= MUX_v_8_2_2(8'b00000000, (out_data_out[103:96]),
          ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0);
      act_write_data_data_0_11_lpi_1_dfm_4 <= MUX_v_8_2_2(8'b00000000, (out_data_out[95:88]),
          ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0);
      act_write_data_data_0_10_lpi_1_dfm_4 <= MUX_v_8_2_2(8'b00000000, (out_data_out[87:80]),
          ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0);
      act_write_data_data_0_9_lpi_1_dfm_4 <= MUX_v_8_2_2(8'b00000000, (out_data_out[79:72]),
          ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0);
      act_write_data_data_0_8_lpi_1_dfm_4 <= MUX_v_8_2_2(8'b00000000, (out_data_out[71:64]),
          ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0);
      act_write_data_data_0_7_lpi_1_dfm_4 <= MUX_v_8_2_2(8'b00000000, (out_data_out[63:56]),
          ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0);
      act_write_data_data_0_6_lpi_1_dfm_4 <= MUX_v_8_2_2(8'b00000000, (out_data_out[55:48]),
          ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0);
      act_write_data_data_0_5_lpi_1_dfm_4 <= MUX_v_8_2_2(8'b00000000, (out_data_out[47:40]),
          ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0);
      act_write_data_data_0_4_lpi_1_dfm_4 <= MUX_v_8_2_2(8'b00000000, (out_data_out[39:32]),
          ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0);
      act_write_data_data_0_3_lpi_1_dfm_4 <= MUX_v_8_2_2(8'b00000000, (out_data_out[31:24]),
          ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0);
      act_write_data_data_0_2_lpi_1_dfm_4 <= MUX_v_8_2_2(8'b00000000, (out_data_out[23:16]),
          ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0);
      act_write_data_data_0_1_lpi_1_dfm_4 <= MUX_v_8_2_2(8'b00000000, (out_data_out[15:8]),
          ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0);
      act_write_data_data_0_0_lpi_1_dfm_4 <= MUX_v_8_2_2(8'b00000000, (out_data_out[7:0]),
          ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0);
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      act_read_addrs_lpi_1_dfm_5 <= 5'b00000;
    end
    else if ( ActUnitRun_wen & mux_4_nl ) begin
      act_read_addrs_lpi_1_dfm_5 <= (z_out_7_0[4:0]) & (signext_5_1(~ act_config_is_zero_first_sva))
          & ({{4{ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_cse_1}},
          ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_cse_1});
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_18_enex5
        ) begin
      reg_act_regs_data_3_15_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo <= 1'b1;
    end
    else if ( act_config_inst_regs_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_18_enex5
        ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo <= act_config_inst_regs_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo <= 1'b1;
    end
    else if ( act_config_inst_regs_and_16_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_18_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo <= act_config_inst_regs_and_16_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo <= 1'b1;
    end
    else if ( ActUnitRun_wen | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_18_enex5
        ) begin
      reg_act_config_inst_counter_enexo <= ActUnitRun_wen;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_1 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_19_enex5
        ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_1 <= act_config_inst_regs_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_19_enex5
        ) begin
      reg_act_regs_data_1_14_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_1 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_16_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_19_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_1 <= act_config_inst_regs_and_16_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_2 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_20_enex5
        ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_2 <= act_config_inst_regs_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_2 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_16_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_20_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_2 <= act_config_inst_regs_and_16_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_20_enex5
        ) begin
      reg_act_regs_data_1_13_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_3 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_21_enex5
        ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_3 <= act_config_inst_regs_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_3 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_16_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_21_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_3 <= act_config_inst_regs_and_16_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_21_enex5
        ) begin
      reg_act_regs_data_0_12_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_4 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_22_enex5
        ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_4 <= act_config_inst_regs_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_22_enex5
        ) begin
      reg_act_regs_data_0_11_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_4 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_16_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_22_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_4 <= act_config_inst_regs_and_16_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_5 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_23_enex5
        ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_5 <= act_config_inst_regs_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_5 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_16_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_23_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_5 <= act_config_inst_regs_and_16_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_23_enex5
        ) begin
      reg_act_regs_data_0_10_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_6 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_24_enex5
        ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_6 <= act_config_inst_regs_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_6 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_16_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_24_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_6 <= act_config_inst_regs_and_16_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_24_enex5
        ) begin
      reg_act_regs_data_3_9_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_7 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_25_enex5
        ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_7 <= act_config_inst_regs_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_25_enex5
        ) begin
      reg_act_regs_data_2_8_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_7 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_16_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_25_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_7 <= act_config_inst_regs_and_16_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_8 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_26_enex5
        ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_8 <= act_config_inst_regs_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_8 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_16_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_26_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_8 <= act_config_inst_regs_and_16_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_26_enex5
        ) begin
      reg_act_regs_data_0_7_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_9 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_27_enex5
        ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_9 <= act_config_inst_regs_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_9 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_16_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_27_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_9 <= act_config_inst_regs_and_16_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_27_enex5
        ) begin
      reg_act_regs_data_1_6_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_10 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_28_enex5
        ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_10 <= act_config_inst_regs_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_10 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_16_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_28_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_10 <= act_config_inst_regs_and_16_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_28_enex5
        ) begin
      reg_act_regs_data_3_5_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_11 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_29_enex5
        ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_11 <= act_config_inst_regs_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_29_enex5
        ) begin
      reg_act_regs_data_2_4_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_11 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_16_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_29_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_11 <= act_config_inst_regs_and_16_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_12 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_30_enex5
        ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_12 <= act_config_inst_regs_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_30_enex5
        ) begin
      reg_act_regs_data_3_3_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_12 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_16_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_30_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_12 <= act_config_inst_regs_and_16_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_13 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_31_enex5
        ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_13 <= act_config_inst_regs_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_31_enex5
        ) begin
      reg_act_regs_data_1_2_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_13 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_16_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_31_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_13 <= act_config_inst_regs_and_16_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_14 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_32_enex5
        ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_14 <= act_config_inst_regs_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_32_enex5
        ) begin
      reg_act_regs_data_0_1_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_14 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_16_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_32_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_14 <= act_config_inst_regs_and_16_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_15 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_33_enex5
        ) begin
      reg_act_config_inst_regs_19_sva_dfm_6_enexo_15 <= act_config_inst_regs_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_33_enex5
        ) begin
      reg_act_regs_data_1_0_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk ) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_15 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_16_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_2_for_and_33_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_15 <= act_config_inst_regs_and_16_cse;
    end
  end
  assign while_while_not_nl = ~ or_dcpl_116;
  assign while_while_while_or_nl = MUX_v_5_2_2((z_out_7_0[4:0]), 5'b11111, while_while_not_nl);
  assign mux_19_nl = MUX_s_1_2_2(or_884_itm, and_tmp, act_config_InstIncr_act_config_InstIncr_if_and_svs_1);
  assign and_1554_nl = MUX_v_5_2_2(5'b00000, while_while_while_or_nl, mux_19_nl);
  assign nand_6_nl = ~((fsm_output[2]) & (~ and_tmp));
  assign nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_2_nl = MUX_s_1_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[0]),
      (act_config_inst_regs_16_sva_dfm_6[0]), not_tmp_34);
  assign nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_33_nl = MUX_s_1_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[8]),
      (act_config_inst_regs_1_sva_dfm_5[0]), or_dcpl_27);
  assign nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_5_nl = MUX_s_1_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[8]),
      (act_config_inst_regs_17_sva_dfm_6[0]), not_tmp_34);
  assign while_else_1_while_else_1_nand_nl = ~(act_config_InstIncr_if_act_config_InstIncr_if_if_act_config_InstIncr_if_if_nor_mdf_sva_1
      & act_config_InstIncr_act_config_InstIncr_if_and_svs_1 & is_incr_lpi_1_dfm_2);
  assign act_config_InstIncr_if_act_config_InstIncr_if_and_1_nl = act_config_is_zero_first_sva
      & (~ act_config_InstIncr_if_act_config_InstIncr_if_if_act_config_InstIncr_if_if_nor_mdf_sva_1);
  assign act_config_ActConfigWrite_mux_33_nl = MUX_s_1_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[8]),
      act_config_is_zero_first_sva, act_config_ActConfigRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiWrite_mux_36_nl = MUX_s_1_2_2(act_config_ActConfigWrite_mux_33_nl,
      act_config_is_zero_first_sva, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxi_if_mux_82_nl = MUX_s_1_2_2(act_config_is_zero_first_sva,
      ActUnit_DecodeAxiWrite_mux_36_nl, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign ActUnit_DecodeAxi_mux_88_nl = MUX_s_1_2_2(act_config_is_zero_first_sva,
      ActUnit_DecodeAxi_if_mux_82_nl, rva_in_PopNB_mioi_return_rsc_z_mxwt);
  assign and_1557_nl = act_config_output_counter_sva_mx0c1 & (~ or_887_tmp);
  assign mux_91_nl = MUX_v_8_2_2(act_config_output_counter_sva, z_out_7_0, and_1557_nl);
  assign not_235_nl = ~ or_887_tmp;
  assign or_960_nl = is_start_sva | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt) | (~
      rva_in_PopNB_mioi_return_rsc_z_mxwt) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10:8]!=3'b001)
      | not_tmp_67;
  assign mux_156_nl = MUX_s_1_2_2(or_tmp_791, mux_tmp_118, is_start_sva);
  assign and_1734_nl = or_958_cse & or_tmp_791;
  assign and_1733_nl = or_957_cse & or_tmp_791;
  assign mux_149_nl = MUX_s_1_2_2(and_1734_nl, and_1733_nl, act_config_inst_counter_sva[0]);
  assign and_1732_nl = or_956_cse & or_tmp_791;
  assign and_1731_nl = or_955_cse & or_tmp_791;
  assign mux_148_nl = MUX_s_1_2_2(and_1732_nl, and_1731_nl, act_config_inst_counter_sva[0]);
  assign mux_150_nl = MUX_s_1_2_2(mux_149_nl, mux_148_nl, act_config_inst_counter_sva[1]);
  assign and_1730_nl = or_954_cse & or_tmp_791;
  assign and_1729_nl = or_953_cse & or_tmp_791;
  assign mux_146_nl = MUX_s_1_2_2(and_1730_nl, and_1729_nl, act_config_inst_counter_sva[0]);
  assign and_1728_nl = or_952_cse & or_tmp_791;
  assign and_1727_nl = or_951_cse & or_tmp_791;
  assign mux_145_nl = MUX_s_1_2_2(and_1728_nl, and_1727_nl, act_config_inst_counter_sva[0]);
  assign mux_147_nl = MUX_s_1_2_2(mux_146_nl, mux_145_nl, act_config_inst_counter_sva[1]);
  assign mux_151_nl = MUX_s_1_2_2(mux_150_nl, mux_147_nl, act_config_inst_counter_sva[2]);
  assign and_1726_nl = or_950_cse & or_tmp_791;
  assign and_1725_nl = or_949_cse & or_tmp_791;
  assign mux_142_nl = MUX_s_1_2_2(and_1726_nl, and_1725_nl, act_config_inst_counter_sva[0]);
  assign and_1724_nl = or_948_cse & or_tmp_791;
  assign and_1723_nl = or_947_cse & or_tmp_791;
  assign mux_141_nl = MUX_s_1_2_2(and_1724_nl, and_1723_nl, act_config_inst_counter_sva[0]);
  assign mux_143_nl = MUX_s_1_2_2(mux_142_nl, mux_141_nl, act_config_inst_counter_sva[1]);
  assign and_1722_nl = or_946_cse & or_tmp_791;
  assign and_1721_nl = or_945_cse & or_tmp_791;
  assign mux_139_nl = MUX_s_1_2_2(and_1722_nl, and_1721_nl, act_config_inst_counter_sva[0]);
  assign and_1720_nl = or_944_cse & or_tmp_791;
  assign and_1719_nl = or_943_cse & or_tmp_791;
  assign mux_138_nl = MUX_s_1_2_2(and_1720_nl, and_1719_nl, act_config_inst_counter_sva[0]);
  assign mux_140_nl = MUX_s_1_2_2(mux_139_nl, mux_138_nl, act_config_inst_counter_sva[1]);
  assign mux_144_nl = MUX_s_1_2_2(mux_143_nl, mux_140_nl, act_config_inst_counter_sva[2]);
  assign mux_152_nl = MUX_s_1_2_2(mux_151_nl, mux_144_nl, act_config_inst_counter_sva[3]);
  assign and_1718_nl = or_942_cse & or_tmp_791;
  assign and_1717_nl = or_941_cse & or_tmp_791;
  assign mux_134_nl = MUX_s_1_2_2(and_1718_nl, and_1717_nl, act_config_inst_counter_sva[0]);
  assign and_1716_nl = or_940_cse & or_tmp_791;
  assign and_1715_nl = or_939_cse & or_tmp_791;
  assign mux_133_nl = MUX_s_1_2_2(and_1716_nl, and_1715_nl, act_config_inst_counter_sva[0]);
  assign mux_135_nl = MUX_s_1_2_2(mux_134_nl, mux_133_nl, act_config_inst_counter_sva[1]);
  assign and_1714_nl = or_938_cse & or_tmp_791;
  assign and_1713_nl = or_937_cse & or_tmp_791;
  assign mux_131_nl = MUX_s_1_2_2(and_1714_nl, and_1713_nl, act_config_inst_counter_sva[0]);
  assign and_1712_nl = or_936_cse & or_tmp_791;
  assign and_1711_nl = or_935_cse & or_tmp_791;
  assign mux_130_nl = MUX_s_1_2_2(and_1712_nl, and_1711_nl, act_config_inst_counter_sva[0]);
  assign mux_132_nl = MUX_s_1_2_2(mux_131_nl, mux_130_nl, act_config_inst_counter_sva[1]);
  assign mux_136_nl = MUX_s_1_2_2(mux_135_nl, mux_132_nl, act_config_inst_counter_sva[2]);
  assign and_1710_nl = or_934_cse & or_tmp_791;
  assign and_1709_nl = or_933_cse & or_tmp_791;
  assign mux_127_nl = MUX_s_1_2_2(and_1710_nl, and_1709_nl, act_config_inst_counter_sva[0]);
  assign and_1708_nl = or_932_cse & or_tmp_791;
  assign and_1707_nl = or_931_cse & or_tmp_791;
  assign mux_126_nl = MUX_s_1_2_2(and_1708_nl, and_1707_nl, act_config_inst_counter_sva[0]);
  assign mux_128_nl = MUX_s_1_2_2(mux_127_nl, mux_126_nl, act_config_inst_counter_sva[1]);
  assign and_1706_nl = or_930_cse & or_tmp_791;
  assign and_1705_nl = or_929_cse & or_tmp_791;
  assign mux_124_nl = MUX_s_1_2_2(and_1706_nl, and_1705_nl, act_config_inst_counter_sva[0]);
  assign and_1704_nl = or_928_cse & or_tmp_791;
  assign and_1703_nl = or_925_cse & or_tmp_791;
  assign mux_123_nl = MUX_s_1_2_2(and_1704_nl, and_1703_nl, act_config_inst_counter_sva[0]);
  assign mux_125_nl = MUX_s_1_2_2(mux_124_nl, mux_123_nl, act_config_inst_counter_sva[1]);
  assign mux_129_nl = MUX_s_1_2_2(mux_128_nl, mux_125_nl, act_config_inst_counter_sva[2]);
  assign mux_137_nl = MUX_s_1_2_2(mux_136_nl, mux_129_nl, act_config_inst_counter_sva[3]);
  assign mux_153_nl = MUX_s_1_2_2(mux_152_nl, mux_137_nl, act_config_inst_counter_sva[4]);
  assign mux_154_nl = MUX_s_1_2_2(or_tmp_791, mux_153_nl, ActUnit_CheckStart_if_ActUnit_CheckStart_if_and_1_cse);
  assign nand_nl = ~(ActUnit_RunInst_switch_lp_equal_tmp_1 & (~ mux_tmp_118));
  assign mux_155_nl = MUX_s_1_2_2(mux_154_nl, nand_nl, is_start_sva);
  assign mux_157_nl = MUX_s_1_2_2(mux_156_nl, mux_155_nl, ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_cse);
  assign mux_158_nl = MUX_s_1_2_2(or_960_nl, mux_157_nl, fsm_output[1]);
  assign nvhls_get_slc_8U_nvhls_nvhls_t_128U_nvuint_t_4_mux_31_nl = MUX_s_1_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[0]),
      (act_config_inst_regs_0_sva_dfm_5[0]), or_dcpl_27);
  assign nor_16_nl = ~((act_config_in_InstFetch_mux_tmp[5]) | (~ mux_tmp_1));
  assign or_1_nl = (act_config_in_InstFetch_mux_tmp[4]) | (act_config_in_InstFetch_mux_tmp[6])
      | (act_config_in_InstFetch_mux_tmp[7]);
  assign mux_4_nl = MUX_s_1_2_2(nor_16_nl, mux_tmp_1, or_1_nl);
  assign operator_8_false_nor_1_nl = ~(or_tmp_756 | (fsm_output[1]));
  assign operator_8_false_operator_8_false_and_1_nl = MUX_v_3_2_2(3'b000, (act_config_output_counter_sva[7:5]),
      operator_8_false_nor_1_nl);
  assign operator_8_false_operator_8_false_mux_2_nl = MUX_v_5_2_2((act_config_output_counter_sva[4:0]),
      act_config_inst_counter_sva, or_tmp_756);
  assign operator_8_false_operator_8_false_mux_3_nl = MUX_v_5_2_2(5'b00001, act_config_buffer_addr_base_sva,
      fsm_output[1]);
  assign nl_z_out_7_0 = ({operator_8_false_operator_8_false_and_1_nl , operator_8_false_operator_8_false_mux_2_nl})
      + conv_u2u_5_8(operator_8_false_operator_8_false_mux_3_nl);
  assign z_out_7_0 = nl_z_out_7_0[7:0];

  function automatic [0:0] MUX1HOT_s_1_1_2;
    input [0:0] input_0;
    input [0:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    MUX1HOT_s_1_1_2 = result;
  end
  endfunction


  function automatic [19:0] MUX1HOT_v_20_3_2;
    input [19:0] input_2;
    input [19:0] input_1;
    input [19:0] input_0;
    input [2:0] sel;
    reg [19:0] result;
  begin
    result = input_0 & {20{sel[0]}};
    result = result | ( input_1 & {20{sel[1]}});
    result = result | ( input_2 & {20{sel[2]}});
    MUX1HOT_v_20_3_2 = result;
  end
  endfunction


  function automatic [19:0] MUX1HOT_v_20_5_2;
    input [19:0] input_4;
    input [19:0] input_3;
    input [19:0] input_2;
    input [19:0] input_1;
    input [19:0] input_0;
    input [4:0] sel;
    reg [19:0] result;
  begin
    result = input_0 & {20{sel[0]}};
    result = result | ( input_1 & {20{sel[1]}});
    result = result | ( input_2 & {20{sel[2]}});
    result = result | ( input_3 & {20{sel[3]}});
    result = result | ( input_4 & {20{sel[4]}});
    MUX1HOT_v_20_5_2 = result;
  end
  endfunction


  function automatic [19:0] MUX1HOT_v_20_9_2;
    input [19:0] input_8;
    input [19:0] input_7;
    input [19:0] input_6;
    input [19:0] input_5;
    input [19:0] input_4;
    input [19:0] input_3;
    input [19:0] input_2;
    input [19:0] input_1;
    input [19:0] input_0;
    input [8:0] sel;
    reg [19:0] result;
  begin
    result = input_0 & {20{sel[0]}};
    result = result | ( input_1 & {20{sel[1]}});
    result = result | ( input_2 & {20{sel[2]}});
    result = result | ( input_3 & {20{sel[3]}});
    result = result | ( input_4 & {20{sel[4]}});
    result = result | ( input_5 & {20{sel[5]}});
    result = result | ( input_6 & {20{sel[6]}});
    result = result | ( input_7 & {20{sel[7]}});
    result = result | ( input_8 & {20{sel[8]}});
    MUX1HOT_v_20_9_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_4_2;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [3:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    result = result | ( input_3 & {3{sel[3]}});
    MUX1HOT_v_3_4_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_4_2;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [3:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | ( input_1 & {5{sel[1]}});
    result = result | ( input_2 & {5{sel[2]}});
    result = result | ( input_3 & {5{sel[3]}});
    MUX1HOT_v_5_4_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_4_2;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [3:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | ( input_1 & {6{sel[1]}});
    result = result | ( input_2 & {6{sel[2]}});
    result = result | ( input_3 & {6{sel[3]}});
    MUX1HOT_v_6_4_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_4_2;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [3:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    result = result | ( input_3 & {8{sel[3]}});
    MUX1HOT_v_8_4_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [19:0] MUX_v_20_4_2;
    input [19:0] input_0;
    input [19:0] input_1;
    input [19:0] input_2;
    input [19:0] input_3;
    input [1:0] sel;
    reg [19:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_20_4_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_32_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [1:0] input_2;
    input [1:0] input_3;
    input [1:0] input_4;
    input [1:0] input_5;
    input [1:0] input_6;
    input [1:0] input_7;
    input [1:0] input_8;
    input [1:0] input_9;
    input [1:0] input_10;
    input [1:0] input_11;
    input [1:0] input_12;
    input [1:0] input_13;
    input [1:0] input_14;
    input [1:0] input_15;
    input [1:0] input_16;
    input [1:0] input_17;
    input [1:0] input_18;
    input [1:0] input_19;
    input [1:0] input_20;
    input [1:0] input_21;
    input [1:0] input_22;
    input [1:0] input_23;
    input [1:0] input_24;
    input [1:0] input_25;
    input [1:0] input_26;
    input [1:0] input_27;
    input [1:0] input_28;
    input [1:0] input_29;
    input [1:0] input_30;
    input [1:0] input_31;
    input [4:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      5'b00000 : begin
        result = input_0;
      end
      5'b00001 : begin
        result = input_1;
      end
      5'b00010 : begin
        result = input_2;
      end
      5'b00011 : begin
        result = input_3;
      end
      5'b00100 : begin
        result = input_4;
      end
      5'b00101 : begin
        result = input_5;
      end
      5'b00110 : begin
        result = input_6;
      end
      5'b00111 : begin
        result = input_7;
      end
      5'b01000 : begin
        result = input_8;
      end
      5'b01001 : begin
        result = input_9;
      end
      5'b01010 : begin
        result = input_10;
      end
      5'b01011 : begin
        result = input_11;
      end
      5'b01100 : begin
        result = input_12;
      end
      5'b01101 : begin
        result = input_13;
      end
      5'b01110 : begin
        result = input_14;
      end
      5'b01111 : begin
        result = input_15;
      end
      5'b10000 : begin
        result = input_16;
      end
      5'b10001 : begin
        result = input_17;
      end
      5'b10010 : begin
        result = input_18;
      end
      5'b10011 : begin
        result = input_19;
      end
      5'b10100 : begin
        result = input_20;
      end
      5'b10101 : begin
        result = input_21;
      end
      5'b10110 : begin
        result = input_22;
      end
      5'b10111 : begin
        result = input_23;
      end
      5'b11000 : begin
        result = input_24;
      end
      5'b11001 : begin
        result = input_25;
      end
      5'b11010 : begin
        result = input_26;
      end
      5'b11011 : begin
        result = input_27;
      end
      5'b11100 : begin
        result = input_28;
      end
      5'b11101 : begin
        result = input_29;
      end
      5'b11110 : begin
        result = input_30;
      end
      default : begin
        result = input_31;
      end
    endcase
    MUX_v_2_32_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_32_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [7:0] input_8;
    input [7:0] input_9;
    input [7:0] input_10;
    input [7:0] input_11;
    input [7:0] input_12;
    input [7:0] input_13;
    input [7:0] input_14;
    input [7:0] input_15;
    input [7:0] input_16;
    input [7:0] input_17;
    input [7:0] input_18;
    input [7:0] input_19;
    input [7:0] input_20;
    input [7:0] input_21;
    input [7:0] input_22;
    input [7:0] input_23;
    input [7:0] input_24;
    input [7:0] input_25;
    input [7:0] input_26;
    input [7:0] input_27;
    input [7:0] input_28;
    input [7:0] input_29;
    input [7:0] input_30;
    input [7:0] input_31;
    input [4:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      5'b00000 : begin
        result = input_0;
      end
      5'b00001 : begin
        result = input_1;
      end
      5'b00010 : begin
        result = input_2;
      end
      5'b00011 : begin
        result = input_3;
      end
      5'b00100 : begin
        result = input_4;
      end
      5'b00101 : begin
        result = input_5;
      end
      5'b00110 : begin
        result = input_6;
      end
      5'b00111 : begin
        result = input_7;
      end
      5'b01000 : begin
        result = input_8;
      end
      5'b01001 : begin
        result = input_9;
      end
      5'b01010 : begin
        result = input_10;
      end
      5'b01011 : begin
        result = input_11;
      end
      5'b01100 : begin
        result = input_12;
      end
      5'b01101 : begin
        result = input_13;
      end
      5'b01110 : begin
        result = input_14;
      end
      5'b01111 : begin
        result = input_15;
      end
      5'b10000 : begin
        result = input_16;
      end
      5'b10001 : begin
        result = input_17;
      end
      5'b10010 : begin
        result = input_18;
      end
      5'b10011 : begin
        result = input_19;
      end
      5'b10100 : begin
        result = input_20;
      end
      5'b10101 : begin
        result = input_21;
      end
      5'b10110 : begin
        result = input_22;
      end
      5'b10111 : begin
        result = input_23;
      end
      5'b11000 : begin
        result = input_24;
      end
      5'b11001 : begin
        result = input_25;
      end
      5'b11010 : begin
        result = input_26;
      end
      5'b11011 : begin
        result = input_27;
      end
      5'b11100 : begin
        result = input_28;
      end
      5'b11101 : begin
        result = input_29;
      end
      5'b11110 : begin
        result = input_30;
      end
      default : begin
        result = input_31;
      end
    endcase
    MUX_v_8_32_2 = result;
  end
  endfunction


  function automatic [19:0] signext_20_1;
    input [0:0] vector;
  begin
    signext_20_1= {{19{vector[0]}}, vector};
  end
  endfunction


  function automatic [1:0] signext_2_1;
    input [0:0] vector;
  begin
    signext_2_1= {{1{vector[0]}}, vector};
  end
  endfunction


  function automatic [2:0] signext_3_1;
    input [0:0] vector;
  begin
    signext_3_1= {{2{vector[0]}}, vector};
  end
  endfunction


  function automatic [4:0] signext_5_1;
    input [0:0] vector;
  begin
    signext_5_1= {{4{vector[0]}}, vector};
  end
  endfunction


  function automatic [6:0] signext_7_1;
    input [0:0] vector;
  begin
    signext_7_1= {{6{vector[0]}}, vector};
  end
  endfunction


  function automatic [7:0] signext_8_1;
    input [0:0] vector;
  begin
    signext_8_1= {{7{vector[0]}}, vector};
  end
  endfunction


  function automatic [6:0] conv_u2s_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2s_6_7 =  {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_5_8 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_8 = {{3{1'b0}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit
// ------------------------------------------------------------------


module ActUnit (
  clk, rst, start_val, start_rdy, start_msg, act_port_val, act_port_rdy, act_port_msg,
      rva_in_val, rva_in_rdy, rva_in_msg, rva_out_val, rva_out_rdy, rva_out_msg,
      output_port_val, output_port_rdy, output_port_msg, done_val, done_rdy, done_msg
);
  input clk;
  input rst;
  input start_val;
  output start_rdy;
  input start_msg;
  input act_port_val;
  output act_port_rdy;
  input [319:0] act_port_msg;
  input rva_in_val;
  output rva_in_rdy;
  input [168:0] rva_in_msg;
  output rva_out_val;
  input rva_out_rdy;
  output [127:0] rva_out_msg;
  output output_port_val;
  input output_port_rdy;
  output [137:0] output_port_msg;
  output done_val;
  input done_rdy;
  output done_msg;

    // helpful signals for verification

    wire is_start = run.is_start_sva;
    wire [2:0] state = is_start ? (run.fsm_output[1]? 3'b010:3'b001) : 3'b000;

    // Act_config
    wire act_config_is_valid = run.act_config_is_valid_sva;
    wire act_config_is_zero_first = run.act_config_is_zero_first_sva;
    wire [2:0] act_config_adpfloat_bias = run.act_config_adpfloat_bias_sva;
    wire [5:0] act_config_num_inst = run.act_config_num_inst_sva;
    wire [7:0] act_config_num_output = run.act_config_num_output_sva;
    wire [4:0] act_config_buffer_addr_base = run.act_config_buffer_addr_base_sva;
    wire [7:0] act_config_output_addr_base = run.act_config_output_addr_base_sva;
    wire [4:0] act_config_inst_counter = run.act_config_inst_counter_sva;
    wire [7:0] act_config_output_counter = run.act_config_output_counter_sva;



  // Interconnect Declarations for Component Instantiations 
  ActUnit_ActUnit_ActUnitRun run (
      .clk(clk),
      .rst(rst),
      .start_val(start_val),
      .start_rdy(start_rdy),
      .start_msg(start_msg),
      .act_port_val(act_port_val),
      .act_port_rdy(act_port_rdy),
      .act_port_msg(act_port_msg),
      .rva_in_val(rva_in_val),
      .rva_in_rdy(rva_in_rdy),
      .rva_in_msg(rva_in_msg),
      .rva_out_val(rva_out_val),
      .rva_out_rdy(rva_out_rdy),
      .rva_out_msg(rva_out_msg),
      .output_port_val(output_port_val),
      .output_port_rdy(output_port_rdy),
      .output_port_msg(output_port_msg),
      .done_val(done_val),
      .done_rdy(done_rdy),
      .done_msg(done_msg)
    );
endmodule



