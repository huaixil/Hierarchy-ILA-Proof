module DATAPATH(
__ILA_DATAPATH_grant__,
alu_op,
bit_addr,
bit_in,
clk,
cy_sel,
nondet_des1_func_n3936,
nondet_desCy_func_n3988,
nondet_des_acc_func_n3499,
nondet_div_des1_n4958,
nondet_div_des2_n4955,
nondet_mul_des1_n4947,
nondet_mul_des2_n4944,
nondet_psw_next_func_n3704,
op2,
op3,
p,
pc,
psw_set,
ram_rd_sel,
ram_wr_sel,
rd_addr,
rst,
src_sel1,
src_sel2,
src_sel3,
wr,
wr_addr,
wr_ind,
wr_sfr,
__ILA_DATAPATH_acc_decode__,
__ILA_DATAPATH_decode_of_alu_add__,
__ILA_DATAPATH_decode_of_alu_and__,
__ILA_DATAPATH_decode_of_alu_da__,
__ILA_DATAPATH_decode_of_alu_div__,
__ILA_DATAPATH_decode_of_alu_inc__,
__ILA_DATAPATH_decode_of_alu_mul__,
__ILA_DATAPATH_decode_of_alu_not__,
__ILA_DATAPATH_decode_of_alu_or__,
__ILA_DATAPATH_decode_of_alu_rl__,
__ILA_DATAPATH_decode_of_alu_rlc__,
__ILA_DATAPATH_decode_of_alu_rr__,
__ILA_DATAPATH_decode_of_alu_rrc__,
__ILA_DATAPATH_decode_of_alu_sub__,
__ILA_DATAPATH_decode_of_alu_xch__,
__ILA_DATAPATH_decode_of_alu_xor__,
__ILA_DATAPATH_decode_of_no_wr__,
__ILA_DATAPATH_decode_of_read_data__,
__ILA_DATAPATH_decode_of_wr_ram__,
__ILA_DATAPATH_decode_of_wr_sfr__,
__ILA_DATAPATH_decode_of_wr_sfr_ram__,
__ILA_DATAPATH_valid__,
bit_addr_r,
wait_data,
bit_address,
ram_rd_data,
sfr_rd_data,
sfr_bit_rd_data,
ram_bit_rd_data,
rd_addr_r,
wr_addr_r,
wr_bit_r,
ram_wr_sel_r,
sfr_wr_addr_r,
rd_ind,
acc,
b_reg,
sp,
pop,
dptr_hi,
dptr_lo,
psw,
p0,
p1,
p2,
p3,
tcon,
scon,
ip,
ie,
pcon,
sbuf,
th0,
th1,
tl0,
tl1,
tmod,
op2_reg,
op3_reg,
iram_0,
iram_1,
iram_2,
iram_3,
iram_4,
iram_5,
iram_6,
iram_7,
iram_8,
iram_9,
iram_10,
iram_11,
iram_12,
iram_13,
iram_14,
iram_15,
iram_16,
iram_17,
iram_18,
iram_19,
iram_20,
iram_21,
iram_22,
iram_23,
iram_24,
iram_25,
iram_26,
iram_27,
iram_28,
iram_29,
iram_30,
iram_31,
iram_32,
iram_33,
iram_34,
iram_35,
iram_36,
iram_37,
iram_38,
iram_39,
iram_40,
iram_41,
iram_42,
iram_43,
iram_44,
iram_45,
iram_46,
iram_47,
iram_48,
iram_49,
iram_50,
iram_51,
iram_52,
iram_53,
iram_54,
iram_55,
iram_56,
iram_57,
iram_58,
iram_59,
iram_60,
iram_61,
iram_62,
iram_63,
iram_64,
iram_65,
iram_66,
iram_67,
iram_68,
iram_69,
iram_70,
iram_71,
iram_72,
iram_73,
iram_74,
iram_75,
iram_76,
iram_77,
iram_78,
iram_79,
iram_80,
iram_81,
iram_82,
iram_83,
iram_84,
iram_85,
iram_86,
iram_87,
iram_88,
iram_89,
iram_90,
iram_91,
iram_92,
iram_93,
iram_94,
iram_95,
iram_96,
iram_97,
iram_98,
iram_99,
iram_100,
iram_101,
iram_102,
iram_103,
iram_104,
iram_105,
iram_106,
iram_107,
iram_108,
iram_109,
iram_110,
iram_111,
iram_112,
iram_113,
iram_114,
iram_115,
iram_116,
iram_117,
iram_118,
iram_119,
iram_120,
iram_121,
iram_122,
iram_123,
iram_124,
iram_125,
iram_126,
iram_127,
iram_128,
iram_129,
iram_130,
iram_131,
iram_132,
iram_133,
iram_134,
iram_135,
iram_136,
iram_137,
iram_138,
iram_139,
iram_140,
iram_141,
iram_142,
iram_143,
iram_144,
iram_145,
iram_146,
iram_147,
iram_148,
iram_149,
iram_150,
iram_151,
iram_152,
iram_153,
iram_154,
iram_155,
iram_156,
iram_157,
iram_158,
iram_159,
iram_160,
iram_161,
iram_162,
iram_163,
iram_164,
iram_165,
iram_166,
iram_167,
iram_168,
iram_169,
iram_170,
iram_171,
iram_172,
iram_173,
iram_174,
iram_175,
iram_176,
iram_177,
iram_178,
iram_179,
iram_180,
iram_181,
iram_182,
iram_183,
iram_184,
iram_185,
iram_186,
iram_187,
iram_188,
iram_189,
iram_190,
iram_191,
iram_192,
iram_193,
iram_194,
iram_195,
iram_196,
iram_197,
iram_198,
iram_199,
iram_200,
iram_201,
iram_202,
iram_203,
iram_204,
iram_205,
iram_206,
iram_207,
iram_208,
iram_209,
iram_210,
iram_211,
iram_212,
iram_213,
iram_214,
iram_215,
iram_216,
iram_217,
iram_218,
iram_219,
iram_220,
iram_221,
iram_222,
iram_223,
iram_224,
iram_225,
iram_226,
iram_227,
iram_228,
iram_229,
iram_230,
iram_231,
iram_232,
iram_233,
iram_234,
iram_235,
iram_236,
iram_237,
iram_238,
iram_239,
iram_240,
iram_241,
iram_242,
iram_243,
iram_244,
iram_245,
iram_246,
iram_247,
iram_248,
iram_249,
iram_250,
iram_251,
iram_252,
iram_253,
iram_254,
iram_255
);
input     [19:0] __ILA_DATAPATH_grant__;
input      [3:0] alu_op;
input            bit_addr;
input            bit_in;
input            clk;
input      [1:0] cy_sel;
input      [7:0] nondet_des1_func_n3936;
input            nondet_desCy_func_n3988;
input      [7:0] nondet_des_acc_func_n3499;
input      [7:0] nondet_div_des1_n4958;
input      [7:0] nondet_div_des2_n4955;
input      [7:0] nondet_mul_des1_n4947;
input      [7:0] nondet_mul_des2_n4944;
input      [7:0] nondet_psw_next_func_n3704;
input      [7:0] op2;
input      [7:0] op3;
input            p;
input     [15:0] pc;
input      [1:0] psw_set;
input      [2:0] ram_rd_sel;
input      [2:0] ram_wr_sel;
input      [7:0] rd_addr;
input            rst;
input      [2:0] src_sel1;
input      [1:0] src_sel2;
input            src_sel3;
input            wr;
input      [7:0] wr_addr;
input            wr_ind;
input      [1:0] wr_sfr;
output     [19:0] __ILA_DATAPATH_acc_decode__;
output            __ILA_DATAPATH_decode_of_alu_add__;
output            __ILA_DATAPATH_decode_of_alu_and__;
output            __ILA_DATAPATH_decode_of_alu_da__;
output            __ILA_DATAPATH_decode_of_alu_div__;
output            __ILA_DATAPATH_decode_of_alu_inc__;
output            __ILA_DATAPATH_decode_of_alu_mul__;
output            __ILA_DATAPATH_decode_of_alu_not__;
output            __ILA_DATAPATH_decode_of_alu_or__;
output            __ILA_DATAPATH_decode_of_alu_rl__;
output            __ILA_DATAPATH_decode_of_alu_rlc__;
output            __ILA_DATAPATH_decode_of_alu_rr__;
output            __ILA_DATAPATH_decode_of_alu_rrc__;
output            __ILA_DATAPATH_decode_of_alu_sub__;
output            __ILA_DATAPATH_decode_of_alu_xch__;
output            __ILA_DATAPATH_decode_of_alu_xor__;
output            __ILA_DATAPATH_decode_of_no_wr__;
output            __ILA_DATAPATH_decode_of_read_data__;
output            __ILA_DATAPATH_decode_of_wr_ram__;
output            __ILA_DATAPATH_decode_of_wr_sfr__;
output            __ILA_DATAPATH_decode_of_wr_sfr_ram__;
output            __ILA_DATAPATH_valid__;
output reg            bit_addr_r;
output reg            wait_data;
output reg      [2:0] bit_address;
output reg      [7:0] ram_rd_data;
output reg      [7:0] sfr_rd_data;
output reg            sfr_bit_rd_data;
output reg            ram_bit_rd_data;
output reg            rd_addr_r;
output reg      [7:0] wr_addr_r;
output reg            wr_bit_r;
output reg      [2:0] ram_wr_sel_r;
output reg      [7:0] sfr_wr_addr_r;
output reg            rd_ind;
output reg      [7:0] acc;
output reg      [7:0] b_reg;
output reg      [7:0] sp;
output reg            pop;
output reg      [7:0] dptr_hi;
output reg      [7:0] dptr_lo;
output reg      [6:0] psw;
output reg      [7:0] p0;
output reg      [7:0] p1;
output reg      [7:0] p2;
output reg      [7:0] p3;
output reg      [7:0] tcon;
output reg      [7:0] scon;
output reg      [7:0] ip;
output reg      [7:0] ie;
output reg      [7:0] pcon;
output reg      [7:0] sbuf;
output reg      [7:0] th0;
output reg      [7:0] th1;
output reg      [7:0] tl0;
output reg      [7:0] tl1;
output reg      [7:0] tmod;
output reg      [7:0] op2_reg;
output reg      [7:0] op3_reg;
output reg      [7:0] iram_0;
output reg      [7:0] iram_1;
output reg      [7:0] iram_2;
output reg      [7:0] iram_3;
output reg      [7:0] iram_4;
output reg      [7:0] iram_5;
output reg      [7:0] iram_6;
output reg      [7:0] iram_7;
output reg      [7:0] iram_8;
output reg      [7:0] iram_9;
output reg      [7:0] iram_10;
output reg      [7:0] iram_11;
output reg      [7:0] iram_12;
output reg      [7:0] iram_13;
output reg      [7:0] iram_14;
output reg      [7:0] iram_15;
output reg      [7:0] iram_16;
output reg      [7:0] iram_17;
output reg      [7:0] iram_18;
output reg      [7:0] iram_19;
output reg      [7:0] iram_20;
output reg      [7:0] iram_21;
output reg      [7:0] iram_22;
output reg      [7:0] iram_23;
output reg      [7:0] iram_24;
output reg      [7:0] iram_25;
output reg      [7:0] iram_26;
output reg      [7:0] iram_27;
output reg      [7:0] iram_28;
output reg      [7:0] iram_29;
output reg      [7:0] iram_30;
output reg      [7:0] iram_31;
output reg      [7:0] iram_32;
output reg      [7:0] iram_33;
output reg      [7:0] iram_34;
output reg      [7:0] iram_35;
output reg      [7:0] iram_36;
output reg      [7:0] iram_37;
output reg      [7:0] iram_38;
output reg      [7:0] iram_39;
output reg      [7:0] iram_40;
output reg      [7:0] iram_41;
output reg      [7:0] iram_42;
output reg      [7:0] iram_43;
output reg      [7:0] iram_44;
output reg      [7:0] iram_45;
output reg      [7:0] iram_46;
output reg      [7:0] iram_47;
output reg      [7:0] iram_48;
output reg      [7:0] iram_49;
output reg      [7:0] iram_50;
output reg      [7:0] iram_51;
output reg      [7:0] iram_52;
output reg      [7:0] iram_53;
output reg      [7:0] iram_54;
output reg      [7:0] iram_55;
output reg      [7:0] iram_56;
output reg      [7:0] iram_57;
output reg      [7:0] iram_58;
output reg      [7:0] iram_59;
output reg      [7:0] iram_60;
output reg      [7:0] iram_61;
output reg      [7:0] iram_62;
output reg      [7:0] iram_63;
output reg      [7:0] iram_64;
output reg      [7:0] iram_65;
output reg      [7:0] iram_66;
output reg      [7:0] iram_67;
output reg      [7:0] iram_68;
output reg      [7:0] iram_69;
output reg      [7:0] iram_70;
output reg      [7:0] iram_71;
output reg      [7:0] iram_72;
output reg      [7:0] iram_73;
output reg      [7:0] iram_74;
output reg      [7:0] iram_75;
output reg      [7:0] iram_76;
output reg      [7:0] iram_77;
output reg      [7:0] iram_78;
output reg      [7:0] iram_79;
output reg      [7:0] iram_80;
output reg      [7:0] iram_81;
output reg      [7:0] iram_82;
output reg      [7:0] iram_83;
output reg      [7:0] iram_84;
output reg      [7:0] iram_85;
output reg      [7:0] iram_86;
output reg      [7:0] iram_87;
output reg      [7:0] iram_88;
output reg      [7:0] iram_89;
output reg      [7:0] iram_90;
output reg      [7:0] iram_91;
output reg      [7:0] iram_92;
output reg      [7:0] iram_93;
output reg      [7:0] iram_94;
output reg      [7:0] iram_95;
output reg      [7:0] iram_96;
output reg      [7:0] iram_97;
output reg      [7:0] iram_98;
output reg      [7:0] iram_99;
output reg      [7:0] iram_100;
output reg      [7:0] iram_101;
output reg      [7:0] iram_102;
output reg      [7:0] iram_103;
output reg      [7:0] iram_104;
output reg      [7:0] iram_105;
output reg      [7:0] iram_106;
output reg      [7:0] iram_107;
output reg      [7:0] iram_108;
output reg      [7:0] iram_109;
output reg      [7:0] iram_110;
output reg      [7:0] iram_111;
output reg      [7:0] iram_112;
output reg      [7:0] iram_113;
output reg      [7:0] iram_114;
output reg      [7:0] iram_115;
output reg      [7:0] iram_116;
output reg      [7:0] iram_117;
output reg      [7:0] iram_118;
output reg      [7:0] iram_119;
output reg      [7:0] iram_120;
output reg      [7:0] iram_121;
output reg      [7:0] iram_122;
output reg      [7:0] iram_123;
output reg      [7:0] iram_124;
output reg      [7:0] iram_125;
output reg      [7:0] iram_126;
output reg      [7:0] iram_127;
output reg      [7:0] iram_128;
output reg      [7:0] iram_129;
output reg      [7:0] iram_130;
output reg      [7:0] iram_131;
output reg      [7:0] iram_132;
output reg      [7:0] iram_133;
output reg      [7:0] iram_134;
output reg      [7:0] iram_135;
output reg      [7:0] iram_136;
output reg      [7:0] iram_137;
output reg      [7:0] iram_138;
output reg      [7:0] iram_139;
output reg      [7:0] iram_140;
output reg      [7:0] iram_141;
output reg      [7:0] iram_142;
output reg      [7:0] iram_143;
output reg      [7:0] iram_144;
output reg      [7:0] iram_145;
output reg      [7:0] iram_146;
output reg      [7:0] iram_147;
output reg      [7:0] iram_148;
output reg      [7:0] iram_149;
output reg      [7:0] iram_150;
output reg      [7:0] iram_151;
output reg      [7:0] iram_152;
output reg      [7:0] iram_153;
output reg      [7:0] iram_154;
output reg      [7:0] iram_155;
output reg      [7:0] iram_156;
output reg      [7:0] iram_157;
output reg      [7:0] iram_158;
output reg      [7:0] iram_159;
output reg      [7:0] iram_160;
output reg      [7:0] iram_161;
output reg      [7:0] iram_162;
output reg      [7:0] iram_163;
output reg      [7:0] iram_164;
output reg      [7:0] iram_165;
output reg      [7:0] iram_166;
output reg      [7:0] iram_167;
output reg      [7:0] iram_168;
output reg      [7:0] iram_169;
output reg      [7:0] iram_170;
output reg      [7:0] iram_171;
output reg      [7:0] iram_172;
output reg      [7:0] iram_173;
output reg      [7:0] iram_174;
output reg      [7:0] iram_175;
output reg      [7:0] iram_176;
output reg      [7:0] iram_177;
output reg      [7:0] iram_178;
output reg      [7:0] iram_179;
output reg      [7:0] iram_180;
output reg      [7:0] iram_181;
output reg      [7:0] iram_182;
output reg      [7:0] iram_183;
output reg      [7:0] iram_184;
output reg      [7:0] iram_185;
output reg      [7:0] iram_186;
output reg      [7:0] iram_187;
output reg      [7:0] iram_188;
output reg      [7:0] iram_189;
output reg      [7:0] iram_190;
output reg      [7:0] iram_191;
output reg      [7:0] iram_192;
output reg      [7:0] iram_193;
output reg      [7:0] iram_194;
output reg      [7:0] iram_195;
output reg      [7:0] iram_196;
output reg      [7:0] iram_197;
output reg      [7:0] iram_198;
output reg      [7:0] iram_199;
output reg      [7:0] iram_200;
output reg      [7:0] iram_201;
output reg      [7:0] iram_202;
output reg      [7:0] iram_203;
output reg      [7:0] iram_204;
output reg      [7:0] iram_205;
output reg      [7:0] iram_206;
output reg      [7:0] iram_207;
output reg      [7:0] iram_208;
output reg      [7:0] iram_209;
output reg      [7:0] iram_210;
output reg      [7:0] iram_211;
output reg      [7:0] iram_212;
output reg      [7:0] iram_213;
output reg      [7:0] iram_214;
output reg      [7:0] iram_215;
output reg      [7:0] iram_216;
output reg      [7:0] iram_217;
output reg      [7:0] iram_218;
output reg      [7:0] iram_219;
output reg      [7:0] iram_220;
output reg      [7:0] iram_221;
output reg      [7:0] iram_222;
output reg      [7:0] iram_223;
output reg      [7:0] iram_224;
output reg      [7:0] iram_225;
output reg      [7:0] iram_226;
output reg      [7:0] iram_227;
output reg      [7:0] iram_228;
output reg      [7:0] iram_229;
output reg      [7:0] iram_230;
output reg      [7:0] iram_231;
output reg      [7:0] iram_232;
output reg      [7:0] iram_233;
output reg      [7:0] iram_234;
output reg      [7:0] iram_235;
output reg      [7:0] iram_236;
output reg      [7:0] iram_237;
output reg      [7:0] iram_238;
output reg      [7:0] iram_239;
output reg      [7:0] iram_240;
output reg      [7:0] iram_241;
output reg      [7:0] iram_242;
output reg      [7:0] iram_243;
output reg      [7:0] iram_244;
output reg      [7:0] iram_245;
output reg      [7:0] iram_246;
output reg      [7:0] iram_247;
output reg      [7:0] iram_248;
output reg      [7:0] iram_249;
output reg      [7:0] iram_250;
output reg      [7:0] iram_251;
output reg      [7:0] iram_252;
output reg      [7:0] iram_253;
output reg      [7:0] iram_254;
output reg      [7:0] iram_255;
wire     [19:0] __ILA_DATAPATH_acc_decode__;
wire            __ILA_DATAPATH_decode_of_alu_add__;
wire            __ILA_DATAPATH_decode_of_alu_and__;
wire            __ILA_DATAPATH_decode_of_alu_da__;
wire            __ILA_DATAPATH_decode_of_alu_div__;
wire            __ILA_DATAPATH_decode_of_alu_inc__;
wire            __ILA_DATAPATH_decode_of_alu_mul__;
wire            __ILA_DATAPATH_decode_of_alu_not__;
wire            __ILA_DATAPATH_decode_of_alu_or__;
wire            __ILA_DATAPATH_decode_of_alu_rl__;
wire            __ILA_DATAPATH_decode_of_alu_rlc__;
wire            __ILA_DATAPATH_decode_of_alu_rr__;
wire            __ILA_DATAPATH_decode_of_alu_rrc__;
wire            __ILA_DATAPATH_decode_of_alu_sub__;
wire            __ILA_DATAPATH_decode_of_alu_xch__;
wire            __ILA_DATAPATH_decode_of_alu_xor__;
wire            __ILA_DATAPATH_decode_of_no_wr__;
wire            __ILA_DATAPATH_decode_of_read_data__;
wire            __ILA_DATAPATH_decode_of_wr_ram__;
wire            __ILA_DATAPATH_decode_of_wr_sfr__;
wire            __ILA_DATAPATH_decode_of_wr_sfr_ram__;
wire     [19:0] __ILA_DATAPATH_grant__;
wire            __ILA_DATAPATH_valid__;
wire      [3:0] alu_op;
wire            bit_addr;
wire            bit_in;
wire     [15:0] bv_16_1_n4830;
wire            bv_1_0_n53;
wire            bv_1_1_n34;
wire      [1:0] bv_2_0_n4771;
wire      [1:0] bv_2_1_n3501;
wire      [1:0] bv_2_2_n3505;
wire      [1:0] bv_2_3_n3495;
wire      [2:0] bv_3_0_n46;
wire      [2:0] bv_3_1_n3667;
wire      [2:0] bv_3_2_n3664;
wire      [2:0] bv_3_3_n3517;
wire      [2:0] bv_3_4_n3659;
wire      [2:0] bv_3_5_n3656;
wire      [2:0] bv_3_6_n3653;
wire      [2:0] bv_3_7_n3557;
wire      [3:0] bv_4_0_n30;
wire      [3:0] bv_4_10_n16;
wire      [3:0] bv_4_11_n18;
wire      [3:0] bv_4_12_n20;
wire      [3:0] bv_4_13_n22;
wire      [3:0] bv_4_14_n2;
wire      [3:0] bv_4_15_n24;
wire      [3:0] bv_4_1_n28;
wire      [3:0] bv_4_2_n12;
wire      [3:0] bv_4_3_n8;
wire      [3:0] bv_4_4_n10;
wire      [3:0] bv_4_5_n6;
wire      [3:0] bv_4_6_n4;
wire      [3:0] bv_4_7_n0;
wire      [3:0] bv_4_8_n26;
wire      [3:0] bv_4_9_n14;
wire      [4:0] bv_5_16_n3727;
wire      [4:0] bv_5_18_n3751;
wire      [4:0] bv_5_20_n3775;
wire      [4:0] bv_5_21_n3871;
wire      [4:0] bv_5_22_n3799;
wire      [4:0] bv_5_23_n3847;
wire      [4:0] bv_5_26_n3701;
wire      [4:0] bv_5_28_n3647;
wire      [4:0] bv_5_30_n3823;
wire      [4:0] bv_5_6_n4912;
wire      [6:0] bv_7_0_n3520;
wire      [7:0] bv_8_0_n69;
wire      [7:0] bv_8_100_n269;
wire      [7:0] bv_8_101_n271;
wire      [7:0] bv_8_102_n273;
wire      [7:0] bv_8_103_n275;
wire      [7:0] bv_8_104_n277;
wire      [7:0] bv_8_105_n279;
wire      [7:0] bv_8_106_n281;
wire      [7:0] bv_8_107_n283;
wire      [7:0] bv_8_108_n285;
wire      [7:0] bv_8_109_n287;
wire      [7:0] bv_8_10_n89;
wire      [7:0] bv_8_110_n289;
wire      [7:0] bv_8_111_n291;
wire      [7:0] bv_8_112_n293;
wire      [7:0] bv_8_113_n295;
wire      [7:0] bv_8_114_n297;
wire      [7:0] bv_8_115_n299;
wire      [7:0] bv_8_116_n301;
wire      [7:0] bv_8_117_n303;
wire      [7:0] bv_8_118_n305;
wire      [7:0] bv_8_119_n307;
wire      [7:0] bv_8_11_n91;
wire      [7:0] bv_8_120_n309;
wire      [7:0] bv_8_121_n311;
wire      [7:0] bv_8_122_n313;
wire      [7:0] bv_8_123_n315;
wire      [7:0] bv_8_124_n317;
wire      [7:0] bv_8_125_n319;
wire      [7:0] bv_8_126_n321;
wire      [7:0] bv_8_127_n323;
wire      [7:0] bv_8_128_n325;
wire      [7:0] bv_8_129_n327;
wire      [7:0] bv_8_12_n93;
wire      [7:0] bv_8_130_n329;
wire      [7:0] bv_8_131_n331;
wire      [7:0] bv_8_132_n333;
wire      [7:0] bv_8_133_n335;
wire      [7:0] bv_8_134_n337;
wire      [7:0] bv_8_135_n339;
wire      [7:0] bv_8_136_n341;
wire      [7:0] bv_8_137_n343;
wire      [7:0] bv_8_138_n345;
wire      [7:0] bv_8_139_n347;
wire      [7:0] bv_8_13_n95;
wire      [7:0] bv_8_140_n349;
wire      [7:0] bv_8_141_n351;
wire      [7:0] bv_8_142_n353;
wire      [7:0] bv_8_143_n355;
wire      [7:0] bv_8_144_n357;
wire      [7:0] bv_8_145_n359;
wire      [7:0] bv_8_146_n361;
wire      [7:0] bv_8_147_n363;
wire      [7:0] bv_8_148_n365;
wire      [7:0] bv_8_149_n367;
wire      [7:0] bv_8_14_n97;
wire      [7:0] bv_8_150_n369;
wire      [7:0] bv_8_151_n371;
wire      [7:0] bv_8_152_n373;
wire      [7:0] bv_8_153_n375;
wire      [7:0] bv_8_154_n377;
wire      [7:0] bv_8_155_n379;
wire      [7:0] bv_8_156_n381;
wire      [7:0] bv_8_157_n383;
wire      [7:0] bv_8_158_n385;
wire      [7:0] bv_8_159_n387;
wire      [7:0] bv_8_15_n99;
wire      [7:0] bv_8_160_n389;
wire      [7:0] bv_8_161_n391;
wire      [7:0] bv_8_162_n393;
wire      [7:0] bv_8_163_n395;
wire      [7:0] bv_8_164_n397;
wire      [7:0] bv_8_165_n399;
wire      [7:0] bv_8_166_n401;
wire      [7:0] bv_8_167_n403;
wire      [7:0] bv_8_168_n405;
wire      [7:0] bv_8_169_n407;
wire      [7:0] bv_8_16_n101;
wire      [7:0] bv_8_170_n409;
wire      [7:0] bv_8_171_n411;
wire      [7:0] bv_8_172_n413;
wire      [7:0] bv_8_173_n415;
wire      [7:0] bv_8_174_n417;
wire      [7:0] bv_8_175_n419;
wire      [7:0] bv_8_176_n421;
wire      [7:0] bv_8_177_n423;
wire      [7:0] bv_8_178_n425;
wire      [7:0] bv_8_179_n427;
wire      [7:0] bv_8_17_n103;
wire      [7:0] bv_8_180_n429;
wire      [7:0] bv_8_181_n431;
wire      [7:0] bv_8_182_n433;
wire      [7:0] bv_8_183_n435;
wire      [7:0] bv_8_184_n437;
wire      [7:0] bv_8_185_n439;
wire      [7:0] bv_8_186_n441;
wire      [7:0] bv_8_187_n443;
wire      [7:0] bv_8_188_n445;
wire      [7:0] bv_8_189_n447;
wire      [7:0] bv_8_18_n105;
wire      [7:0] bv_8_190_n449;
wire      [7:0] bv_8_191_n451;
wire      [7:0] bv_8_192_n453;
wire      [7:0] bv_8_193_n455;
wire      [7:0] bv_8_194_n457;
wire      [7:0] bv_8_195_n459;
wire      [7:0] bv_8_196_n461;
wire      [7:0] bv_8_197_n463;
wire      [7:0] bv_8_198_n465;
wire      [7:0] bv_8_199_n467;
wire      [7:0] bv_8_19_n107;
wire      [7:0] bv_8_1_n71;
wire      [7:0] bv_8_200_n469;
wire      [7:0] bv_8_201_n471;
wire      [7:0] bv_8_202_n473;
wire      [7:0] bv_8_203_n475;
wire      [7:0] bv_8_204_n477;
wire      [7:0] bv_8_205_n479;
wire      [7:0] bv_8_206_n481;
wire      [7:0] bv_8_207_n483;
wire      [7:0] bv_8_208_n485;
wire      [7:0] bv_8_209_n487;
wire      [7:0] bv_8_20_n109;
wire      [7:0] bv_8_210_n489;
wire      [7:0] bv_8_211_n491;
wire      [7:0] bv_8_212_n493;
wire      [7:0] bv_8_213_n495;
wire      [7:0] bv_8_214_n497;
wire      [7:0] bv_8_215_n499;
wire      [7:0] bv_8_216_n501;
wire      [7:0] bv_8_217_n503;
wire      [7:0] bv_8_218_n505;
wire      [7:0] bv_8_219_n507;
wire      [7:0] bv_8_21_n111;
wire      [7:0] bv_8_220_n509;
wire      [7:0] bv_8_221_n511;
wire      [7:0] bv_8_222_n513;
wire      [7:0] bv_8_223_n515;
wire      [7:0] bv_8_224_n517;
wire      [7:0] bv_8_225_n519;
wire      [7:0] bv_8_226_n521;
wire      [7:0] bv_8_227_n523;
wire      [7:0] bv_8_228_n525;
wire      [7:0] bv_8_229_n527;
wire      [7:0] bv_8_22_n113;
wire      [7:0] bv_8_230_n529;
wire      [7:0] bv_8_231_n531;
wire      [7:0] bv_8_232_n533;
wire      [7:0] bv_8_233_n535;
wire      [7:0] bv_8_234_n537;
wire      [7:0] bv_8_235_n539;
wire      [7:0] bv_8_236_n541;
wire      [7:0] bv_8_237_n543;
wire      [7:0] bv_8_238_n545;
wire      [7:0] bv_8_239_n547;
wire      [7:0] bv_8_23_n115;
wire      [7:0] bv_8_240_n549;
wire      [7:0] bv_8_241_n551;
wire      [7:0] bv_8_242_n553;
wire      [7:0] bv_8_243_n555;
wire      [7:0] bv_8_244_n557;
wire      [7:0] bv_8_245_n559;
wire      [7:0] bv_8_246_n561;
wire      [7:0] bv_8_247_n563;
wire      [7:0] bv_8_248_n565;
wire      [7:0] bv_8_249_n567;
wire      [7:0] bv_8_24_n117;
wire      [7:0] bv_8_250_n569;
wire      [7:0] bv_8_251_n571;
wire      [7:0] bv_8_252_n573;
wire      [7:0] bv_8_253_n575;
wire      [7:0] bv_8_254_n577;
wire      [7:0] bv_8_255_n29279;
wire      [7:0] bv_8_25_n119;
wire      [7:0] bv_8_26_n121;
wire      [7:0] bv_8_27_n123;
wire      [7:0] bv_8_28_n125;
wire      [7:0] bv_8_29_n127;
wire      [7:0] bv_8_2_n73;
wire      [7:0] bv_8_30_n129;
wire      [7:0] bv_8_31_n131;
wire      [7:0] bv_8_32_n133;
wire      [7:0] bv_8_33_n135;
wire      [7:0] bv_8_34_n137;
wire      [7:0] bv_8_35_n139;
wire      [7:0] bv_8_36_n141;
wire      [7:0] bv_8_37_n143;
wire      [7:0] bv_8_38_n145;
wire      [7:0] bv_8_39_n147;
wire      [7:0] bv_8_3_n75;
wire      [7:0] bv_8_40_n149;
wire      [7:0] bv_8_41_n151;
wire      [7:0] bv_8_42_n153;
wire      [7:0] bv_8_43_n155;
wire      [7:0] bv_8_44_n157;
wire      [7:0] bv_8_45_n159;
wire      [7:0] bv_8_46_n161;
wire      [7:0] bv_8_47_n163;
wire      [7:0] bv_8_48_n165;
wire      [7:0] bv_8_49_n167;
wire      [7:0] bv_8_4_n77;
wire      [7:0] bv_8_50_n169;
wire      [7:0] bv_8_51_n171;
wire      [7:0] bv_8_52_n173;
wire      [7:0] bv_8_53_n175;
wire      [7:0] bv_8_54_n177;
wire      [7:0] bv_8_55_n179;
wire      [7:0] bv_8_56_n181;
wire      [7:0] bv_8_57_n183;
wire      [7:0] bv_8_58_n185;
wire      [7:0] bv_8_59_n187;
wire      [7:0] bv_8_5_n79;
wire      [7:0] bv_8_60_n189;
wire      [7:0] bv_8_61_n191;
wire      [7:0] bv_8_62_n193;
wire      [7:0] bv_8_63_n195;
wire      [7:0] bv_8_64_n197;
wire      [7:0] bv_8_65_n199;
wire      [7:0] bv_8_66_n201;
wire      [7:0] bv_8_67_n203;
wire      [7:0] bv_8_68_n205;
wire      [7:0] bv_8_69_n207;
wire      [7:0] bv_8_6_n81;
wire      [7:0] bv_8_70_n209;
wire      [7:0] bv_8_71_n211;
wire      [7:0] bv_8_72_n213;
wire      [7:0] bv_8_73_n215;
wire      [7:0] bv_8_74_n217;
wire      [7:0] bv_8_75_n219;
wire      [7:0] bv_8_76_n221;
wire      [7:0] bv_8_77_n223;
wire      [7:0] bv_8_78_n225;
wire      [7:0] bv_8_79_n227;
wire      [7:0] bv_8_7_n83;
wire      [7:0] bv_8_80_n229;
wire      [7:0] bv_8_81_n231;
wire      [7:0] bv_8_82_n233;
wire      [7:0] bv_8_83_n235;
wire      [7:0] bv_8_84_n237;
wire      [7:0] bv_8_85_n239;
wire      [7:0] bv_8_86_n241;
wire      [7:0] bv_8_87_n243;
wire      [7:0] bv_8_88_n245;
wire      [7:0] bv_8_89_n247;
wire      [7:0] bv_8_8_n85;
wire      [7:0] bv_8_90_n249;
wire      [7:0] bv_8_91_n251;
wire      [7:0] bv_8_92_n253;
wire      [7:0] bv_8_93_n255;
wire      [7:0] bv_8_94_n257;
wire      [7:0] bv_8_95_n259;
wire      [7:0] bv_8_96_n261;
wire      [7:0] bv_8_97_n263;
wire      [7:0] bv_8_98_n265;
wire      [7:0] bv_8_99_n267;
wire      [7:0] bv_8_9_n87;
wire            clk;
wire      [1:0] cy_sel;
wire            n1;
wire            n100;
wire            n1000;
wire            n10000;
wire            n10001;
wire            n10002;
wire            n10003;
wire      [7:0] n10004;
wire            n10005;
wire            n10006;
wire            n10007;
wire            n10008;
wire            n10009;
wire            n1001;
wire      [7:0] n10010;
wire            n10011;
wire            n10012;
wire            n10013;
wire            n10014;
wire            n10015;
wire      [7:0] n10016;
wire            n10017;
wire            n10018;
wire            n10019;
wire            n1002;
wire            n10020;
wire            n10021;
wire      [7:0] n10022;
wire            n10023;
wire            n10024;
wire            n10025;
wire            n10026;
wire            n10027;
wire      [7:0] n10028;
wire            n10029;
wire            n1003;
wire            n10030;
wire            n10031;
wire            n10032;
wire            n10033;
wire      [7:0] n10034;
wire            n10035;
wire            n10036;
wire            n10037;
wire            n10038;
wire            n10039;
wire            n1004;
wire      [7:0] n10040;
wire            n10041;
wire            n10042;
wire            n10043;
wire            n10044;
wire            n10045;
wire      [7:0] n10046;
wire            n10047;
wire            n10048;
wire            n10049;
wire            n1005;
wire            n10050;
wire            n10051;
wire      [7:0] n10052;
wire            n10053;
wire            n10054;
wire            n10055;
wire            n10056;
wire            n10057;
wire      [7:0] n10058;
wire            n10059;
wire            n1006;
wire            n10060;
wire            n10061;
wire            n10062;
wire            n10063;
wire      [7:0] n10064;
wire            n10065;
wire            n10066;
wire            n10067;
wire            n10068;
wire            n10069;
wire            n1007;
wire      [7:0] n10070;
wire            n10071;
wire            n10072;
wire            n10073;
wire            n10074;
wire            n10075;
wire      [7:0] n10076;
wire            n10077;
wire            n10078;
wire            n10079;
wire            n1008;
wire            n10080;
wire            n10081;
wire      [7:0] n10082;
wire            n10083;
wire            n10084;
wire            n10085;
wire            n10086;
wire            n10087;
wire      [7:0] n10088;
wire            n10089;
wire            n1009;
wire            n10090;
wire            n10091;
wire            n10092;
wire            n10093;
wire      [7:0] n10094;
wire            n10095;
wire            n10096;
wire            n10097;
wire            n10098;
wire            n10099;
wire            n1010;
wire      [7:0] n10100;
wire            n10101;
wire            n10102;
wire            n10103;
wire            n10104;
wire            n10105;
wire      [7:0] n10106;
wire            n10107;
wire            n10108;
wire            n10109;
wire            n1011;
wire            n10110;
wire            n10111;
wire      [7:0] n10112;
wire            n10113;
wire            n10114;
wire            n10115;
wire            n10116;
wire            n10117;
wire      [7:0] n10118;
wire            n10119;
wire            n1012;
wire            n10120;
wire            n10121;
wire            n10122;
wire            n10123;
wire      [7:0] n10124;
wire            n10125;
wire            n10126;
wire            n10127;
wire            n10128;
wire            n10129;
wire            n1013;
wire      [7:0] n10130;
wire            n10131;
wire            n10132;
wire            n10133;
wire            n10134;
wire            n10135;
wire      [7:0] n10136;
wire            n10137;
wire            n10138;
wire            n10139;
wire            n1014;
wire            n10140;
wire            n10141;
wire      [7:0] n10142;
wire            n10143;
wire            n10144;
wire            n10145;
wire            n10146;
wire            n10147;
wire      [7:0] n10148;
wire            n10149;
wire            n1015;
wire            n10150;
wire            n10151;
wire            n10152;
wire            n10153;
wire      [7:0] n10154;
wire            n10155;
wire            n10156;
wire            n10157;
wire            n10158;
wire            n10159;
wire            n1016;
wire      [7:0] n10160;
wire            n10161;
wire            n10162;
wire            n10163;
wire            n10164;
wire            n10165;
wire      [7:0] n10166;
wire            n10167;
wire            n10168;
wire            n10169;
wire            n1017;
wire            n10170;
wire            n10171;
wire      [7:0] n10172;
wire            n10173;
wire            n10174;
wire            n10175;
wire            n10176;
wire            n10177;
wire      [7:0] n10178;
wire            n10179;
wire            n1018;
wire            n10180;
wire            n10181;
wire            n10182;
wire            n10183;
wire      [7:0] n10184;
wire            n10185;
wire            n10186;
wire            n10187;
wire            n10188;
wire            n10189;
wire            n1019;
wire      [7:0] n10190;
wire            n10191;
wire            n10192;
wire            n10193;
wire            n10194;
wire            n10195;
wire      [7:0] n10196;
wire            n10197;
wire            n10198;
wire            n10199;
wire            n102;
wire            n1020;
wire            n10200;
wire            n10201;
wire      [7:0] n10202;
wire            n10203;
wire            n10204;
wire            n10205;
wire            n10206;
wire            n10207;
wire      [7:0] n10208;
wire            n10209;
wire            n1021;
wire            n10210;
wire            n10211;
wire            n10212;
wire            n10213;
wire      [7:0] n10214;
wire            n10215;
wire            n10216;
wire            n10217;
wire            n10218;
wire            n10219;
wire            n1022;
wire      [7:0] n10220;
wire            n10221;
wire            n10222;
wire            n10223;
wire            n10224;
wire            n10225;
wire      [7:0] n10226;
wire            n10227;
wire            n10228;
wire            n10229;
wire            n1023;
wire            n10230;
wire            n10231;
wire      [7:0] n10232;
wire            n10233;
wire            n10234;
wire            n10235;
wire            n10236;
wire            n10237;
wire      [7:0] n10238;
wire            n10239;
wire            n1024;
wire            n10240;
wire            n10241;
wire            n10242;
wire            n10243;
wire      [7:0] n10244;
wire            n10245;
wire            n10246;
wire            n10247;
wire            n10248;
wire            n10249;
wire            n1025;
wire      [7:0] n10250;
wire            n10251;
wire            n10252;
wire            n10253;
wire            n10254;
wire            n10255;
wire      [7:0] n10256;
wire            n10257;
wire            n10258;
wire            n10259;
wire            n1026;
wire            n10260;
wire            n10261;
wire      [7:0] n10262;
wire            n10263;
wire            n10264;
wire            n10265;
wire            n10266;
wire            n10267;
wire      [7:0] n10268;
wire            n10269;
wire            n1027;
wire            n10270;
wire            n10271;
wire            n10272;
wire            n10273;
wire      [7:0] n10274;
wire            n10275;
wire            n10276;
wire            n10277;
wire            n10278;
wire            n10279;
wire            n1028;
wire      [7:0] n10280;
wire            n10281;
wire            n10282;
wire            n10283;
wire            n10284;
wire            n10285;
wire      [7:0] n10286;
wire            n10287;
wire            n10288;
wire            n10289;
wire            n1029;
wire            n10290;
wire            n10291;
wire      [7:0] n10292;
wire            n10293;
wire            n10294;
wire            n10295;
wire            n10296;
wire            n10297;
wire      [7:0] n10298;
wire            n10299;
wire            n1030;
wire            n10300;
wire            n10301;
wire            n10302;
wire            n10303;
wire      [7:0] n10304;
wire            n10305;
wire            n10306;
wire            n10307;
wire            n10308;
wire            n10309;
wire            n1031;
wire      [7:0] n10310;
wire            n10311;
wire            n10312;
wire            n10313;
wire            n10314;
wire            n10315;
wire      [7:0] n10316;
wire            n10317;
wire            n10318;
wire            n10319;
wire            n1032;
wire            n10320;
wire            n10321;
wire      [7:0] n10322;
wire            n10323;
wire            n10324;
wire            n10325;
wire            n10326;
wire            n10327;
wire      [7:0] n10328;
wire            n10329;
wire            n1033;
wire            n10330;
wire            n10331;
wire            n10332;
wire            n10333;
wire      [7:0] n10334;
wire            n10335;
wire            n10336;
wire            n10337;
wire            n10338;
wire            n10339;
wire            n1034;
wire      [7:0] n10340;
wire            n10341;
wire            n10342;
wire            n10343;
wire            n10344;
wire            n10345;
wire      [7:0] n10346;
wire            n10347;
wire            n10348;
wire            n10349;
wire            n1035;
wire            n10350;
wire            n10351;
wire      [7:0] n10352;
wire            n10353;
wire            n10354;
wire            n10355;
wire            n10356;
wire            n10357;
wire      [7:0] n10358;
wire            n10359;
wire            n1036;
wire            n10360;
wire            n10361;
wire            n10362;
wire            n10363;
wire      [7:0] n10364;
wire            n10365;
wire            n10366;
wire            n10367;
wire            n10368;
wire            n10369;
wire            n1037;
wire      [7:0] n10370;
wire            n10371;
wire            n10372;
wire            n10373;
wire            n10374;
wire            n10375;
wire      [7:0] n10376;
wire            n10377;
wire            n10378;
wire            n10379;
wire            n1038;
wire            n10380;
wire            n10381;
wire      [7:0] n10382;
wire            n10383;
wire            n10384;
wire            n10385;
wire            n10386;
wire            n10387;
wire      [7:0] n10388;
wire            n10389;
wire            n1039;
wire            n10390;
wire            n10391;
wire            n10392;
wire            n10393;
wire      [7:0] n10394;
wire            n10395;
wire            n10396;
wire            n10397;
wire            n10398;
wire            n10399;
wire            n104;
wire            n1040;
wire      [7:0] n10400;
wire            n10401;
wire            n10402;
wire            n10403;
wire            n10404;
wire            n10405;
wire      [7:0] n10406;
wire            n10407;
wire            n10408;
wire            n10409;
wire            n1041;
wire            n10410;
wire            n10411;
wire      [7:0] n10412;
wire            n10413;
wire            n10414;
wire            n10415;
wire            n10416;
wire            n10417;
wire      [7:0] n10418;
wire            n10419;
wire            n1042;
wire            n10420;
wire            n10421;
wire            n10422;
wire            n10423;
wire      [7:0] n10424;
wire            n10425;
wire            n10426;
wire            n10427;
wire            n10428;
wire            n10429;
wire            n1043;
wire      [7:0] n10430;
wire            n10431;
wire            n10432;
wire            n10433;
wire            n10434;
wire            n10435;
wire      [7:0] n10436;
wire            n10437;
wire            n10438;
wire            n10439;
wire            n1044;
wire            n10440;
wire            n10441;
wire      [7:0] n10442;
wire            n10443;
wire            n10444;
wire            n10445;
wire            n10446;
wire            n10447;
wire      [7:0] n10448;
wire            n10449;
wire            n1045;
wire            n10450;
wire            n10451;
wire            n10452;
wire            n10453;
wire      [7:0] n10454;
wire            n10455;
wire            n10456;
wire            n10457;
wire            n10458;
wire            n10459;
wire            n1046;
wire      [7:0] n10460;
wire            n10461;
wire            n10462;
wire            n10463;
wire            n10464;
wire            n10465;
wire      [7:0] n10466;
wire            n10467;
wire            n10468;
wire            n10469;
wire            n1047;
wire            n10470;
wire            n10471;
wire      [7:0] n10472;
wire            n10473;
wire            n10474;
wire            n10475;
wire            n10476;
wire            n10477;
wire      [7:0] n10478;
wire            n10479;
wire            n1048;
wire            n10480;
wire            n10481;
wire            n10482;
wire            n10483;
wire      [7:0] n10484;
wire            n10485;
wire            n10486;
wire            n10487;
wire            n10488;
wire            n10489;
wire            n1049;
wire      [7:0] n10490;
wire            n10491;
wire            n10492;
wire            n10493;
wire            n10494;
wire            n10495;
wire      [7:0] n10496;
wire            n10497;
wire            n10498;
wire            n10499;
wire            n1050;
wire            n10500;
wire            n10501;
wire      [7:0] n10502;
wire            n10503;
wire            n10504;
wire            n10505;
wire            n10506;
wire            n10507;
wire      [7:0] n10508;
wire            n10509;
wire            n1051;
wire            n10510;
wire            n10511;
wire            n10512;
wire            n10513;
wire      [7:0] n10514;
wire            n10515;
wire            n10516;
wire            n10517;
wire            n10518;
wire            n10519;
wire            n1052;
wire      [7:0] n10520;
wire            n10521;
wire            n10522;
wire            n10523;
wire            n10524;
wire            n10525;
wire      [7:0] n10526;
wire            n10527;
wire            n10528;
wire            n10529;
wire            n1053;
wire            n10530;
wire            n10531;
wire      [7:0] n10532;
wire            n10533;
wire            n10534;
wire            n10535;
wire            n10536;
wire            n10537;
wire      [7:0] n10538;
wire            n10539;
wire            n1054;
wire            n10540;
wire            n10541;
wire            n10542;
wire            n10543;
wire      [7:0] n10544;
wire            n10545;
wire            n10546;
wire            n10547;
wire            n10548;
wire            n10549;
wire            n1055;
wire      [7:0] n10550;
wire            n10551;
wire            n10552;
wire            n10553;
wire            n10554;
wire            n10555;
wire      [7:0] n10556;
wire            n10557;
wire            n10558;
wire            n10559;
wire            n1056;
wire            n10560;
wire            n10561;
wire      [7:0] n10562;
wire            n10563;
wire            n10564;
wire            n10565;
wire            n10566;
wire            n10567;
wire      [7:0] n10568;
wire            n10569;
wire            n1057;
wire            n10570;
wire            n10571;
wire            n10572;
wire            n10573;
wire      [7:0] n10574;
wire            n10575;
wire            n10576;
wire            n10577;
wire            n10578;
wire            n10579;
wire            n1058;
wire      [7:0] n10580;
wire            n10581;
wire            n10582;
wire            n10583;
wire            n10584;
wire            n10585;
wire      [7:0] n10586;
wire            n10587;
wire            n10588;
wire            n10589;
wire            n1059;
wire            n10590;
wire            n10591;
wire      [7:0] n10592;
wire            n10593;
wire            n10594;
wire            n10595;
wire            n10596;
wire            n10597;
wire      [7:0] n10598;
wire            n10599;
wire            n106;
wire            n1060;
wire            n10600;
wire            n10601;
wire            n10602;
wire            n10603;
wire      [7:0] n10604;
wire            n10605;
wire            n10606;
wire            n10607;
wire            n10608;
wire            n10609;
wire            n1061;
wire      [7:0] n10610;
wire            n10611;
wire            n10612;
wire            n10613;
wire            n10614;
wire            n10615;
wire      [7:0] n10616;
wire            n10617;
wire            n10618;
wire            n10619;
wire            n1062;
wire            n10620;
wire            n10621;
wire      [7:0] n10622;
wire            n10623;
wire            n10624;
wire            n10625;
wire            n10626;
wire            n10627;
wire      [7:0] n10628;
wire            n10629;
wire            n1063;
wire            n10630;
wire            n10631;
wire            n10632;
wire            n10633;
wire      [7:0] n10634;
wire            n10635;
wire            n10636;
wire            n10637;
wire            n10638;
wire            n10639;
wire            n1064;
wire      [7:0] n10640;
wire            n10641;
wire            n10642;
wire            n10643;
wire            n10644;
wire            n10645;
wire      [7:0] n10646;
wire            n10647;
wire            n10648;
wire            n10649;
wire            n1065;
wire            n10650;
wire            n10651;
wire      [7:0] n10652;
wire            n10653;
wire            n10654;
wire            n10655;
wire            n10656;
wire            n10657;
wire      [7:0] n10658;
wire            n10659;
wire            n1066;
wire            n10660;
wire            n10661;
wire            n10662;
wire            n10663;
wire      [7:0] n10664;
wire            n10665;
wire            n10666;
wire            n10667;
wire            n10668;
wire            n10669;
wire            n1067;
wire      [7:0] n10670;
wire            n10671;
wire            n10672;
wire            n10673;
wire            n10674;
wire            n10675;
wire      [7:0] n10676;
wire            n10677;
wire            n10678;
wire            n10679;
wire            n1068;
wire            n10680;
wire            n10681;
wire      [7:0] n10682;
wire            n10683;
wire            n10684;
wire            n10685;
wire            n10686;
wire            n10687;
wire      [7:0] n10688;
wire            n10689;
wire            n1069;
wire            n10690;
wire            n10691;
wire            n10692;
wire            n10693;
wire      [7:0] n10694;
wire            n10695;
wire            n10696;
wire            n10697;
wire            n10698;
wire            n10699;
wire            n1070;
wire      [7:0] n10700;
wire            n10701;
wire            n10702;
wire            n10703;
wire            n10704;
wire            n10705;
wire      [7:0] n10706;
wire            n10707;
wire            n10708;
wire            n10709;
wire            n1071;
wire            n10710;
wire            n10711;
wire      [7:0] n10712;
wire            n10713;
wire            n10714;
wire            n10715;
wire            n10716;
wire            n10717;
wire      [7:0] n10718;
wire            n10719;
wire            n1072;
wire            n10720;
wire            n10721;
wire            n10722;
wire            n10723;
wire      [7:0] n10724;
wire            n10725;
wire            n10726;
wire            n10727;
wire            n10728;
wire            n10729;
wire            n1073;
wire      [7:0] n10730;
wire            n10731;
wire            n10732;
wire            n10733;
wire            n10734;
wire            n10735;
wire      [7:0] n10736;
wire            n10737;
wire            n10738;
wire            n10739;
wire            n1074;
wire            n10740;
wire            n10741;
wire      [7:0] n10742;
wire            n10743;
wire            n10744;
wire            n10745;
wire            n10746;
wire            n10747;
wire      [7:0] n10748;
wire            n10749;
wire            n1075;
wire            n10750;
wire            n10751;
wire            n10752;
wire            n10753;
wire      [7:0] n10754;
wire            n10755;
wire            n10756;
wire            n10757;
wire            n10758;
wire            n10759;
wire            n1076;
wire      [7:0] n10760;
wire            n10761;
wire            n10762;
wire            n10763;
wire            n10764;
wire            n10765;
wire      [7:0] n10766;
wire            n10767;
wire            n10768;
wire            n10769;
wire            n1077;
wire            n10770;
wire            n10771;
wire      [7:0] n10772;
wire            n10773;
wire            n10774;
wire            n10775;
wire            n10776;
wire            n10777;
wire      [7:0] n10778;
wire            n10779;
wire            n1078;
wire            n10780;
wire            n10781;
wire            n10782;
wire            n10783;
wire      [7:0] n10784;
wire            n10785;
wire            n10786;
wire            n10787;
wire            n10788;
wire            n10789;
wire            n1079;
wire      [7:0] n10790;
wire            n10791;
wire            n10792;
wire            n10793;
wire            n10794;
wire            n10795;
wire      [7:0] n10796;
wire            n10797;
wire            n10798;
wire            n10799;
wire            n108;
wire            n1080;
wire            n10800;
wire            n10801;
wire      [7:0] n10802;
wire            n10803;
wire            n10804;
wire            n10805;
wire            n10806;
wire            n10807;
wire      [7:0] n10808;
wire            n10809;
wire            n1081;
wire            n10810;
wire            n10811;
wire            n10812;
wire            n10813;
wire      [7:0] n10814;
wire            n10815;
wire            n10816;
wire            n10817;
wire            n10818;
wire            n10819;
wire            n1082;
wire      [7:0] n10820;
wire            n10821;
wire            n10822;
wire            n10823;
wire            n10824;
wire            n10825;
wire      [7:0] n10826;
wire            n10827;
wire            n10828;
wire            n10829;
wire            n1083;
wire            n10830;
wire            n10831;
wire      [7:0] n10832;
wire            n10833;
wire            n10834;
wire            n10835;
wire            n10836;
wire            n10837;
wire      [7:0] n10838;
wire            n10839;
wire            n1084;
wire            n10840;
wire            n10841;
wire            n10842;
wire            n10843;
wire      [7:0] n10844;
wire            n10845;
wire            n10846;
wire            n10847;
wire            n10848;
wire            n10849;
wire            n1085;
wire      [7:0] n10850;
wire            n10851;
wire            n10852;
wire            n10853;
wire            n10854;
wire            n10855;
wire      [7:0] n10856;
wire            n10857;
wire            n10858;
wire            n10859;
wire            n1086;
wire            n10860;
wire            n10861;
wire      [7:0] n10862;
wire            n10863;
wire            n10864;
wire            n10865;
wire            n10866;
wire            n10867;
wire      [7:0] n10868;
wire            n10869;
wire            n1087;
wire            n10870;
wire            n10871;
wire            n10872;
wire            n10873;
wire      [7:0] n10874;
wire            n10875;
wire            n10876;
wire            n10877;
wire            n10878;
wire            n10879;
wire            n1088;
wire      [7:0] n10880;
wire            n10881;
wire            n10882;
wire            n10883;
wire            n10884;
wire            n10885;
wire      [7:0] n10886;
wire            n10887;
wire            n10888;
wire            n10889;
wire      [7:0] n1089;
wire            n10890;
wire            n10891;
wire      [7:0] n10892;
wire            n10893;
wire            n10894;
wire            n10895;
wire            n10896;
wire            n10897;
wire      [7:0] n10898;
wire            n10899;
wire      [7:0] n1090;
wire            n10900;
wire            n10901;
wire            n10902;
wire            n10903;
wire      [7:0] n10904;
wire            n10905;
wire            n10906;
wire            n10907;
wire            n10908;
wire            n10909;
wire      [7:0] n1091;
wire      [7:0] n10910;
wire            n10911;
wire            n10912;
wire            n10913;
wire            n10914;
wire            n10915;
wire      [7:0] n10916;
wire            n10917;
wire            n10918;
wire            n10919;
wire      [7:0] n1092;
wire            n10920;
wire            n10921;
wire      [7:0] n10922;
wire            n10923;
wire            n10924;
wire            n10925;
wire            n10926;
wire            n10927;
wire      [7:0] n10928;
wire            n10929;
wire      [7:0] n1093;
wire            n10930;
wire            n10931;
wire            n10932;
wire            n10933;
wire      [7:0] n10934;
wire            n10935;
wire            n10936;
wire            n10937;
wire            n10938;
wire            n10939;
wire      [7:0] n1094;
wire      [7:0] n10940;
wire            n10941;
wire            n10942;
wire            n10943;
wire            n10944;
wire            n10945;
wire      [7:0] n10946;
wire            n10947;
wire            n10948;
wire            n10949;
wire      [7:0] n1095;
wire            n10950;
wire            n10951;
wire      [7:0] n10952;
wire            n10953;
wire            n10954;
wire            n10955;
wire            n10956;
wire            n10957;
wire      [7:0] n10958;
wire            n10959;
wire      [7:0] n1096;
wire            n10960;
wire            n10961;
wire            n10962;
wire            n10963;
wire      [7:0] n10964;
wire            n10965;
wire            n10966;
wire            n10967;
wire            n10968;
wire            n10969;
wire      [7:0] n1097;
wire      [7:0] n10970;
wire            n10971;
wire            n10972;
wire            n10973;
wire            n10974;
wire            n10975;
wire      [7:0] n10976;
wire            n10977;
wire            n10978;
wire            n10979;
wire      [7:0] n1098;
wire            n10980;
wire            n10981;
wire      [7:0] n10982;
wire            n10983;
wire            n10984;
wire            n10985;
wire            n10986;
wire            n10987;
wire      [7:0] n10988;
wire            n10989;
wire      [7:0] n1099;
wire            n10990;
wire            n10991;
wire            n10992;
wire            n10993;
wire      [7:0] n10994;
wire            n10995;
wire            n10996;
wire            n10997;
wire            n10998;
wire            n10999;
wire            n11;
wire            n110;
wire      [7:0] n1100;
wire      [7:0] n11000;
wire            n11001;
wire            n11002;
wire            n11003;
wire            n11004;
wire            n11005;
wire      [7:0] n11006;
wire            n11007;
wire            n11008;
wire            n11009;
wire      [7:0] n1101;
wire            n11010;
wire            n11011;
wire      [7:0] n11012;
wire            n11013;
wire            n11014;
wire            n11015;
wire            n11016;
wire            n11017;
wire      [7:0] n11018;
wire            n11019;
wire      [7:0] n1102;
wire            n11020;
wire            n11021;
wire            n11022;
wire            n11023;
wire      [7:0] n11024;
wire            n11025;
wire            n11026;
wire            n11027;
wire            n11028;
wire            n11029;
wire      [7:0] n1103;
wire      [7:0] n11030;
wire            n11031;
wire            n11032;
wire            n11033;
wire            n11034;
wire            n11035;
wire      [7:0] n11036;
wire            n11037;
wire            n11038;
wire            n11039;
wire      [7:0] n1104;
wire            n11040;
wire            n11041;
wire      [7:0] n11042;
wire            n11043;
wire            n11044;
wire            n11045;
wire            n11046;
wire            n11047;
wire      [7:0] n11048;
wire            n11049;
wire      [7:0] n1105;
wire            n11050;
wire            n11051;
wire            n11052;
wire            n11053;
wire      [7:0] n11054;
wire            n11055;
wire            n11056;
wire            n11057;
wire            n11058;
wire            n11059;
wire      [7:0] n1106;
wire      [7:0] n11060;
wire            n11061;
wire            n11062;
wire            n11063;
wire            n11064;
wire            n11065;
wire      [7:0] n11066;
wire            n11067;
wire            n11068;
wire            n11069;
wire      [7:0] n1107;
wire            n11070;
wire            n11071;
wire      [7:0] n11072;
wire            n11073;
wire            n11074;
wire            n11075;
wire            n11076;
wire            n11077;
wire      [7:0] n11078;
wire            n11079;
wire      [7:0] n1108;
wire            n11080;
wire            n11081;
wire            n11082;
wire            n11083;
wire      [7:0] n11084;
wire            n11085;
wire            n11086;
wire            n11087;
wire            n11088;
wire            n11089;
wire      [7:0] n1109;
wire      [7:0] n11090;
wire            n11091;
wire            n11092;
wire            n11093;
wire            n11094;
wire            n11095;
wire      [7:0] n11096;
wire            n11097;
wire            n11098;
wire            n11099;
wire      [7:0] n1110;
wire            n11100;
wire            n11101;
wire      [7:0] n11102;
wire            n11103;
wire            n11104;
wire            n11105;
wire            n11106;
wire            n11107;
wire      [7:0] n11108;
wire            n11109;
wire      [7:0] n1111;
wire            n11110;
wire            n11111;
wire            n11112;
wire            n11113;
wire      [7:0] n11114;
wire            n11115;
wire            n11116;
wire            n11117;
wire            n11118;
wire            n11119;
wire      [7:0] n1112;
wire      [7:0] n11120;
wire            n11121;
wire            n11122;
wire            n11123;
wire            n11124;
wire            n11125;
wire      [7:0] n11126;
wire            n11127;
wire            n11128;
wire            n11129;
wire      [7:0] n1113;
wire            n11130;
wire            n11131;
wire      [7:0] n11132;
wire            n11133;
wire            n11134;
wire            n11135;
wire            n11136;
wire            n11137;
wire      [7:0] n11138;
wire            n11139;
wire      [7:0] n1114;
wire            n11140;
wire            n11141;
wire            n11142;
wire            n11143;
wire      [7:0] n11144;
wire            n11145;
wire            n11146;
wire            n11147;
wire            n11148;
wire            n11149;
wire      [7:0] n1115;
wire      [7:0] n11150;
wire            n11151;
wire            n11152;
wire            n11153;
wire            n11154;
wire            n11155;
wire      [7:0] n11156;
wire            n11157;
wire            n11158;
wire            n11159;
wire      [7:0] n1116;
wire            n11160;
wire            n11161;
wire      [7:0] n11162;
wire            n11163;
wire            n11164;
wire            n11165;
wire            n11166;
wire            n11167;
wire      [7:0] n11168;
wire            n11169;
wire      [7:0] n1117;
wire            n11170;
wire            n11171;
wire            n11172;
wire            n11173;
wire      [7:0] n11174;
wire            n11175;
wire            n11176;
wire            n11177;
wire            n11178;
wire            n11179;
wire      [7:0] n1118;
wire      [7:0] n11180;
wire            n11181;
wire            n11182;
wire            n11183;
wire            n11184;
wire            n11185;
wire      [7:0] n11186;
wire            n11187;
wire            n11188;
wire            n11189;
wire      [7:0] n1119;
wire            n11190;
wire            n11191;
wire      [7:0] n11192;
wire            n11193;
wire            n11194;
wire            n11195;
wire            n11196;
wire            n11197;
wire      [7:0] n11198;
wire            n11199;
wire            n112;
wire      [7:0] n1120;
wire            n11200;
wire            n11201;
wire            n11202;
wire            n11203;
wire      [7:0] n11204;
wire            n11205;
wire            n11206;
wire            n11207;
wire            n11208;
wire            n11209;
wire      [7:0] n1121;
wire      [7:0] n11210;
wire            n11211;
wire            n11212;
wire            n11213;
wire            n11214;
wire            n11215;
wire      [7:0] n11216;
wire            n11217;
wire            n11218;
wire            n11219;
wire      [7:0] n1122;
wire            n11220;
wire            n11221;
wire      [7:0] n11222;
wire            n11223;
wire            n11224;
wire            n11225;
wire            n11226;
wire            n11227;
wire      [7:0] n11228;
wire            n11229;
wire      [7:0] n1123;
wire            n11230;
wire            n11231;
wire            n11232;
wire            n11233;
wire      [7:0] n11234;
wire            n11235;
wire            n11236;
wire            n11237;
wire            n11238;
wire            n11239;
wire      [7:0] n1124;
wire      [7:0] n11240;
wire            n11241;
wire            n11242;
wire            n11243;
wire            n11244;
wire            n11245;
wire      [7:0] n11246;
wire            n11247;
wire            n11248;
wire            n11249;
wire      [7:0] n1125;
wire            n11250;
wire            n11251;
wire      [7:0] n11252;
wire            n11253;
wire            n11254;
wire            n11255;
wire            n11256;
wire            n11257;
wire      [7:0] n11258;
wire            n11259;
wire      [7:0] n1126;
wire            n11260;
wire            n11261;
wire            n11262;
wire            n11263;
wire      [7:0] n11264;
wire            n11265;
wire            n11266;
wire            n11267;
wire            n11268;
wire            n11269;
wire      [7:0] n1127;
wire      [7:0] n11270;
wire            n11271;
wire            n11272;
wire            n11273;
wire            n11274;
wire            n11275;
wire      [7:0] n11276;
wire            n11277;
wire            n11278;
wire            n11279;
wire      [7:0] n1128;
wire            n11280;
wire            n11281;
wire      [7:0] n11282;
wire            n11283;
wire            n11284;
wire            n11285;
wire            n11286;
wire            n11287;
wire      [7:0] n11288;
wire            n11289;
wire      [7:0] n1129;
wire            n11290;
wire            n11291;
wire            n11292;
wire            n11293;
wire      [7:0] n11294;
wire            n11295;
wire            n11296;
wire            n11297;
wire            n11298;
wire            n11299;
wire      [7:0] n1130;
wire      [7:0] n11300;
wire            n11301;
wire            n11302;
wire            n11303;
wire            n11304;
wire            n11305;
wire      [7:0] n11306;
wire            n11307;
wire            n11308;
wire            n11309;
wire      [7:0] n1131;
wire            n11310;
wire            n11311;
wire      [7:0] n11312;
wire            n11313;
wire            n11314;
wire            n11315;
wire            n11316;
wire            n11317;
wire      [7:0] n11318;
wire            n11319;
wire      [7:0] n1132;
wire            n11320;
wire            n11321;
wire            n11322;
wire            n11323;
wire      [7:0] n11324;
wire            n11325;
wire            n11326;
wire            n11327;
wire            n11328;
wire            n11329;
wire      [7:0] n1133;
wire      [7:0] n11330;
wire            n11331;
wire            n11332;
wire            n11333;
wire            n11334;
wire            n11335;
wire      [7:0] n11336;
wire            n11337;
wire            n11338;
wire            n11339;
wire      [7:0] n1134;
wire            n11340;
wire            n11341;
wire      [7:0] n11342;
wire            n11343;
wire            n11344;
wire            n11345;
wire            n11346;
wire            n11347;
wire      [7:0] n11348;
wire            n11349;
wire      [7:0] n1135;
wire            n11350;
wire            n11351;
wire            n11352;
wire            n11353;
wire      [7:0] n11354;
wire            n11355;
wire            n11356;
wire            n11357;
wire            n11358;
wire            n11359;
wire      [7:0] n1136;
wire      [7:0] n11360;
wire            n11361;
wire            n11362;
wire            n11363;
wire            n11364;
wire            n11365;
wire      [7:0] n11366;
wire            n11367;
wire            n11368;
wire            n11369;
wire      [7:0] n1137;
wire            n11370;
wire            n11371;
wire      [7:0] n11372;
wire            n11373;
wire            n11374;
wire            n11375;
wire            n11376;
wire            n11377;
wire      [7:0] n11378;
wire            n11379;
wire      [7:0] n1138;
wire            n11380;
wire            n11381;
wire            n11382;
wire            n11383;
wire      [7:0] n11384;
wire            n11385;
wire            n11386;
wire            n11387;
wire            n11388;
wire            n11389;
wire      [7:0] n1139;
wire      [7:0] n11390;
wire            n11391;
wire            n11392;
wire            n11393;
wire            n11394;
wire            n11395;
wire      [7:0] n11396;
wire            n11397;
wire            n11398;
wire            n11399;
wire            n114;
wire      [7:0] n1140;
wire            n11400;
wire            n11401;
wire      [7:0] n11402;
wire            n11403;
wire            n11404;
wire            n11405;
wire            n11406;
wire            n11407;
wire      [7:0] n11408;
wire            n11409;
wire      [7:0] n1141;
wire            n11410;
wire            n11411;
wire            n11412;
wire            n11413;
wire      [7:0] n11414;
wire            n11415;
wire            n11416;
wire            n11417;
wire            n11418;
wire            n11419;
wire      [7:0] n1142;
wire      [7:0] n11420;
wire            n11421;
wire            n11422;
wire            n11423;
wire            n11424;
wire            n11425;
wire      [7:0] n11426;
wire            n11427;
wire            n11428;
wire            n11429;
wire      [7:0] n1143;
wire            n11430;
wire            n11431;
wire      [7:0] n11432;
wire            n11433;
wire            n11434;
wire            n11435;
wire            n11436;
wire            n11437;
wire      [7:0] n11438;
wire            n11439;
wire      [7:0] n1144;
wire            n11440;
wire            n11441;
wire            n11442;
wire            n11443;
wire      [7:0] n11444;
wire            n11445;
wire            n11446;
wire            n11447;
wire            n11448;
wire            n11449;
wire      [7:0] n1145;
wire      [7:0] n11450;
wire            n11451;
wire            n11452;
wire            n11453;
wire            n11454;
wire            n11455;
wire      [7:0] n11456;
wire            n11457;
wire            n11458;
wire            n11459;
wire      [7:0] n1146;
wire            n11460;
wire            n11461;
wire      [7:0] n11462;
wire            n11463;
wire            n11464;
wire            n11465;
wire            n11466;
wire            n11467;
wire      [7:0] n11468;
wire            n11469;
wire      [7:0] n1147;
wire            n11470;
wire            n11471;
wire            n11472;
wire            n11473;
wire      [7:0] n11474;
wire            n11475;
wire            n11476;
wire            n11477;
wire            n11478;
wire            n11479;
wire      [7:0] n1148;
wire      [7:0] n11480;
wire            n11481;
wire            n11482;
wire            n11483;
wire            n11484;
wire            n11485;
wire      [7:0] n11486;
wire            n11487;
wire            n11488;
wire            n11489;
wire      [7:0] n1149;
wire            n11490;
wire            n11491;
wire      [7:0] n11492;
wire            n11493;
wire            n11494;
wire            n11495;
wire            n11496;
wire            n11497;
wire      [7:0] n11498;
wire            n11499;
wire      [7:0] n1150;
wire            n11500;
wire            n11501;
wire            n11502;
wire            n11503;
wire      [7:0] n11504;
wire            n11505;
wire            n11506;
wire            n11507;
wire            n11508;
wire            n11509;
wire      [7:0] n1151;
wire      [7:0] n11510;
wire            n11511;
wire            n11512;
wire            n11513;
wire            n11514;
wire            n11515;
wire      [7:0] n11516;
wire            n11517;
wire            n11518;
wire            n11519;
wire      [7:0] n1152;
wire            n11520;
wire            n11521;
wire      [7:0] n11522;
wire            n11523;
wire            n11524;
wire            n11525;
wire            n11526;
wire            n11527;
wire      [7:0] n11528;
wire            n11529;
wire      [7:0] n1153;
wire            n11530;
wire            n11531;
wire            n11532;
wire            n11533;
wire      [7:0] n11534;
wire            n11535;
wire            n11536;
wire            n11537;
wire            n11538;
wire            n11539;
wire      [7:0] n1154;
wire      [7:0] n11540;
wire            n11541;
wire            n11542;
wire            n11543;
wire            n11544;
wire            n11545;
wire      [7:0] n11546;
wire            n11547;
wire            n11548;
wire            n11549;
wire      [7:0] n1155;
wire            n11550;
wire            n11551;
wire      [7:0] n11552;
wire            n11553;
wire            n11554;
wire            n11555;
wire            n11556;
wire            n11557;
wire      [7:0] n11558;
wire            n11559;
wire      [7:0] n1156;
wire            n11560;
wire            n11561;
wire            n11562;
wire            n11563;
wire      [7:0] n11564;
wire            n11565;
wire            n11566;
wire            n11567;
wire            n11568;
wire            n11569;
wire      [7:0] n1157;
wire      [7:0] n11570;
wire            n11571;
wire            n11572;
wire            n11573;
wire            n11574;
wire            n11575;
wire      [7:0] n11576;
wire            n11577;
wire            n11578;
wire            n11579;
wire      [7:0] n1158;
wire            n11580;
wire            n11581;
wire      [7:0] n11582;
wire            n11583;
wire            n11584;
wire            n11585;
wire            n11586;
wire            n11587;
wire      [7:0] n11588;
wire            n11589;
wire      [7:0] n1159;
wire            n11590;
wire            n11591;
wire            n11592;
wire            n11593;
wire      [7:0] n11594;
wire            n11595;
wire            n11596;
wire            n11597;
wire            n11598;
wire            n11599;
wire            n116;
wire      [7:0] n1160;
wire      [7:0] n11600;
wire            n11601;
wire            n11602;
wire            n11603;
wire            n11604;
wire            n11605;
wire      [7:0] n11606;
wire            n11607;
wire            n11608;
wire            n11609;
wire      [7:0] n1161;
wire            n11610;
wire            n11611;
wire      [7:0] n11612;
wire            n11613;
wire            n11614;
wire            n11615;
wire            n11616;
wire            n11617;
wire      [7:0] n11618;
wire            n11619;
wire      [7:0] n1162;
wire            n11620;
wire            n11621;
wire            n11622;
wire            n11623;
wire      [7:0] n11624;
wire            n11625;
wire            n11626;
wire            n11627;
wire            n11628;
wire            n11629;
wire      [7:0] n1163;
wire      [7:0] n11630;
wire            n11631;
wire            n11632;
wire            n11633;
wire            n11634;
wire            n11635;
wire      [7:0] n11636;
wire            n11637;
wire            n11638;
wire            n11639;
wire      [7:0] n1164;
wire            n11640;
wire            n11641;
wire      [7:0] n11642;
wire            n11643;
wire            n11644;
wire            n11645;
wire            n11646;
wire            n11647;
wire      [7:0] n11648;
wire            n11649;
wire      [7:0] n1165;
wire            n11650;
wire            n11651;
wire            n11652;
wire            n11653;
wire      [7:0] n11654;
wire            n11655;
wire            n11656;
wire            n11657;
wire            n11658;
wire            n11659;
wire      [7:0] n1166;
wire      [7:0] n11660;
wire            n11661;
wire            n11662;
wire            n11663;
wire            n11664;
wire            n11665;
wire      [7:0] n11666;
wire            n11667;
wire            n11668;
wire            n11669;
wire      [7:0] n1167;
wire            n11670;
wire            n11671;
wire      [7:0] n11672;
wire            n11673;
wire            n11674;
wire            n11675;
wire            n11676;
wire            n11677;
wire      [7:0] n11678;
wire            n11679;
wire      [7:0] n1168;
wire            n11680;
wire            n11681;
wire            n11682;
wire            n11683;
wire      [7:0] n11684;
wire            n11685;
wire            n11686;
wire            n11687;
wire            n11688;
wire            n11689;
wire      [7:0] n1169;
wire      [7:0] n11690;
wire            n11691;
wire            n11692;
wire            n11693;
wire            n11694;
wire            n11695;
wire      [7:0] n11696;
wire            n11697;
wire            n11698;
wire            n11699;
wire      [7:0] n1170;
wire            n11700;
wire            n11701;
wire      [7:0] n11702;
wire            n11703;
wire            n11704;
wire            n11705;
wire            n11706;
wire            n11707;
wire      [7:0] n11708;
wire            n11709;
wire      [7:0] n1171;
wire            n11710;
wire            n11711;
wire            n11712;
wire            n11713;
wire      [7:0] n11714;
wire            n11715;
wire            n11716;
wire            n11717;
wire            n11718;
wire            n11719;
wire      [7:0] n1172;
wire      [7:0] n11720;
wire            n11721;
wire            n11722;
wire            n11723;
wire            n11724;
wire            n11725;
wire      [7:0] n11726;
wire            n11727;
wire            n11728;
wire            n11729;
wire      [7:0] n1173;
wire            n11730;
wire            n11731;
wire      [7:0] n11732;
wire            n11733;
wire            n11734;
wire            n11735;
wire            n11736;
wire            n11737;
wire      [7:0] n11738;
wire            n11739;
wire      [7:0] n1174;
wire            n11740;
wire            n11741;
wire            n11742;
wire            n11743;
wire      [7:0] n11744;
wire            n11745;
wire            n11746;
wire            n11747;
wire            n11748;
wire            n11749;
wire      [7:0] n1175;
wire      [7:0] n11750;
wire            n11751;
wire            n11752;
wire            n11753;
wire            n11754;
wire            n11755;
wire      [7:0] n11756;
wire            n11757;
wire            n11758;
wire            n11759;
wire      [7:0] n1176;
wire            n11760;
wire            n11761;
wire      [7:0] n11762;
wire            n11763;
wire            n11764;
wire            n11765;
wire            n11766;
wire            n11767;
wire      [7:0] n11768;
wire            n11769;
wire      [7:0] n1177;
wire            n11770;
wire            n11771;
wire            n11772;
wire            n11773;
wire      [7:0] n11774;
wire            n11775;
wire            n11776;
wire            n11777;
wire            n11778;
wire            n11779;
wire      [7:0] n1178;
wire      [7:0] n11780;
wire            n11781;
wire            n11782;
wire            n11783;
wire            n11784;
wire            n11785;
wire      [7:0] n11786;
wire            n11787;
wire            n11788;
wire            n11789;
wire      [7:0] n1179;
wire            n11790;
wire            n11791;
wire      [7:0] n11792;
wire            n11793;
wire            n11794;
wire            n11795;
wire            n11796;
wire            n11797;
wire      [7:0] n11798;
wire            n11799;
wire            n118;
wire      [7:0] n1180;
wire            n11800;
wire            n11801;
wire            n11802;
wire            n11803;
wire      [7:0] n11804;
wire            n11805;
wire            n11806;
wire            n11807;
wire            n11808;
wire            n11809;
wire      [7:0] n1181;
wire      [7:0] n11810;
wire            n11811;
wire            n11812;
wire            n11813;
wire            n11814;
wire            n11815;
wire      [7:0] n11816;
wire            n11817;
wire            n11818;
wire            n11819;
wire      [7:0] n1182;
wire            n11820;
wire            n11821;
wire      [7:0] n11822;
wire            n11823;
wire            n11824;
wire            n11825;
wire            n11826;
wire            n11827;
wire      [7:0] n11828;
wire            n11829;
wire      [7:0] n1183;
wire            n11830;
wire            n11831;
wire            n11832;
wire            n11833;
wire      [7:0] n11834;
wire            n11835;
wire            n11836;
wire            n11837;
wire            n11838;
wire            n11839;
wire      [7:0] n1184;
wire      [7:0] n11840;
wire            n11841;
wire            n11842;
wire            n11843;
wire            n11844;
wire            n11845;
wire      [7:0] n11846;
wire            n11847;
wire            n11848;
wire            n11849;
wire      [7:0] n1185;
wire            n11850;
wire            n11851;
wire      [7:0] n11852;
wire            n11853;
wire            n11854;
wire            n11855;
wire            n11856;
wire            n11857;
wire      [7:0] n11858;
wire            n11859;
wire      [7:0] n1186;
wire            n11860;
wire            n11861;
wire            n11862;
wire            n11863;
wire      [7:0] n11864;
wire            n11865;
wire            n11866;
wire            n11867;
wire            n11868;
wire            n11869;
wire      [7:0] n1187;
wire      [7:0] n11870;
wire            n11871;
wire            n11872;
wire            n11873;
wire            n11874;
wire            n11875;
wire      [7:0] n11876;
wire            n11877;
wire            n11878;
wire            n11879;
wire      [7:0] n1188;
wire            n11880;
wire            n11881;
wire      [7:0] n11882;
wire            n11883;
wire            n11884;
wire            n11885;
wire            n11886;
wire            n11887;
wire      [7:0] n11888;
wire            n11889;
wire      [7:0] n1189;
wire            n11890;
wire            n11891;
wire            n11892;
wire            n11893;
wire      [7:0] n11894;
wire            n11895;
wire            n11896;
wire            n11897;
wire            n11898;
wire            n11899;
wire      [7:0] n1190;
wire      [7:0] n11900;
wire            n11901;
wire            n11902;
wire            n11903;
wire            n11904;
wire            n11905;
wire      [7:0] n11906;
wire            n11907;
wire            n11908;
wire            n11909;
wire      [7:0] n1191;
wire            n11910;
wire            n11911;
wire      [7:0] n11912;
wire            n11913;
wire            n11914;
wire            n11915;
wire            n11916;
wire            n11917;
wire      [7:0] n11918;
wire            n11919;
wire      [7:0] n1192;
wire            n11920;
wire            n11921;
wire            n11922;
wire            n11923;
wire      [7:0] n11924;
wire            n11925;
wire            n11926;
wire            n11927;
wire            n11928;
wire            n11929;
wire      [7:0] n1193;
wire      [7:0] n11930;
wire            n11931;
wire            n11932;
wire            n11933;
wire            n11934;
wire            n11935;
wire      [7:0] n11936;
wire            n11937;
wire            n11938;
wire            n11939;
wire      [7:0] n1194;
wire            n11940;
wire            n11941;
wire      [7:0] n11942;
wire            n11943;
wire            n11944;
wire            n11945;
wire            n11946;
wire            n11947;
wire      [7:0] n11948;
wire            n11949;
wire      [7:0] n1195;
wire            n11950;
wire            n11951;
wire            n11952;
wire            n11953;
wire      [7:0] n11954;
wire            n11955;
wire            n11956;
wire            n11957;
wire            n11958;
wire            n11959;
wire      [7:0] n1196;
wire      [7:0] n11960;
wire            n11961;
wire            n11962;
wire            n11963;
wire            n11964;
wire            n11965;
wire      [7:0] n11966;
wire            n11967;
wire            n11968;
wire            n11969;
wire      [7:0] n1197;
wire            n11970;
wire            n11971;
wire      [7:0] n11972;
wire            n11973;
wire            n11974;
wire            n11975;
wire            n11976;
wire            n11977;
wire      [7:0] n11978;
wire            n11979;
wire      [7:0] n1198;
wire            n11980;
wire            n11981;
wire            n11982;
wire            n11983;
wire      [7:0] n11984;
wire            n11985;
wire            n11986;
wire            n11987;
wire            n11988;
wire            n11989;
wire      [7:0] n1199;
wire      [7:0] n11990;
wire            n11991;
wire            n11992;
wire            n11993;
wire            n11994;
wire            n11995;
wire      [7:0] n11996;
wire            n11997;
wire            n11998;
wire            n11999;
wire            n120;
wire      [7:0] n1200;
wire            n12000;
wire            n12001;
wire      [7:0] n12002;
wire            n12003;
wire            n12004;
wire            n12005;
wire            n12006;
wire            n12007;
wire      [7:0] n12008;
wire            n12009;
wire      [7:0] n1201;
wire            n12010;
wire            n12011;
wire            n12012;
wire            n12013;
wire      [7:0] n12014;
wire            n12015;
wire            n12016;
wire            n12017;
wire            n12018;
wire            n12019;
wire      [7:0] n1202;
wire      [7:0] n12020;
wire            n12021;
wire            n12022;
wire            n12023;
wire            n12024;
wire            n12025;
wire      [7:0] n12026;
wire            n12027;
wire            n12028;
wire            n12029;
wire      [7:0] n1203;
wire            n12030;
wire            n12031;
wire      [7:0] n12032;
wire            n12033;
wire            n12034;
wire            n12035;
wire            n12036;
wire            n12037;
wire      [7:0] n12038;
wire            n12039;
wire      [7:0] n1204;
wire            n12040;
wire            n12041;
wire            n12042;
wire            n12043;
wire      [7:0] n12044;
wire            n12045;
wire            n12046;
wire            n12047;
wire            n12048;
wire            n12049;
wire      [7:0] n1205;
wire      [7:0] n12050;
wire            n12051;
wire            n12052;
wire            n12053;
wire            n12054;
wire            n12055;
wire      [7:0] n12056;
wire            n12057;
wire            n12058;
wire            n12059;
wire      [7:0] n1206;
wire            n12060;
wire            n12061;
wire      [7:0] n12062;
wire            n12063;
wire            n12064;
wire            n12065;
wire            n12066;
wire            n12067;
wire      [7:0] n12068;
wire            n12069;
wire      [7:0] n1207;
wire            n12070;
wire            n12071;
wire            n12072;
wire            n12073;
wire      [7:0] n12074;
wire            n12075;
wire            n12076;
wire            n12077;
wire            n12078;
wire            n12079;
wire      [7:0] n1208;
wire      [7:0] n12080;
wire            n12081;
wire            n12082;
wire            n12083;
wire            n12084;
wire            n12085;
wire      [7:0] n12086;
wire            n12087;
wire            n12088;
wire            n12089;
wire      [7:0] n1209;
wire            n12090;
wire            n12091;
wire      [7:0] n12092;
wire            n12093;
wire            n12094;
wire            n12095;
wire            n12096;
wire            n12097;
wire      [7:0] n12098;
wire            n12099;
wire      [7:0] n1210;
wire            n12100;
wire            n12101;
wire            n12102;
wire            n12103;
wire      [7:0] n12104;
wire            n12105;
wire            n12106;
wire            n12107;
wire            n12108;
wire            n12109;
wire      [7:0] n1211;
wire      [7:0] n12110;
wire            n12111;
wire            n12112;
wire            n12113;
wire            n12114;
wire            n12115;
wire      [7:0] n12116;
wire            n12117;
wire            n12118;
wire            n12119;
wire      [7:0] n1212;
wire            n12120;
wire            n12121;
wire      [7:0] n12122;
wire            n12123;
wire            n12124;
wire            n12125;
wire            n12126;
wire            n12127;
wire      [7:0] n12128;
wire            n12129;
wire      [7:0] n1213;
wire            n12130;
wire            n12131;
wire            n12132;
wire            n12133;
wire      [7:0] n12134;
wire            n12135;
wire            n12136;
wire            n12137;
wire            n12138;
wire            n12139;
wire      [7:0] n1214;
wire      [7:0] n12140;
wire            n12141;
wire            n12142;
wire            n12143;
wire            n12144;
wire            n12145;
wire      [7:0] n12146;
wire            n12147;
wire            n12148;
wire            n12149;
wire      [7:0] n1215;
wire            n12150;
wire            n12151;
wire      [7:0] n12152;
wire            n12153;
wire            n12154;
wire            n12155;
wire            n12156;
wire            n12157;
wire      [7:0] n12158;
wire            n12159;
wire      [7:0] n1216;
wire            n12160;
wire            n12161;
wire            n12162;
wire            n12163;
wire      [7:0] n12164;
wire            n12165;
wire            n12166;
wire            n12167;
wire            n12168;
wire            n12169;
wire      [7:0] n1217;
wire      [7:0] n12170;
wire            n12171;
wire            n12172;
wire            n12173;
wire            n12174;
wire            n12175;
wire      [7:0] n12176;
wire            n12177;
wire            n12178;
wire            n12179;
wire      [7:0] n1218;
wire            n12180;
wire            n12181;
wire      [7:0] n12182;
wire            n12183;
wire            n12184;
wire            n12185;
wire            n12186;
wire            n12187;
wire      [7:0] n12188;
wire            n12189;
wire      [7:0] n1219;
wire            n12190;
wire            n12191;
wire            n12192;
wire            n12193;
wire      [7:0] n12194;
wire            n12195;
wire            n12196;
wire            n12197;
wire            n12198;
wire            n12199;
wire            n122;
wire      [7:0] n1220;
wire      [7:0] n12200;
wire            n12201;
wire            n12202;
wire            n12203;
wire            n12204;
wire            n12205;
wire      [7:0] n12206;
wire            n12207;
wire            n12208;
wire            n12209;
wire      [7:0] n1221;
wire            n12210;
wire            n12211;
wire      [7:0] n12212;
wire            n12213;
wire            n12214;
wire            n12215;
wire            n12216;
wire            n12217;
wire      [7:0] n12218;
wire            n12219;
wire      [7:0] n1222;
wire            n12220;
wire            n12221;
wire            n12222;
wire            n12223;
wire      [7:0] n12224;
wire            n12225;
wire            n12226;
wire            n12227;
wire            n12228;
wire            n12229;
wire      [7:0] n1223;
wire      [7:0] n12230;
wire            n12231;
wire            n12232;
wire            n12233;
wire            n12234;
wire            n12235;
wire      [7:0] n12236;
wire            n12237;
wire            n12238;
wire            n12239;
wire      [7:0] n1224;
wire            n12240;
wire            n12241;
wire      [7:0] n12242;
wire            n12243;
wire            n12244;
wire            n12245;
wire            n12246;
wire            n12247;
wire      [7:0] n12248;
wire            n12249;
wire      [7:0] n1225;
wire            n12250;
wire            n12251;
wire            n12252;
wire            n12253;
wire      [7:0] n12254;
wire            n12255;
wire            n12256;
wire            n12257;
wire            n12258;
wire            n12259;
wire      [7:0] n1226;
wire      [7:0] n12260;
wire            n12261;
wire            n12262;
wire            n12263;
wire            n12264;
wire            n12265;
wire      [7:0] n12266;
wire            n12267;
wire            n12268;
wire            n12269;
wire      [7:0] n1227;
wire            n12270;
wire            n12271;
wire      [7:0] n12272;
wire            n12273;
wire            n12274;
wire            n12275;
wire            n12276;
wire            n12277;
wire      [7:0] n12278;
wire            n12279;
wire      [7:0] n1228;
wire            n12280;
wire            n12281;
wire            n12282;
wire            n12283;
wire      [7:0] n12284;
wire            n12285;
wire            n12286;
wire            n12287;
wire            n12288;
wire            n12289;
wire      [7:0] n1229;
wire      [7:0] n12290;
wire            n12291;
wire            n12292;
wire            n12293;
wire            n12294;
wire            n12295;
wire      [7:0] n12296;
wire            n12297;
wire            n12298;
wire            n12299;
wire      [7:0] n1230;
wire            n12300;
wire            n12301;
wire      [7:0] n12302;
wire            n12303;
wire            n12304;
wire            n12305;
wire            n12306;
wire            n12307;
wire      [7:0] n12308;
wire            n12309;
wire      [7:0] n1231;
wire            n12310;
wire            n12311;
wire            n12312;
wire            n12313;
wire      [7:0] n12314;
wire            n12315;
wire            n12316;
wire            n12317;
wire            n12318;
wire            n12319;
wire      [7:0] n1232;
wire      [7:0] n12320;
wire            n12321;
wire            n12322;
wire            n12323;
wire            n12324;
wire            n12325;
wire      [7:0] n12326;
wire            n12327;
wire            n12328;
wire            n12329;
wire      [7:0] n1233;
wire            n12330;
wire            n12331;
wire      [7:0] n12332;
wire            n12333;
wire            n12334;
wire            n12335;
wire            n12336;
wire            n12337;
wire      [7:0] n12338;
wire            n12339;
wire      [7:0] n1234;
wire            n12340;
wire            n12341;
wire            n12342;
wire            n12343;
wire      [7:0] n12344;
wire            n12345;
wire            n12346;
wire            n12347;
wire            n12348;
wire            n12349;
wire      [7:0] n1235;
wire      [7:0] n12350;
wire            n12351;
wire            n12352;
wire            n12353;
wire            n12354;
wire            n12355;
wire      [7:0] n12356;
wire            n12357;
wire            n12358;
wire            n12359;
wire      [7:0] n1236;
wire            n12360;
wire            n12361;
wire      [7:0] n12362;
wire            n12363;
wire            n12364;
wire            n12365;
wire            n12366;
wire            n12367;
wire      [7:0] n12368;
wire            n12369;
wire      [7:0] n1237;
wire            n12370;
wire            n12371;
wire            n12372;
wire            n12373;
wire      [7:0] n12374;
wire            n12375;
wire            n12376;
wire            n12377;
wire            n12378;
wire            n12379;
wire      [7:0] n1238;
wire      [7:0] n12380;
wire            n12381;
wire            n12382;
wire            n12383;
wire            n12384;
wire            n12385;
wire      [7:0] n12386;
wire            n12387;
wire            n12388;
wire            n12389;
wire      [7:0] n1239;
wire            n12390;
wire            n12391;
wire      [7:0] n12392;
wire            n12393;
wire            n12394;
wire            n12395;
wire            n12396;
wire            n12397;
wire      [7:0] n12398;
wire            n12399;
wire            n124;
wire      [7:0] n1240;
wire            n12400;
wire            n12401;
wire            n12402;
wire            n12403;
wire      [7:0] n12404;
wire            n12405;
wire            n12406;
wire            n12407;
wire            n12408;
wire            n12409;
wire      [7:0] n1241;
wire      [7:0] n12410;
wire            n12411;
wire            n12412;
wire            n12413;
wire            n12414;
wire            n12415;
wire      [7:0] n12416;
wire            n12417;
wire            n12418;
wire            n12419;
wire      [7:0] n1242;
wire            n12420;
wire            n12421;
wire      [7:0] n12422;
wire            n12423;
wire            n12424;
wire            n12425;
wire            n12426;
wire            n12427;
wire      [7:0] n12428;
wire            n12429;
wire      [7:0] n1243;
wire            n12430;
wire            n12431;
wire            n12432;
wire            n12433;
wire      [7:0] n12434;
wire            n12435;
wire            n12436;
wire            n12437;
wire            n12438;
wire            n12439;
wire      [7:0] n1244;
wire      [7:0] n12440;
wire            n12441;
wire            n12442;
wire            n12443;
wire            n12444;
wire            n12445;
wire      [7:0] n12446;
wire            n12447;
wire            n12448;
wire            n12449;
wire      [7:0] n1245;
wire            n12450;
wire            n12451;
wire      [7:0] n12452;
wire            n12453;
wire            n12454;
wire            n12455;
wire            n12456;
wire            n12457;
wire      [7:0] n12458;
wire            n12459;
wire      [7:0] n1246;
wire            n12460;
wire            n12461;
wire            n12462;
wire            n12463;
wire      [7:0] n12464;
wire            n12465;
wire            n12466;
wire            n12467;
wire            n12468;
wire            n12469;
wire      [7:0] n1247;
wire      [7:0] n12470;
wire            n12471;
wire            n12472;
wire            n12473;
wire            n12474;
wire            n12475;
wire      [7:0] n12476;
wire            n12477;
wire            n12478;
wire            n12479;
wire      [7:0] n1248;
wire            n12480;
wire            n12481;
wire      [7:0] n12482;
wire            n12483;
wire            n12484;
wire            n12485;
wire            n12486;
wire            n12487;
wire      [7:0] n12488;
wire            n12489;
wire      [7:0] n1249;
wire            n12490;
wire            n12491;
wire            n12492;
wire            n12493;
wire      [7:0] n12494;
wire            n12495;
wire            n12496;
wire            n12497;
wire            n12498;
wire            n12499;
wire      [7:0] n1250;
wire      [7:0] n12500;
wire            n12501;
wire            n12502;
wire            n12503;
wire            n12504;
wire            n12505;
wire      [7:0] n12506;
wire            n12507;
wire            n12508;
wire            n12509;
wire      [7:0] n1251;
wire            n12510;
wire            n12511;
wire      [7:0] n12512;
wire            n12513;
wire            n12514;
wire            n12515;
wire            n12516;
wire            n12517;
wire      [7:0] n12518;
wire            n12519;
wire      [7:0] n1252;
wire            n12520;
wire            n12521;
wire            n12522;
wire            n12523;
wire      [7:0] n12524;
wire            n12525;
wire            n12526;
wire            n12527;
wire            n12528;
wire            n12529;
wire      [7:0] n1253;
wire      [7:0] n12530;
wire            n12531;
wire            n12532;
wire            n12533;
wire            n12534;
wire            n12535;
wire      [7:0] n12536;
wire            n12537;
wire            n12538;
wire            n12539;
wire      [7:0] n1254;
wire            n12540;
wire            n12541;
wire      [7:0] n12542;
wire            n12543;
wire            n12544;
wire            n12545;
wire            n12546;
wire            n12547;
wire      [7:0] n12548;
wire            n12549;
wire      [7:0] n1255;
wire            n12550;
wire            n12551;
wire            n12552;
wire            n12553;
wire      [7:0] n12554;
wire            n12555;
wire            n12556;
wire            n12557;
wire            n12558;
wire            n12559;
wire      [7:0] n1256;
wire      [7:0] n12560;
wire            n12561;
wire            n12562;
wire            n12563;
wire            n12564;
wire            n12565;
wire      [7:0] n12566;
wire            n12567;
wire            n12568;
wire            n12569;
wire      [7:0] n1257;
wire            n12570;
wire            n12571;
wire      [7:0] n12572;
wire            n12573;
wire            n12574;
wire            n12575;
wire            n12576;
wire            n12577;
wire      [7:0] n12578;
wire            n12579;
wire      [7:0] n1258;
wire            n12580;
wire            n12581;
wire            n12582;
wire            n12583;
wire      [7:0] n12584;
wire            n12585;
wire            n12586;
wire            n12587;
wire            n12588;
wire            n12589;
wire      [7:0] n1259;
wire      [7:0] n12590;
wire            n12591;
wire            n12592;
wire            n12593;
wire            n12594;
wire            n12595;
wire      [7:0] n12596;
wire            n12597;
wire            n12598;
wire            n12599;
wire            n126;
wire      [7:0] n1260;
wire            n12600;
wire            n12601;
wire      [7:0] n12602;
wire            n12603;
wire            n12604;
wire            n12605;
wire            n12606;
wire            n12607;
wire      [7:0] n12608;
wire            n12609;
wire      [7:0] n1261;
wire            n12610;
wire            n12611;
wire            n12612;
wire            n12613;
wire      [7:0] n12614;
wire            n12615;
wire            n12616;
wire            n12617;
wire            n12618;
wire            n12619;
wire      [7:0] n1262;
wire      [7:0] n12620;
wire            n12621;
wire            n12622;
wire            n12623;
wire            n12624;
wire            n12625;
wire      [7:0] n12626;
wire            n12627;
wire            n12628;
wire            n12629;
wire      [7:0] n1263;
wire            n12630;
wire            n12631;
wire      [7:0] n12632;
wire            n12633;
wire            n12634;
wire            n12635;
wire            n12636;
wire            n12637;
wire      [7:0] n12638;
wire            n12639;
wire      [7:0] n1264;
wire            n12640;
wire            n12641;
wire            n12642;
wire            n12643;
wire      [7:0] n12644;
wire            n12645;
wire            n12646;
wire            n12647;
wire            n12648;
wire            n12649;
wire      [7:0] n1265;
wire      [7:0] n12650;
wire            n12651;
wire            n12652;
wire            n12653;
wire            n12654;
wire            n12655;
wire      [7:0] n12656;
wire            n12657;
wire            n12658;
wire            n12659;
wire      [7:0] n1266;
wire            n12660;
wire            n12661;
wire      [7:0] n12662;
wire            n12663;
wire            n12664;
wire            n12665;
wire            n12666;
wire            n12667;
wire      [7:0] n12668;
wire            n12669;
wire      [7:0] n1267;
wire            n12670;
wire            n12671;
wire            n12672;
wire            n12673;
wire      [7:0] n12674;
wire            n12675;
wire            n12676;
wire            n12677;
wire            n12678;
wire            n12679;
wire      [7:0] n1268;
wire      [7:0] n12680;
wire            n12681;
wire            n12682;
wire            n12683;
wire            n12684;
wire            n12685;
wire      [7:0] n12686;
wire            n12687;
wire            n12688;
wire            n12689;
wire      [7:0] n1269;
wire            n12690;
wire            n12691;
wire      [7:0] n12692;
wire            n12693;
wire            n12694;
wire            n12695;
wire            n12696;
wire            n12697;
wire      [7:0] n12698;
wire            n12699;
wire      [7:0] n1270;
wire            n12700;
wire            n12701;
wire            n12702;
wire            n12703;
wire      [7:0] n12704;
wire            n12705;
wire            n12706;
wire            n12707;
wire            n12708;
wire            n12709;
wire      [7:0] n1271;
wire      [7:0] n12710;
wire            n12711;
wire            n12712;
wire            n12713;
wire            n12714;
wire            n12715;
wire      [7:0] n12716;
wire            n12717;
wire            n12718;
wire            n12719;
wire      [7:0] n1272;
wire            n12720;
wire            n12721;
wire      [7:0] n12722;
wire            n12723;
wire            n12724;
wire            n12725;
wire            n12726;
wire            n12727;
wire      [7:0] n12728;
wire            n12729;
wire      [7:0] n1273;
wire            n12730;
wire            n12731;
wire            n12732;
wire            n12733;
wire      [7:0] n12734;
wire            n12735;
wire            n12736;
wire            n12737;
wire            n12738;
wire            n12739;
wire      [7:0] n1274;
wire      [7:0] n12740;
wire            n12741;
wire            n12742;
wire            n12743;
wire            n12744;
wire            n12745;
wire      [7:0] n12746;
wire            n12747;
wire            n12748;
wire            n12749;
wire      [7:0] n1275;
wire            n12750;
wire            n12751;
wire      [7:0] n12752;
wire            n12753;
wire            n12754;
wire            n12755;
wire            n12756;
wire            n12757;
wire      [7:0] n12758;
wire            n12759;
wire      [7:0] n1276;
wire            n12760;
wire            n12761;
wire            n12762;
wire            n12763;
wire      [7:0] n12764;
wire            n12765;
wire            n12766;
wire            n12767;
wire            n12768;
wire            n12769;
wire      [7:0] n1277;
wire      [7:0] n12770;
wire            n12771;
wire            n12772;
wire            n12773;
wire            n12774;
wire            n12775;
wire      [7:0] n12776;
wire            n12777;
wire            n12778;
wire            n12779;
wire      [7:0] n1278;
wire            n12780;
wire            n12781;
wire      [7:0] n12782;
wire            n12783;
wire            n12784;
wire            n12785;
wire            n12786;
wire            n12787;
wire      [7:0] n12788;
wire            n12789;
wire      [7:0] n1279;
wire            n12790;
wire            n12791;
wire            n12792;
wire            n12793;
wire      [7:0] n12794;
wire            n12795;
wire            n12796;
wire            n12797;
wire            n12798;
wire            n12799;
wire            n128;
wire      [7:0] n1280;
wire      [7:0] n12800;
wire            n12801;
wire            n12802;
wire            n12803;
wire            n12804;
wire            n12805;
wire      [7:0] n12806;
wire            n12807;
wire            n12808;
wire            n12809;
wire      [7:0] n1281;
wire            n12810;
wire            n12811;
wire      [7:0] n12812;
wire            n12813;
wire            n12814;
wire            n12815;
wire            n12816;
wire            n12817;
wire      [7:0] n12818;
wire            n12819;
wire      [7:0] n1282;
wire            n12820;
wire            n12821;
wire            n12822;
wire            n12823;
wire      [7:0] n12824;
wire            n12825;
wire            n12826;
wire            n12827;
wire            n12828;
wire            n12829;
wire      [7:0] n1283;
wire      [7:0] n12830;
wire            n12831;
wire            n12832;
wire            n12833;
wire            n12834;
wire            n12835;
wire      [7:0] n12836;
wire            n12837;
wire            n12838;
wire            n12839;
wire      [7:0] n1284;
wire            n12840;
wire            n12841;
wire      [7:0] n12842;
wire            n12843;
wire            n12844;
wire            n12845;
wire            n12846;
wire            n12847;
wire      [7:0] n12848;
wire            n12849;
wire      [7:0] n1285;
wire            n12850;
wire            n12851;
wire            n12852;
wire            n12853;
wire      [7:0] n12854;
wire            n12855;
wire            n12856;
wire            n12857;
wire            n12858;
wire            n12859;
wire      [7:0] n1286;
wire      [7:0] n12860;
wire            n12861;
wire            n12862;
wire            n12863;
wire            n12864;
wire            n12865;
wire      [7:0] n12866;
wire            n12867;
wire            n12868;
wire            n12869;
wire      [7:0] n1287;
wire            n12870;
wire            n12871;
wire      [7:0] n12872;
wire            n12873;
wire            n12874;
wire            n12875;
wire            n12876;
wire            n12877;
wire      [7:0] n12878;
wire            n12879;
wire      [7:0] n1288;
wire            n12880;
wire            n12881;
wire            n12882;
wire            n12883;
wire      [7:0] n12884;
wire            n12885;
wire            n12886;
wire            n12887;
wire            n12888;
wire            n12889;
wire      [7:0] n1289;
wire      [7:0] n12890;
wire            n12891;
wire            n12892;
wire            n12893;
wire            n12894;
wire            n12895;
wire      [7:0] n12896;
wire            n12897;
wire            n12898;
wire            n12899;
wire      [7:0] n1290;
wire            n12900;
wire            n12901;
wire      [7:0] n12902;
wire            n12903;
wire            n12904;
wire            n12905;
wire            n12906;
wire            n12907;
wire      [7:0] n12908;
wire            n12909;
wire      [7:0] n1291;
wire            n12910;
wire            n12911;
wire            n12912;
wire            n12913;
wire      [7:0] n12914;
wire            n12915;
wire            n12916;
wire            n12917;
wire            n12918;
wire            n12919;
wire      [7:0] n1292;
wire      [7:0] n12920;
wire            n12921;
wire            n12922;
wire            n12923;
wire            n12924;
wire            n12925;
wire      [7:0] n12926;
wire            n12927;
wire            n12928;
wire            n12929;
wire      [7:0] n1293;
wire            n12930;
wire            n12931;
wire      [7:0] n12932;
wire            n12933;
wire            n12934;
wire            n12935;
wire            n12936;
wire            n12937;
wire      [7:0] n12938;
wire            n12939;
wire      [7:0] n1294;
wire            n12940;
wire            n12941;
wire            n12942;
wire            n12943;
wire      [7:0] n12944;
wire            n12945;
wire            n12946;
wire            n12947;
wire            n12948;
wire            n12949;
wire      [7:0] n1295;
wire      [7:0] n12950;
wire            n12951;
wire            n12952;
wire            n12953;
wire            n12954;
wire            n12955;
wire      [7:0] n12956;
wire            n12957;
wire            n12958;
wire            n12959;
wire      [7:0] n1296;
wire            n12960;
wire            n12961;
wire      [7:0] n12962;
wire            n12963;
wire            n12964;
wire            n12965;
wire            n12966;
wire            n12967;
wire      [7:0] n12968;
wire            n12969;
wire      [7:0] n1297;
wire            n12970;
wire            n12971;
wire            n12972;
wire            n12973;
wire      [7:0] n12974;
wire            n12975;
wire            n12976;
wire            n12977;
wire            n12978;
wire            n12979;
wire      [7:0] n1298;
wire      [7:0] n12980;
wire            n12981;
wire            n12982;
wire            n12983;
wire            n12984;
wire            n12985;
wire      [7:0] n12986;
wire            n12987;
wire            n12988;
wire            n12989;
wire      [7:0] n1299;
wire            n12990;
wire            n12991;
wire      [7:0] n12992;
wire            n12993;
wire            n12994;
wire            n12995;
wire            n12996;
wire            n12997;
wire      [7:0] n12998;
wire            n12999;
wire            n13;
wire            n130;
wire      [7:0] n1300;
wire            n13000;
wire            n13001;
wire            n13002;
wire            n13003;
wire      [7:0] n13004;
wire            n13005;
wire            n13006;
wire            n13007;
wire            n13008;
wire            n13009;
wire      [7:0] n1301;
wire      [7:0] n13010;
wire            n13011;
wire            n13012;
wire            n13013;
wire            n13014;
wire            n13015;
wire      [7:0] n13016;
wire            n13017;
wire            n13018;
wire            n13019;
wire      [7:0] n1302;
wire            n13020;
wire            n13021;
wire      [7:0] n13022;
wire            n13023;
wire            n13024;
wire            n13025;
wire            n13026;
wire            n13027;
wire      [7:0] n13028;
wire            n13029;
wire      [7:0] n1303;
wire            n13030;
wire            n13031;
wire            n13032;
wire            n13033;
wire      [7:0] n13034;
wire            n13035;
wire            n13036;
wire            n13037;
wire            n13038;
wire            n13039;
wire      [7:0] n1304;
wire      [7:0] n13040;
wire            n13041;
wire            n13042;
wire            n13043;
wire            n13044;
wire            n13045;
wire      [7:0] n13046;
wire            n13047;
wire            n13048;
wire            n13049;
wire      [7:0] n1305;
wire            n13050;
wire            n13051;
wire      [7:0] n13052;
wire            n13053;
wire            n13054;
wire            n13055;
wire            n13056;
wire            n13057;
wire      [7:0] n13058;
wire            n13059;
wire      [7:0] n1306;
wire            n13060;
wire            n13061;
wire            n13062;
wire            n13063;
wire      [7:0] n13064;
wire            n13065;
wire            n13066;
wire            n13067;
wire            n13068;
wire            n13069;
wire      [7:0] n1307;
wire      [7:0] n13070;
wire            n13071;
wire            n13072;
wire            n13073;
wire            n13074;
wire            n13075;
wire      [7:0] n13076;
wire            n13077;
wire            n13078;
wire            n13079;
wire      [7:0] n1308;
wire            n13080;
wire            n13081;
wire      [7:0] n13082;
wire            n13083;
wire            n13084;
wire            n13085;
wire            n13086;
wire            n13087;
wire      [7:0] n13088;
wire            n13089;
wire      [7:0] n1309;
wire            n13090;
wire            n13091;
wire            n13092;
wire            n13093;
wire      [7:0] n13094;
wire            n13095;
wire            n13096;
wire            n13097;
wire            n13098;
wire            n13099;
wire      [7:0] n1310;
wire      [7:0] n13100;
wire            n13101;
wire            n13102;
wire            n13103;
wire            n13104;
wire            n13105;
wire      [7:0] n13106;
wire            n13107;
wire            n13108;
wire            n13109;
wire      [7:0] n1311;
wire            n13110;
wire            n13111;
wire      [7:0] n13112;
wire            n13113;
wire            n13114;
wire            n13115;
wire            n13116;
wire            n13117;
wire      [7:0] n13118;
wire            n13119;
wire      [7:0] n1312;
wire            n13120;
wire            n13121;
wire            n13122;
wire            n13123;
wire      [7:0] n13124;
wire            n13125;
wire            n13126;
wire            n13127;
wire            n13128;
wire            n13129;
wire      [7:0] n1313;
wire      [7:0] n13130;
wire            n13131;
wire            n13132;
wire            n13133;
wire            n13134;
wire            n13135;
wire      [7:0] n13136;
wire            n13137;
wire            n13138;
wire            n13139;
wire      [7:0] n1314;
wire            n13140;
wire            n13141;
wire      [7:0] n13142;
wire            n13143;
wire            n13144;
wire            n13145;
wire            n13146;
wire            n13147;
wire      [7:0] n13148;
wire            n13149;
wire      [7:0] n1315;
wire            n13150;
wire            n13151;
wire            n13152;
wire            n13153;
wire      [7:0] n13154;
wire            n13155;
wire            n13156;
wire            n13157;
wire            n13158;
wire            n13159;
wire      [7:0] n1316;
wire      [7:0] n13160;
wire            n13161;
wire            n13162;
wire            n13163;
wire            n13164;
wire            n13165;
wire      [7:0] n13166;
wire            n13167;
wire            n13168;
wire            n13169;
wire      [7:0] n1317;
wire            n13170;
wire            n13171;
wire      [7:0] n13172;
wire            n13173;
wire            n13174;
wire            n13175;
wire            n13176;
wire            n13177;
wire      [7:0] n13178;
wire            n13179;
wire      [7:0] n1318;
wire            n13180;
wire            n13181;
wire            n13182;
wire            n13183;
wire      [7:0] n13184;
wire            n13185;
wire            n13186;
wire            n13187;
wire            n13188;
wire            n13189;
wire      [7:0] n1319;
wire      [7:0] n13190;
wire            n13191;
wire            n13192;
wire            n13193;
wire            n13194;
wire            n13195;
wire      [7:0] n13196;
wire            n13197;
wire            n13198;
wire            n13199;
wire            n132;
wire      [7:0] n1320;
wire            n13200;
wire            n13201;
wire      [7:0] n13202;
wire            n13203;
wire            n13204;
wire            n13205;
wire            n13206;
wire            n13207;
wire      [7:0] n13208;
wire            n13209;
wire      [7:0] n1321;
wire            n13210;
wire            n13211;
wire            n13212;
wire            n13213;
wire      [7:0] n13214;
wire            n13215;
wire            n13216;
wire            n13217;
wire            n13218;
wire            n13219;
wire      [7:0] n1322;
wire      [7:0] n13220;
wire            n13221;
wire            n13222;
wire            n13223;
wire            n13224;
wire            n13225;
wire      [7:0] n13226;
wire            n13227;
wire            n13228;
wire            n13229;
wire      [7:0] n1323;
wire            n13230;
wire            n13231;
wire      [7:0] n13232;
wire            n13233;
wire            n13234;
wire            n13235;
wire            n13236;
wire            n13237;
wire      [7:0] n13238;
wire            n13239;
wire      [7:0] n1324;
wire            n13240;
wire            n13241;
wire            n13242;
wire            n13243;
wire      [7:0] n13244;
wire            n13245;
wire            n13246;
wire            n13247;
wire            n13248;
wire            n13249;
wire      [7:0] n1325;
wire      [7:0] n13250;
wire            n13251;
wire            n13252;
wire            n13253;
wire            n13254;
wire            n13255;
wire      [7:0] n13256;
wire            n13257;
wire            n13258;
wire            n13259;
wire      [7:0] n1326;
wire            n13260;
wire            n13261;
wire      [7:0] n13262;
wire            n13263;
wire            n13264;
wire            n13265;
wire            n13266;
wire            n13267;
wire      [7:0] n13268;
wire            n13269;
wire      [7:0] n1327;
wire            n13270;
wire            n13271;
wire            n13272;
wire            n13273;
wire      [7:0] n13274;
wire            n13275;
wire            n13276;
wire            n13277;
wire            n13278;
wire            n13279;
wire      [7:0] n1328;
wire      [7:0] n13280;
wire            n13281;
wire            n13282;
wire            n13283;
wire            n13284;
wire            n13285;
wire      [7:0] n13286;
wire            n13287;
wire            n13288;
wire            n13289;
wire      [7:0] n1329;
wire            n13290;
wire            n13291;
wire      [7:0] n13292;
wire            n13293;
wire            n13294;
wire            n13295;
wire            n13296;
wire            n13297;
wire      [7:0] n13298;
wire            n13299;
wire      [7:0] n1330;
wire            n13300;
wire            n13301;
wire            n13302;
wire            n13303;
wire      [7:0] n13304;
wire            n13305;
wire            n13306;
wire            n13307;
wire            n13308;
wire            n13309;
wire      [7:0] n1331;
wire      [7:0] n13310;
wire            n13311;
wire            n13312;
wire            n13313;
wire            n13314;
wire            n13315;
wire      [7:0] n13316;
wire            n13317;
wire            n13318;
wire            n13319;
wire      [7:0] n1332;
wire            n13320;
wire            n13321;
wire      [7:0] n13322;
wire            n13323;
wire            n13324;
wire            n13325;
wire            n13326;
wire            n13327;
wire      [7:0] n13328;
wire            n13329;
wire      [7:0] n1333;
wire            n13330;
wire            n13331;
wire            n13332;
wire            n13333;
wire      [7:0] n13334;
wire            n13335;
wire            n13336;
wire            n13337;
wire            n13338;
wire            n13339;
wire      [7:0] n1334;
wire      [7:0] n13340;
wire            n13341;
wire            n13342;
wire            n13343;
wire            n13344;
wire            n13345;
wire      [7:0] n13346;
wire            n13347;
wire            n13348;
wire            n13349;
wire      [7:0] n1335;
wire            n13350;
wire            n13351;
wire      [7:0] n13352;
wire            n13353;
wire            n13354;
wire            n13355;
wire            n13356;
wire            n13357;
wire      [7:0] n13358;
wire            n13359;
wire      [7:0] n1336;
wire            n13360;
wire            n13361;
wire            n13362;
wire            n13363;
wire      [7:0] n13364;
wire            n13365;
wire            n13366;
wire            n13367;
wire            n13368;
wire            n13369;
wire      [7:0] n1337;
wire      [7:0] n13370;
wire            n13371;
wire            n13372;
wire            n13373;
wire            n13374;
wire            n13375;
wire      [7:0] n13376;
wire            n13377;
wire            n13378;
wire            n13379;
wire      [7:0] n1338;
wire            n13380;
wire            n13381;
wire      [7:0] n13382;
wire            n13383;
wire            n13384;
wire            n13385;
wire            n13386;
wire            n13387;
wire      [7:0] n13388;
wire            n13389;
wire      [7:0] n1339;
wire            n13390;
wire            n13391;
wire            n13392;
wire            n13393;
wire      [7:0] n13394;
wire            n13395;
wire            n13396;
wire            n13397;
wire            n13398;
wire            n13399;
wire            n134;
wire      [7:0] n1340;
wire      [7:0] n13400;
wire            n13401;
wire            n13402;
wire            n13403;
wire            n13404;
wire            n13405;
wire      [7:0] n13406;
wire            n13407;
wire            n13408;
wire            n13409;
wire      [7:0] n1341;
wire            n13410;
wire            n13411;
wire      [7:0] n13412;
wire            n13413;
wire            n13414;
wire            n13415;
wire            n13416;
wire            n13417;
wire      [7:0] n13418;
wire            n13419;
wire      [7:0] n1342;
wire            n13420;
wire            n13421;
wire            n13422;
wire            n13423;
wire      [7:0] n13424;
wire            n13425;
wire            n13426;
wire            n13427;
wire            n13428;
wire            n13429;
wire      [7:0] n1343;
wire      [7:0] n13430;
wire            n13431;
wire            n13432;
wire            n13433;
wire            n13434;
wire            n13435;
wire      [7:0] n13436;
wire            n13437;
wire            n13438;
wire            n13439;
wire      [7:0] n1344;
wire            n13440;
wire            n13441;
wire      [7:0] n13442;
wire            n13443;
wire            n13444;
wire            n13445;
wire            n13446;
wire            n13447;
wire      [7:0] n13448;
wire            n13449;
wire            n1345;
wire            n13450;
wire            n13451;
wire            n13452;
wire            n13453;
wire      [7:0] n13454;
wire            n13455;
wire            n13456;
wire            n13457;
wire            n13458;
wire            n13459;
wire            n1346;
wire      [7:0] n13460;
wire            n13461;
wire            n13462;
wire            n13463;
wire            n13464;
wire            n13465;
wire      [7:0] n13466;
wire            n13467;
wire            n13468;
wire            n13469;
wire      [3:0] n1347;
wire            n13470;
wire            n13471;
wire      [7:0] n13472;
wire            n13473;
wire            n13474;
wire            n13475;
wire            n13476;
wire            n13477;
wire      [7:0] n13478;
wire            n13479;
wire      [4:0] n1348;
wire            n13480;
wire            n13481;
wire            n13482;
wire            n13483;
wire      [7:0] n13484;
wire            n13485;
wire            n13486;
wire            n13487;
wire            n13488;
wire            n13489;
wire      [7:0] n1349;
wire      [7:0] n13490;
wire            n13491;
wire            n13492;
wire            n13493;
wire            n13494;
wire            n13495;
wire      [7:0] n13496;
wire            n13497;
wire            n13498;
wire            n13499;
wire      [3:0] n1350;
wire            n13500;
wire            n13501;
wire      [7:0] n13502;
wire            n13503;
wire            n13504;
wire            n13505;
wire            n13506;
wire            n13507;
wire      [7:0] n13508;
wire            n13509;
wire      [7:0] n1351;
wire            n13510;
wire            n13511;
wire            n13512;
wire            n13513;
wire      [7:0] n13514;
wire            n13515;
wire            n13516;
wire            n13517;
wire            n13518;
wire            n13519;
wire      [7:0] n1352;
wire      [7:0] n13520;
wire            n13521;
wire            n13522;
wire            n13523;
wire            n13524;
wire            n13525;
wire      [7:0] n13526;
wire            n13527;
wire            n13528;
wire            n13529;
wire      [7:0] n1353;
wire            n13530;
wire            n13531;
wire      [7:0] n13532;
wire            n13533;
wire            n13534;
wire            n13535;
wire            n13536;
wire            n13537;
wire      [7:0] n13538;
wire            n13539;
wire      [7:0] n1354;
wire            n13540;
wire            n13541;
wire            n13542;
wire            n13543;
wire      [7:0] n13544;
wire            n13545;
wire            n13546;
wire            n13547;
wire            n13548;
wire            n13549;
wire            n1355;
wire      [7:0] n13550;
wire            n13551;
wire            n13552;
wire            n13553;
wire            n13554;
wire            n13555;
wire      [7:0] n13556;
wire            n13557;
wire            n13558;
wire            n13559;
wire            n1356;
wire            n13560;
wire            n13561;
wire      [7:0] n13562;
wire            n13563;
wire            n13564;
wire            n13565;
wire            n13566;
wire            n13567;
wire      [7:0] n13568;
wire            n13569;
wire            n1357;
wire            n13570;
wire            n13571;
wire            n13572;
wire            n13573;
wire      [7:0] n13574;
wire            n13575;
wire            n13576;
wire            n13577;
wire            n13578;
wire            n13579;
wire            n1358;
wire      [7:0] n13580;
wire            n13581;
wire            n13582;
wire            n13583;
wire            n13584;
wire            n13585;
wire      [7:0] n13586;
wire            n13587;
wire            n13588;
wire            n13589;
wire            n1359;
wire            n13590;
wire            n13591;
wire      [7:0] n13592;
wire            n13593;
wire            n13594;
wire            n13595;
wire            n13596;
wire            n13597;
wire      [7:0] n13598;
wire            n13599;
wire            n136;
wire            n1360;
wire            n13600;
wire            n13601;
wire            n13602;
wire            n13603;
wire      [7:0] n13604;
wire            n13605;
wire            n13606;
wire            n13607;
wire            n13608;
wire            n13609;
wire            n1361;
wire      [7:0] n13610;
wire            n13611;
wire            n13612;
wire            n13613;
wire            n13614;
wire            n13615;
wire      [7:0] n13616;
wire            n13617;
wire            n13618;
wire            n13619;
wire            n1362;
wire            n13620;
wire            n13621;
wire      [7:0] n13622;
wire            n13623;
wire            n13624;
wire            n13625;
wire            n13626;
wire            n13627;
wire      [7:0] n13628;
wire            n13629;
wire            n1363;
wire            n13630;
wire            n13631;
wire            n13632;
wire            n13633;
wire      [7:0] n13634;
wire            n13635;
wire            n13636;
wire            n13637;
wire            n13638;
wire            n13639;
wire            n1364;
wire      [7:0] n13640;
wire            n13641;
wire            n13642;
wire            n13643;
wire            n13644;
wire            n13645;
wire      [7:0] n13646;
wire            n13647;
wire            n13648;
wire            n13649;
wire            n1365;
wire            n13650;
wire            n13651;
wire      [7:0] n13652;
wire            n13653;
wire            n13654;
wire            n13655;
wire            n13656;
wire            n13657;
wire      [7:0] n13658;
wire            n13659;
wire            n1366;
wire            n13660;
wire            n13661;
wire            n13662;
wire            n13663;
wire      [7:0] n13664;
wire            n13665;
wire            n13666;
wire            n13667;
wire            n13668;
wire            n13669;
wire            n1367;
wire      [7:0] n13670;
wire            n13671;
wire            n13672;
wire            n13673;
wire            n13674;
wire            n13675;
wire      [7:0] n13676;
wire            n13677;
wire            n13678;
wire            n13679;
wire            n1368;
wire            n13680;
wire            n13681;
wire      [7:0] n13682;
wire            n13683;
wire            n13684;
wire            n13685;
wire            n13686;
wire            n13687;
wire      [7:0] n13688;
wire            n13689;
wire            n1369;
wire            n13690;
wire            n13691;
wire            n13692;
wire            n13693;
wire      [7:0] n13694;
wire            n13695;
wire            n13696;
wire            n13697;
wire            n13698;
wire            n13699;
wire            n1370;
wire      [7:0] n13700;
wire            n13701;
wire            n13702;
wire            n13703;
wire            n13704;
wire            n13705;
wire      [7:0] n13706;
wire            n13707;
wire            n13708;
wire            n13709;
wire            n1371;
wire            n13710;
wire            n13711;
wire      [7:0] n13712;
wire            n13713;
wire            n13714;
wire            n13715;
wire            n13716;
wire            n13717;
wire      [7:0] n13718;
wire            n13719;
wire            n1372;
wire            n13720;
wire            n13721;
wire            n13722;
wire            n13723;
wire      [7:0] n13724;
wire            n13725;
wire            n13726;
wire            n13727;
wire            n13728;
wire            n13729;
wire            n1373;
wire      [7:0] n13730;
wire            n13731;
wire            n13732;
wire            n13733;
wire            n13734;
wire            n13735;
wire      [7:0] n13736;
wire            n13737;
wire            n13738;
wire            n13739;
wire            n1374;
wire            n13740;
wire            n13741;
wire      [7:0] n13742;
wire            n13743;
wire            n13744;
wire            n13745;
wire            n13746;
wire            n13747;
wire      [7:0] n13748;
wire            n13749;
wire            n1375;
wire            n13750;
wire            n13751;
wire            n13752;
wire            n13753;
wire      [7:0] n13754;
wire            n13755;
wire            n13756;
wire            n13757;
wire            n13758;
wire            n13759;
wire            n1376;
wire      [7:0] n13760;
wire            n13761;
wire            n13762;
wire            n13763;
wire            n13764;
wire            n13765;
wire      [7:0] n13766;
wire            n13767;
wire            n13768;
wire            n13769;
wire            n1377;
wire            n13770;
wire            n13771;
wire      [7:0] n13772;
wire            n13773;
wire            n13774;
wire            n13775;
wire            n13776;
wire            n13777;
wire      [7:0] n13778;
wire            n13779;
wire            n1378;
wire            n13780;
wire            n13781;
wire            n13782;
wire            n13783;
wire      [7:0] n13784;
wire            n13785;
wire            n13786;
wire            n13787;
wire            n13788;
wire            n13789;
wire            n1379;
wire      [7:0] n13790;
wire            n13791;
wire            n13792;
wire            n13793;
wire            n13794;
wire            n13795;
wire      [7:0] n13796;
wire            n13797;
wire            n13798;
wire            n13799;
wire            n138;
wire            n1380;
wire            n13800;
wire            n13801;
wire      [7:0] n13802;
wire            n13803;
wire            n13804;
wire            n13805;
wire            n13806;
wire            n13807;
wire      [7:0] n13808;
wire            n13809;
wire            n1381;
wire            n13810;
wire            n13811;
wire            n13812;
wire            n13813;
wire      [7:0] n13814;
wire            n13815;
wire            n13816;
wire            n13817;
wire            n13818;
wire            n13819;
wire            n1382;
wire      [7:0] n13820;
wire            n13821;
wire            n13822;
wire            n13823;
wire            n13824;
wire            n13825;
wire      [7:0] n13826;
wire            n13827;
wire            n13828;
wire            n13829;
wire            n1383;
wire            n13830;
wire            n13831;
wire      [7:0] n13832;
wire            n13833;
wire            n13834;
wire            n13835;
wire            n13836;
wire            n13837;
wire      [7:0] n13838;
wire            n13839;
wire            n1384;
wire            n13840;
wire            n13841;
wire            n13842;
wire            n13843;
wire      [7:0] n13844;
wire            n13845;
wire            n13846;
wire            n13847;
wire            n13848;
wire            n13849;
wire            n1385;
wire      [7:0] n13850;
wire            n13851;
wire            n13852;
wire            n13853;
wire            n13854;
wire            n13855;
wire      [7:0] n13856;
wire            n13857;
wire            n13858;
wire            n13859;
wire            n1386;
wire            n13860;
wire            n13861;
wire      [7:0] n13862;
wire            n13863;
wire            n13864;
wire            n13865;
wire            n13866;
wire            n13867;
wire      [7:0] n13868;
wire            n13869;
wire            n1387;
wire            n13870;
wire            n13871;
wire            n13872;
wire            n13873;
wire      [7:0] n13874;
wire            n13875;
wire            n13876;
wire            n13877;
wire            n13878;
wire            n13879;
wire            n1388;
wire      [7:0] n13880;
wire            n13881;
wire            n13882;
wire            n13883;
wire            n13884;
wire            n13885;
wire      [7:0] n13886;
wire            n13887;
wire            n13888;
wire            n13889;
wire            n1389;
wire            n13890;
wire            n13891;
wire      [7:0] n13892;
wire            n13893;
wire            n13894;
wire            n13895;
wire            n13896;
wire            n13897;
wire      [7:0] n13898;
wire            n13899;
wire            n1390;
wire            n13900;
wire            n13901;
wire            n13902;
wire            n13903;
wire      [7:0] n13904;
wire            n13905;
wire            n13906;
wire            n13907;
wire            n13908;
wire            n13909;
wire            n1391;
wire      [7:0] n13910;
wire            n13911;
wire            n13912;
wire            n13913;
wire            n13914;
wire            n13915;
wire      [7:0] n13916;
wire            n13917;
wire            n13918;
wire            n13919;
wire            n1392;
wire            n13920;
wire            n13921;
wire      [7:0] n13922;
wire            n13923;
wire            n13924;
wire            n13925;
wire            n13926;
wire            n13927;
wire      [7:0] n13928;
wire            n13929;
wire            n1393;
wire            n13930;
wire            n13931;
wire            n13932;
wire            n13933;
wire      [7:0] n13934;
wire            n13935;
wire            n13936;
wire            n13937;
wire            n13938;
wire            n13939;
wire            n1394;
wire      [7:0] n13940;
wire            n13941;
wire            n13942;
wire            n13943;
wire            n13944;
wire            n13945;
wire      [7:0] n13946;
wire            n13947;
wire            n13948;
wire            n13949;
wire            n1395;
wire            n13950;
wire            n13951;
wire      [7:0] n13952;
wire            n13953;
wire            n13954;
wire            n13955;
wire            n13956;
wire            n13957;
wire      [7:0] n13958;
wire            n13959;
wire            n1396;
wire            n13960;
wire            n13961;
wire            n13962;
wire            n13963;
wire      [7:0] n13964;
wire            n13965;
wire            n13966;
wire            n13967;
wire            n13968;
wire            n13969;
wire            n1397;
wire      [7:0] n13970;
wire            n13971;
wire            n13972;
wire            n13973;
wire            n13974;
wire            n13975;
wire      [7:0] n13976;
wire            n13977;
wire            n13978;
wire            n13979;
wire            n1398;
wire            n13980;
wire            n13981;
wire      [7:0] n13982;
wire            n13983;
wire            n13984;
wire            n13985;
wire            n13986;
wire            n13987;
wire      [7:0] n13988;
wire            n13989;
wire            n1399;
wire            n13990;
wire            n13991;
wire            n13992;
wire            n13993;
wire      [7:0] n13994;
wire            n13995;
wire            n13996;
wire            n13997;
wire            n13998;
wire            n13999;
wire            n140;
wire            n1400;
wire      [7:0] n14000;
wire            n14001;
wire            n14002;
wire            n14003;
wire            n14004;
wire            n14005;
wire      [7:0] n14006;
wire            n14007;
wire            n14008;
wire            n14009;
wire            n1401;
wire            n14010;
wire            n14011;
wire      [7:0] n14012;
wire            n14013;
wire            n14014;
wire            n14015;
wire            n14016;
wire            n14017;
wire      [7:0] n14018;
wire            n14019;
wire            n1402;
wire            n14020;
wire            n14021;
wire            n14022;
wire            n14023;
wire      [7:0] n14024;
wire            n14025;
wire            n14026;
wire            n14027;
wire            n14028;
wire            n14029;
wire            n1403;
wire      [7:0] n14030;
wire            n14031;
wire            n14032;
wire            n14033;
wire            n14034;
wire            n14035;
wire      [7:0] n14036;
wire            n14037;
wire            n14038;
wire            n14039;
wire            n1404;
wire            n14040;
wire            n14041;
wire      [7:0] n14042;
wire            n14043;
wire            n14044;
wire            n14045;
wire            n14046;
wire            n14047;
wire      [7:0] n14048;
wire            n14049;
wire            n1405;
wire            n14050;
wire            n14051;
wire            n14052;
wire            n14053;
wire      [7:0] n14054;
wire            n14055;
wire            n14056;
wire            n14057;
wire            n14058;
wire            n14059;
wire            n1406;
wire      [7:0] n14060;
wire            n14061;
wire            n14062;
wire            n14063;
wire            n14064;
wire            n14065;
wire      [7:0] n14066;
wire            n14067;
wire            n14068;
wire            n14069;
wire            n1407;
wire            n14070;
wire            n14071;
wire      [7:0] n14072;
wire            n14073;
wire            n14074;
wire            n14075;
wire            n14076;
wire            n14077;
wire      [7:0] n14078;
wire            n14079;
wire            n1408;
wire            n14080;
wire            n14081;
wire            n14082;
wire            n14083;
wire      [7:0] n14084;
wire            n14085;
wire            n14086;
wire            n14087;
wire            n14088;
wire            n14089;
wire            n1409;
wire      [7:0] n14090;
wire            n14091;
wire            n14092;
wire            n14093;
wire            n14094;
wire            n14095;
wire      [7:0] n14096;
wire            n14097;
wire            n14098;
wire            n14099;
wire            n1410;
wire            n14100;
wire            n14101;
wire      [7:0] n14102;
wire            n14103;
wire            n14104;
wire            n14105;
wire            n14106;
wire            n14107;
wire      [7:0] n14108;
wire            n14109;
wire            n1411;
wire            n14110;
wire            n14111;
wire            n14112;
wire            n14113;
wire      [7:0] n14114;
wire            n14115;
wire            n14116;
wire            n14117;
wire            n14118;
wire            n14119;
wire            n1412;
wire      [7:0] n14120;
wire            n14121;
wire            n14122;
wire            n14123;
wire            n14124;
wire            n14125;
wire      [7:0] n14126;
wire            n14127;
wire            n14128;
wire            n14129;
wire            n1413;
wire            n14130;
wire            n14131;
wire      [7:0] n14132;
wire            n14133;
wire            n14134;
wire            n14135;
wire            n14136;
wire            n14137;
wire      [7:0] n14138;
wire            n14139;
wire            n1414;
wire            n14140;
wire            n14141;
wire            n14142;
wire            n14143;
wire      [7:0] n14144;
wire            n14145;
wire            n14146;
wire            n14147;
wire            n14148;
wire            n14149;
wire            n1415;
wire      [7:0] n14150;
wire            n14151;
wire            n14152;
wire            n14153;
wire            n14154;
wire            n14155;
wire      [7:0] n14156;
wire            n14157;
wire            n14158;
wire            n14159;
wire            n1416;
wire            n14160;
wire            n14161;
wire      [7:0] n14162;
wire            n14163;
wire            n14164;
wire            n14165;
wire            n14166;
wire            n14167;
wire      [7:0] n14168;
wire            n14169;
wire            n1417;
wire            n14170;
wire            n14171;
wire            n14172;
wire            n14173;
wire      [7:0] n14174;
wire            n14175;
wire            n14176;
wire            n14177;
wire            n14178;
wire            n14179;
wire            n1418;
wire      [7:0] n14180;
wire            n14181;
wire            n14182;
wire            n14183;
wire            n14184;
wire            n14185;
wire      [7:0] n14186;
wire            n14187;
wire            n14188;
wire            n14189;
wire            n1419;
wire            n14190;
wire            n14191;
wire      [7:0] n14192;
wire            n14193;
wire            n14194;
wire            n14195;
wire            n14196;
wire            n14197;
wire      [7:0] n14198;
wire            n14199;
wire            n142;
wire            n1420;
wire            n14200;
wire            n14201;
wire            n14202;
wire            n14203;
wire      [7:0] n14204;
wire            n14205;
wire            n14206;
wire            n14207;
wire            n14208;
wire            n14209;
wire            n1421;
wire      [7:0] n14210;
wire            n14211;
wire            n14212;
wire            n14213;
wire            n14214;
wire            n14215;
wire      [7:0] n14216;
wire            n14217;
wire            n14218;
wire            n14219;
wire            n1422;
wire            n14220;
wire            n14221;
wire      [7:0] n14222;
wire            n14223;
wire            n14224;
wire            n14225;
wire            n14226;
wire            n14227;
wire      [7:0] n14228;
wire            n14229;
wire            n1423;
wire            n14230;
wire            n14231;
wire            n14232;
wire            n14233;
wire      [7:0] n14234;
wire            n14235;
wire            n14236;
wire            n14237;
wire            n14238;
wire            n14239;
wire            n1424;
wire      [7:0] n14240;
wire            n14241;
wire            n14242;
wire            n14243;
wire            n14244;
wire            n14245;
wire      [7:0] n14246;
wire            n14247;
wire            n14248;
wire            n14249;
wire            n1425;
wire            n14250;
wire            n14251;
wire      [7:0] n14252;
wire            n14253;
wire            n14254;
wire            n14255;
wire            n14256;
wire            n14257;
wire      [7:0] n14258;
wire            n14259;
wire            n1426;
wire            n14260;
wire            n14261;
wire            n14262;
wire            n14263;
wire      [7:0] n14264;
wire            n14265;
wire            n14266;
wire            n14267;
wire            n14268;
wire            n14269;
wire            n1427;
wire      [7:0] n14270;
wire            n14271;
wire            n14272;
wire            n14273;
wire            n14274;
wire            n14275;
wire      [7:0] n14276;
wire            n14277;
wire            n14278;
wire            n14279;
wire            n1428;
wire            n14280;
wire            n14281;
wire      [7:0] n14282;
wire            n14283;
wire            n14284;
wire            n14285;
wire            n14286;
wire            n14287;
wire      [7:0] n14288;
wire            n14289;
wire            n1429;
wire            n14290;
wire            n14291;
wire            n14292;
wire            n14293;
wire      [7:0] n14294;
wire            n14295;
wire            n14296;
wire            n14297;
wire            n14298;
wire            n14299;
wire            n1430;
wire      [7:0] n14300;
wire            n14301;
wire            n14302;
wire            n14303;
wire            n14304;
wire            n14305;
wire      [7:0] n14306;
wire            n14307;
wire            n14308;
wire            n14309;
wire            n1431;
wire            n14310;
wire            n14311;
wire      [7:0] n14312;
wire            n14313;
wire            n14314;
wire            n14315;
wire            n14316;
wire            n14317;
wire      [7:0] n14318;
wire            n14319;
wire            n1432;
wire            n14320;
wire            n14321;
wire            n14322;
wire            n14323;
wire      [7:0] n14324;
wire            n14325;
wire            n14326;
wire            n14327;
wire            n14328;
wire            n14329;
wire            n1433;
wire      [7:0] n14330;
wire            n14331;
wire            n14332;
wire            n14333;
wire            n14334;
wire            n14335;
wire      [7:0] n14336;
wire            n14337;
wire            n14338;
wire            n14339;
wire            n1434;
wire            n14340;
wire            n14341;
wire      [7:0] n14342;
wire            n14343;
wire            n14344;
wire            n14345;
wire            n14346;
wire            n14347;
wire      [7:0] n14348;
wire            n14349;
wire            n1435;
wire            n14350;
wire            n14351;
wire            n14352;
wire            n14353;
wire      [7:0] n14354;
wire            n14355;
wire            n14356;
wire            n14357;
wire            n14358;
wire            n14359;
wire            n1436;
wire      [7:0] n14360;
wire            n14361;
wire            n14362;
wire            n14363;
wire            n14364;
wire            n14365;
wire      [7:0] n14366;
wire            n14367;
wire            n14368;
wire            n14369;
wire            n1437;
wire            n14370;
wire            n14371;
wire      [7:0] n14372;
wire            n14373;
wire            n14374;
wire            n14375;
wire            n14376;
wire            n14377;
wire      [7:0] n14378;
wire            n14379;
wire            n1438;
wire            n14380;
wire            n14381;
wire            n14382;
wire            n14383;
wire      [7:0] n14384;
wire            n14385;
wire            n14386;
wire            n14387;
wire            n14388;
wire            n14389;
wire            n1439;
wire      [7:0] n14390;
wire            n14391;
wire            n14392;
wire            n14393;
wire            n14394;
wire            n14395;
wire      [7:0] n14396;
wire            n14397;
wire            n14398;
wire            n14399;
wire            n144;
wire            n1440;
wire            n14400;
wire            n14401;
wire      [7:0] n14402;
wire            n14403;
wire            n14404;
wire            n14405;
wire            n14406;
wire            n14407;
wire      [7:0] n14408;
wire            n14409;
wire            n1441;
wire            n14410;
wire            n14411;
wire            n14412;
wire            n14413;
wire      [7:0] n14414;
wire            n14415;
wire            n14416;
wire            n14417;
wire            n14418;
wire            n14419;
wire            n1442;
wire      [7:0] n14420;
wire            n14421;
wire            n14422;
wire            n14423;
wire            n14424;
wire            n14425;
wire      [7:0] n14426;
wire            n14427;
wire            n14428;
wire            n14429;
wire            n1443;
wire            n14430;
wire            n14431;
wire      [7:0] n14432;
wire            n14433;
wire            n14434;
wire            n14435;
wire            n14436;
wire            n14437;
wire      [7:0] n14438;
wire            n14439;
wire            n1444;
wire            n14440;
wire            n14441;
wire            n14442;
wire            n14443;
wire      [7:0] n14444;
wire            n14445;
wire            n14446;
wire            n14447;
wire            n14448;
wire            n14449;
wire            n1445;
wire      [7:0] n14450;
wire            n14451;
wire            n14452;
wire            n14453;
wire            n14454;
wire            n14455;
wire      [7:0] n14456;
wire            n14457;
wire            n14458;
wire            n14459;
wire            n1446;
wire            n14460;
wire            n14461;
wire      [7:0] n14462;
wire            n14463;
wire            n14464;
wire            n14465;
wire            n14466;
wire            n14467;
wire      [7:0] n14468;
wire            n14469;
wire            n1447;
wire            n14470;
wire            n14471;
wire            n14472;
wire            n14473;
wire      [7:0] n14474;
wire            n14475;
wire            n14476;
wire            n14477;
wire            n14478;
wire            n14479;
wire            n1448;
wire      [7:0] n14480;
wire            n14481;
wire            n14482;
wire            n14483;
wire            n14484;
wire            n14485;
wire      [7:0] n14486;
wire            n14487;
wire            n14488;
wire            n14489;
wire            n1449;
wire            n14490;
wire            n14491;
wire      [7:0] n14492;
wire            n14493;
wire            n14494;
wire            n14495;
wire            n14496;
wire            n14497;
wire      [7:0] n14498;
wire            n14499;
wire            n1450;
wire            n14500;
wire            n14501;
wire            n14502;
wire            n14503;
wire      [7:0] n14504;
wire            n14505;
wire            n14506;
wire            n14507;
wire            n14508;
wire            n14509;
wire            n1451;
wire      [7:0] n14510;
wire            n14511;
wire            n14512;
wire            n14513;
wire            n14514;
wire            n14515;
wire      [7:0] n14516;
wire            n14517;
wire            n14518;
wire            n14519;
wire            n1452;
wire            n14520;
wire            n14521;
wire      [7:0] n14522;
wire            n14523;
wire            n14524;
wire            n14525;
wire            n14526;
wire            n14527;
wire      [7:0] n14528;
wire            n14529;
wire            n1453;
wire            n14530;
wire            n14531;
wire            n14532;
wire            n14533;
wire      [7:0] n14534;
wire            n14535;
wire            n14536;
wire            n14537;
wire            n14538;
wire            n14539;
wire            n1454;
wire      [7:0] n14540;
wire            n14541;
wire            n14542;
wire            n14543;
wire            n14544;
wire            n14545;
wire      [7:0] n14546;
wire            n14547;
wire            n14548;
wire            n14549;
wire            n1455;
wire            n14550;
wire            n14551;
wire      [7:0] n14552;
wire            n14553;
wire            n14554;
wire            n14555;
wire            n14556;
wire            n14557;
wire      [7:0] n14558;
wire            n14559;
wire            n1456;
wire            n14560;
wire            n14561;
wire            n14562;
wire            n14563;
wire      [7:0] n14564;
wire            n14565;
wire            n14566;
wire            n14567;
wire            n14568;
wire            n14569;
wire            n1457;
wire      [7:0] n14570;
wire            n14571;
wire            n14572;
wire            n14573;
wire            n14574;
wire            n14575;
wire      [7:0] n14576;
wire            n14577;
wire            n14578;
wire            n14579;
wire            n1458;
wire            n14580;
wire            n14581;
wire      [7:0] n14582;
wire            n14583;
wire            n14584;
wire            n14585;
wire            n14586;
wire            n14587;
wire      [7:0] n14588;
wire            n14589;
wire            n1459;
wire            n14590;
wire            n14591;
wire            n14592;
wire            n14593;
wire      [7:0] n14594;
wire            n14595;
wire            n14596;
wire            n14597;
wire            n14598;
wire            n14599;
wire            n146;
wire            n1460;
wire      [7:0] n14600;
wire            n14601;
wire            n14602;
wire            n14603;
wire            n14604;
wire            n14605;
wire      [7:0] n14606;
wire            n14607;
wire            n14608;
wire            n14609;
wire            n1461;
wire            n14610;
wire            n14611;
wire      [7:0] n14612;
wire            n14613;
wire            n14614;
wire            n14615;
wire            n14616;
wire            n14617;
wire      [7:0] n14618;
wire            n14619;
wire            n1462;
wire            n14620;
wire            n14621;
wire            n14622;
wire            n14623;
wire      [7:0] n14624;
wire            n14625;
wire            n14626;
wire            n14627;
wire            n14628;
wire            n14629;
wire            n1463;
wire      [7:0] n14630;
wire            n14631;
wire            n14632;
wire            n14633;
wire            n14634;
wire            n14635;
wire      [7:0] n14636;
wire            n14637;
wire            n14638;
wire            n14639;
wire            n1464;
wire            n14640;
wire            n14641;
wire      [7:0] n14642;
wire            n14643;
wire            n14644;
wire            n14645;
wire            n14646;
wire            n14647;
wire      [7:0] n14648;
wire            n14649;
wire            n1465;
wire            n14650;
wire            n14651;
wire            n14652;
wire            n14653;
wire      [7:0] n14654;
wire            n14655;
wire            n14656;
wire            n14657;
wire            n14658;
wire            n14659;
wire            n1466;
wire      [7:0] n14660;
wire            n14661;
wire            n14662;
wire            n14663;
wire            n14664;
wire            n14665;
wire      [7:0] n14666;
wire            n14667;
wire            n14668;
wire            n14669;
wire            n1467;
wire            n14670;
wire            n14671;
wire      [7:0] n14672;
wire            n14673;
wire            n14674;
wire            n14675;
wire            n14676;
wire            n14677;
wire      [7:0] n14678;
wire            n14679;
wire            n1468;
wire            n14680;
wire            n14681;
wire            n14682;
wire            n14683;
wire      [7:0] n14684;
wire            n14685;
wire            n14686;
wire            n14687;
wire            n14688;
wire            n14689;
wire            n1469;
wire      [7:0] n14690;
wire            n14691;
wire            n14692;
wire            n14693;
wire            n14694;
wire            n14695;
wire      [7:0] n14696;
wire            n14697;
wire            n14698;
wire            n14699;
wire            n1470;
wire            n14700;
wire            n14701;
wire      [7:0] n14702;
wire            n14703;
wire            n14704;
wire            n14705;
wire            n14706;
wire            n14707;
wire      [7:0] n14708;
wire            n14709;
wire            n1471;
wire            n14710;
wire            n14711;
wire            n14712;
wire            n14713;
wire      [7:0] n14714;
wire            n14715;
wire            n14716;
wire            n14717;
wire            n14718;
wire            n14719;
wire            n1472;
wire      [7:0] n14720;
wire            n14721;
wire            n14722;
wire            n14723;
wire            n14724;
wire            n14725;
wire      [7:0] n14726;
wire            n14727;
wire            n14728;
wire            n14729;
wire            n1473;
wire            n14730;
wire            n14731;
wire      [7:0] n14732;
wire            n14733;
wire            n14734;
wire            n14735;
wire            n14736;
wire            n14737;
wire      [7:0] n14738;
wire            n14739;
wire            n1474;
wire            n14740;
wire            n14741;
wire            n14742;
wire            n14743;
wire      [7:0] n14744;
wire            n14745;
wire            n14746;
wire            n14747;
wire            n14748;
wire            n14749;
wire            n1475;
wire      [7:0] n14750;
wire            n14751;
wire            n14752;
wire            n14753;
wire            n14754;
wire            n14755;
wire      [7:0] n14756;
wire            n14757;
wire            n14758;
wire            n14759;
wire            n1476;
wire            n14760;
wire            n14761;
wire      [7:0] n14762;
wire            n14763;
wire            n14764;
wire            n14765;
wire            n14766;
wire            n14767;
wire      [7:0] n14768;
wire            n14769;
wire            n1477;
wire            n14770;
wire            n14771;
wire            n14772;
wire            n14773;
wire      [7:0] n14774;
wire            n14775;
wire            n14776;
wire            n14777;
wire            n14778;
wire            n14779;
wire            n1478;
wire      [7:0] n14780;
wire            n14781;
wire            n14782;
wire            n14783;
wire            n14784;
wire            n14785;
wire      [7:0] n14786;
wire            n14787;
wire            n14788;
wire            n14789;
wire            n1479;
wire            n14790;
wire            n14791;
wire      [7:0] n14792;
wire            n14793;
wire            n14794;
wire            n14795;
wire            n14796;
wire            n14797;
wire      [7:0] n14798;
wire            n14799;
wire            n148;
wire            n1480;
wire            n14800;
wire            n14801;
wire            n14802;
wire            n14803;
wire      [7:0] n14804;
wire            n14805;
wire            n14806;
wire            n14807;
wire            n14808;
wire            n14809;
wire            n1481;
wire      [7:0] n14810;
wire            n14811;
wire            n14812;
wire            n14813;
wire            n14814;
wire            n14815;
wire      [7:0] n14816;
wire            n14817;
wire            n14818;
wire            n14819;
wire            n1482;
wire            n14820;
wire            n14821;
wire      [7:0] n14822;
wire            n14823;
wire            n14824;
wire            n14825;
wire            n14826;
wire            n14827;
wire      [7:0] n14828;
wire            n14829;
wire            n1483;
wire            n14830;
wire            n14831;
wire            n14832;
wire            n14833;
wire      [7:0] n14834;
wire            n14835;
wire            n14836;
wire            n14837;
wire            n14838;
wire            n14839;
wire            n1484;
wire      [7:0] n14840;
wire            n14841;
wire            n14842;
wire            n14843;
wire            n14844;
wire            n14845;
wire      [7:0] n14846;
wire            n14847;
wire            n14848;
wire            n14849;
wire            n1485;
wire            n14850;
wire            n14851;
wire      [7:0] n14852;
wire            n14853;
wire            n14854;
wire            n14855;
wire            n14856;
wire            n14857;
wire      [7:0] n14858;
wire            n14859;
wire            n1486;
wire            n14860;
wire            n14861;
wire            n14862;
wire            n14863;
wire      [7:0] n14864;
wire            n14865;
wire            n14866;
wire            n14867;
wire            n14868;
wire            n14869;
wire            n1487;
wire      [7:0] n14870;
wire            n14871;
wire            n14872;
wire            n14873;
wire            n14874;
wire            n14875;
wire      [7:0] n14876;
wire            n14877;
wire            n14878;
wire            n14879;
wire            n1488;
wire            n14880;
wire            n14881;
wire      [7:0] n14882;
wire            n14883;
wire            n14884;
wire            n14885;
wire            n14886;
wire            n14887;
wire      [7:0] n14888;
wire            n14889;
wire            n1489;
wire            n14890;
wire            n14891;
wire            n14892;
wire            n14893;
wire      [7:0] n14894;
wire            n14895;
wire            n14896;
wire            n14897;
wire            n14898;
wire            n14899;
wire            n1490;
wire      [7:0] n14900;
wire            n14901;
wire            n14902;
wire            n14903;
wire            n14904;
wire            n14905;
wire      [7:0] n14906;
wire            n14907;
wire            n14908;
wire            n14909;
wire            n1491;
wire            n14910;
wire            n14911;
wire      [7:0] n14912;
wire            n14913;
wire            n14914;
wire            n14915;
wire            n14916;
wire            n14917;
wire      [7:0] n14918;
wire            n14919;
wire            n1492;
wire            n14920;
wire            n14921;
wire            n14922;
wire            n14923;
wire      [7:0] n14924;
wire            n14925;
wire            n14926;
wire            n14927;
wire            n14928;
wire            n14929;
wire            n1493;
wire      [7:0] n14930;
wire            n14931;
wire            n14932;
wire            n14933;
wire            n14934;
wire            n14935;
wire      [7:0] n14936;
wire            n14937;
wire            n14938;
wire            n14939;
wire            n1494;
wire            n14940;
wire            n14941;
wire      [7:0] n14942;
wire            n14943;
wire            n14944;
wire            n14945;
wire            n14946;
wire            n14947;
wire      [7:0] n14948;
wire            n14949;
wire            n1495;
wire            n14950;
wire            n14951;
wire            n14952;
wire            n14953;
wire      [7:0] n14954;
wire            n14955;
wire            n14956;
wire            n14957;
wire            n14958;
wire            n14959;
wire            n1496;
wire      [7:0] n14960;
wire            n14961;
wire            n14962;
wire            n14963;
wire            n14964;
wire            n14965;
wire      [7:0] n14966;
wire            n14967;
wire            n14968;
wire            n14969;
wire            n1497;
wire            n14970;
wire            n14971;
wire      [7:0] n14972;
wire            n14973;
wire            n14974;
wire            n14975;
wire            n14976;
wire            n14977;
wire      [7:0] n14978;
wire            n14979;
wire            n1498;
wire            n14980;
wire            n14981;
wire            n14982;
wire            n14983;
wire      [7:0] n14984;
wire            n14985;
wire            n14986;
wire            n14987;
wire            n14988;
wire            n14989;
wire            n1499;
wire      [7:0] n14990;
wire            n14991;
wire            n14992;
wire            n14993;
wire            n14994;
wire            n14995;
wire      [7:0] n14996;
wire            n14997;
wire            n14998;
wire            n14999;
wire            n15;
wire            n150;
wire            n1500;
wire            n15000;
wire            n15001;
wire      [7:0] n15002;
wire            n15003;
wire            n15004;
wire            n15005;
wire            n15006;
wire            n15007;
wire      [7:0] n15008;
wire            n15009;
wire            n1501;
wire            n15010;
wire            n15011;
wire            n15012;
wire            n15013;
wire      [7:0] n15014;
wire            n15015;
wire            n15016;
wire            n15017;
wire            n15018;
wire            n15019;
wire            n1502;
wire      [7:0] n15020;
wire            n15021;
wire            n15022;
wire            n15023;
wire            n15024;
wire            n15025;
wire      [7:0] n15026;
wire            n15027;
wire            n15028;
wire            n15029;
wire            n1503;
wire            n15030;
wire            n15031;
wire      [7:0] n15032;
wire            n15033;
wire            n15034;
wire            n15035;
wire            n15036;
wire            n15037;
wire      [7:0] n15038;
wire            n15039;
wire            n1504;
wire            n15040;
wire            n15041;
wire            n15042;
wire            n15043;
wire      [7:0] n15044;
wire            n15045;
wire            n15046;
wire            n15047;
wire            n15048;
wire            n15049;
wire            n1505;
wire      [7:0] n15050;
wire            n15051;
wire            n15052;
wire            n15053;
wire            n15054;
wire            n15055;
wire      [7:0] n15056;
wire            n15057;
wire            n15058;
wire            n15059;
wire            n1506;
wire            n15060;
wire            n15061;
wire      [7:0] n15062;
wire            n15063;
wire            n15064;
wire            n15065;
wire            n15066;
wire            n15067;
wire      [7:0] n15068;
wire            n15069;
wire            n1507;
wire            n15070;
wire            n15071;
wire            n15072;
wire            n15073;
wire      [7:0] n15074;
wire            n15075;
wire            n15076;
wire            n15077;
wire            n15078;
wire            n15079;
wire            n1508;
wire      [7:0] n15080;
wire            n15081;
wire            n15082;
wire            n15083;
wire            n15084;
wire            n15085;
wire      [7:0] n15086;
wire            n15087;
wire            n15088;
wire            n15089;
wire            n1509;
wire            n15090;
wire            n15091;
wire      [7:0] n15092;
wire            n15093;
wire            n15094;
wire            n15095;
wire            n15096;
wire            n15097;
wire      [7:0] n15098;
wire            n15099;
wire            n1510;
wire            n15100;
wire            n15101;
wire            n15102;
wire            n15103;
wire      [7:0] n15104;
wire            n15105;
wire            n15106;
wire            n15107;
wire            n15108;
wire            n15109;
wire            n1511;
wire      [7:0] n15110;
wire            n15111;
wire            n15112;
wire            n15113;
wire            n15114;
wire            n15115;
wire      [7:0] n15116;
wire            n15117;
wire            n15118;
wire            n15119;
wire            n1512;
wire            n15120;
wire            n15121;
wire      [7:0] n15122;
wire            n15123;
wire            n15124;
wire            n15125;
wire            n15126;
wire            n15127;
wire      [7:0] n15128;
wire            n15129;
wire            n1513;
wire            n15130;
wire            n15131;
wire            n15132;
wire            n15133;
wire      [7:0] n15134;
wire            n15135;
wire            n15136;
wire            n15137;
wire            n15138;
wire            n15139;
wire            n1514;
wire      [7:0] n15140;
wire            n15141;
wire            n15142;
wire            n15143;
wire            n15144;
wire            n15145;
wire      [7:0] n15146;
wire            n15147;
wire            n15148;
wire            n15149;
wire            n1515;
wire            n15150;
wire            n15151;
wire      [7:0] n15152;
wire            n15153;
wire            n15154;
wire            n15155;
wire            n15156;
wire            n15157;
wire      [7:0] n15158;
wire            n15159;
wire            n1516;
wire            n15160;
wire            n15161;
wire            n15162;
wire            n15163;
wire      [7:0] n15164;
wire            n15165;
wire            n15166;
wire            n15167;
wire            n15168;
wire            n15169;
wire            n1517;
wire      [7:0] n15170;
wire            n15171;
wire            n15172;
wire            n15173;
wire            n15174;
wire            n15175;
wire      [7:0] n15176;
wire            n15177;
wire            n15178;
wire            n15179;
wire            n1518;
wire            n15180;
wire            n15181;
wire      [7:0] n15182;
wire            n15183;
wire            n15184;
wire            n15185;
wire            n15186;
wire            n15187;
wire      [7:0] n15188;
wire            n15189;
wire            n1519;
wire            n15190;
wire            n15191;
wire            n15192;
wire            n15193;
wire      [7:0] n15194;
wire            n15195;
wire            n15196;
wire            n15197;
wire            n15198;
wire            n15199;
wire            n152;
wire            n1520;
wire      [7:0] n15200;
wire            n15201;
wire            n15202;
wire            n15203;
wire            n15204;
wire            n15205;
wire      [7:0] n15206;
wire            n15207;
wire            n15208;
wire            n15209;
wire            n1521;
wire            n15210;
wire            n15211;
wire      [7:0] n15212;
wire            n15213;
wire            n15214;
wire            n15215;
wire            n15216;
wire            n15217;
wire      [7:0] n15218;
wire            n15219;
wire            n1522;
wire            n15220;
wire            n15221;
wire            n15222;
wire            n15223;
wire      [7:0] n15224;
wire            n15225;
wire            n15226;
wire            n15227;
wire            n15228;
wire            n15229;
wire            n1523;
wire      [7:0] n15230;
wire            n15231;
wire            n15232;
wire            n15233;
wire            n15234;
wire            n15235;
wire      [7:0] n15236;
wire            n15237;
wire            n15238;
wire            n15239;
wire            n1524;
wire            n15240;
wire            n15241;
wire      [7:0] n15242;
wire            n15243;
wire            n15244;
wire            n15245;
wire            n15246;
wire            n15247;
wire      [7:0] n15248;
wire            n15249;
wire            n1525;
wire            n15250;
wire            n15251;
wire            n15252;
wire            n15253;
wire      [7:0] n15254;
wire            n15255;
wire            n15256;
wire            n15257;
wire            n15258;
wire            n15259;
wire            n1526;
wire      [7:0] n15260;
wire            n15261;
wire            n15262;
wire            n15263;
wire            n15264;
wire            n15265;
wire      [7:0] n15266;
wire            n15267;
wire            n15268;
wire            n15269;
wire            n1527;
wire            n15270;
wire            n15271;
wire      [7:0] n15272;
wire            n15273;
wire            n15274;
wire            n15275;
wire            n15276;
wire            n15277;
wire      [7:0] n15278;
wire            n15279;
wire            n1528;
wire            n15280;
wire            n15281;
wire            n15282;
wire            n15283;
wire      [7:0] n15284;
wire            n15285;
wire            n15286;
wire            n15287;
wire            n15288;
wire            n15289;
wire            n1529;
wire      [7:0] n15290;
wire            n15291;
wire            n15292;
wire            n15293;
wire            n15294;
wire            n15295;
wire      [7:0] n15296;
wire            n15297;
wire            n15298;
wire            n15299;
wire            n1530;
wire            n15300;
wire            n15301;
wire      [7:0] n15302;
wire            n15303;
wire            n15304;
wire            n15305;
wire            n15306;
wire            n15307;
wire      [7:0] n15308;
wire            n15309;
wire            n1531;
wire            n15310;
wire            n15311;
wire            n15312;
wire            n15313;
wire      [7:0] n15314;
wire            n15315;
wire            n15316;
wire            n15317;
wire            n15318;
wire            n15319;
wire            n1532;
wire      [7:0] n15320;
wire            n15321;
wire            n15322;
wire            n15323;
wire            n15324;
wire            n15325;
wire      [7:0] n15326;
wire            n15327;
wire            n15328;
wire            n15329;
wire            n1533;
wire            n15330;
wire            n15331;
wire      [7:0] n15332;
wire            n15333;
wire            n15334;
wire            n15335;
wire            n15336;
wire            n15337;
wire      [7:0] n15338;
wire            n15339;
wire            n1534;
wire            n15340;
wire            n15341;
wire            n15342;
wire            n15343;
wire      [7:0] n15344;
wire            n15345;
wire            n15346;
wire            n15347;
wire            n15348;
wire            n15349;
wire            n1535;
wire      [7:0] n15350;
wire            n15351;
wire            n15352;
wire            n15353;
wire            n15354;
wire            n15355;
wire      [7:0] n15356;
wire            n15357;
wire            n15358;
wire            n15359;
wire            n1536;
wire            n15360;
wire            n15361;
wire      [7:0] n15362;
wire            n15363;
wire            n15364;
wire            n15365;
wire            n15366;
wire            n15367;
wire      [7:0] n15368;
wire            n15369;
wire            n1537;
wire            n15370;
wire            n15371;
wire            n15372;
wire            n15373;
wire      [7:0] n15374;
wire            n15375;
wire            n15376;
wire            n15377;
wire            n15378;
wire            n15379;
wire            n1538;
wire      [7:0] n15380;
wire            n15381;
wire            n15382;
wire            n15383;
wire            n15384;
wire            n15385;
wire      [7:0] n15386;
wire            n15387;
wire            n15388;
wire            n15389;
wire            n1539;
wire            n15390;
wire            n15391;
wire      [7:0] n15392;
wire            n15393;
wire            n15394;
wire            n15395;
wire            n15396;
wire            n15397;
wire      [7:0] n15398;
wire            n15399;
wire            n154;
wire            n1540;
wire            n15400;
wire            n15401;
wire            n15402;
wire            n15403;
wire      [7:0] n15404;
wire            n15405;
wire            n15406;
wire            n15407;
wire            n15408;
wire            n15409;
wire            n1541;
wire      [7:0] n15410;
wire            n15411;
wire            n15412;
wire            n15413;
wire            n15414;
wire            n15415;
wire      [7:0] n15416;
wire            n15417;
wire            n15418;
wire            n15419;
wire            n1542;
wire            n15420;
wire            n15421;
wire      [7:0] n15422;
wire            n15423;
wire            n15424;
wire            n15425;
wire            n15426;
wire            n15427;
wire      [7:0] n15428;
wire            n15429;
wire            n1543;
wire            n15430;
wire            n15431;
wire            n15432;
wire            n15433;
wire      [7:0] n15434;
wire            n15435;
wire            n15436;
wire            n15437;
wire            n15438;
wire            n15439;
wire            n1544;
wire      [7:0] n15440;
wire            n15441;
wire            n15442;
wire            n15443;
wire            n15444;
wire            n15445;
wire      [7:0] n15446;
wire            n15447;
wire            n15448;
wire            n15449;
wire            n1545;
wire            n15450;
wire            n15451;
wire      [7:0] n15452;
wire            n15453;
wire            n15454;
wire            n15455;
wire            n15456;
wire            n15457;
wire      [7:0] n15458;
wire            n15459;
wire            n1546;
wire            n15460;
wire            n15461;
wire            n15462;
wire            n15463;
wire      [7:0] n15464;
wire            n15465;
wire            n15466;
wire            n15467;
wire            n15468;
wire            n15469;
wire            n1547;
wire      [7:0] n15470;
wire            n15471;
wire            n15472;
wire            n15473;
wire            n15474;
wire            n15475;
wire      [7:0] n15476;
wire            n15477;
wire            n15478;
wire            n15479;
wire            n1548;
wire            n15480;
wire            n15481;
wire      [7:0] n15482;
wire            n15483;
wire            n15484;
wire            n15485;
wire            n15486;
wire            n15487;
wire      [7:0] n15488;
wire            n15489;
wire            n1549;
wire            n15490;
wire            n15491;
wire            n15492;
wire            n15493;
wire      [7:0] n15494;
wire            n15495;
wire            n15496;
wire            n15497;
wire            n15498;
wire            n15499;
wire            n1550;
wire      [7:0] n15500;
wire            n15501;
wire            n15502;
wire            n15503;
wire            n15504;
wire            n15505;
wire      [7:0] n15506;
wire            n15507;
wire            n15508;
wire            n15509;
wire            n1551;
wire            n15510;
wire            n15511;
wire      [7:0] n15512;
wire            n15513;
wire            n15514;
wire            n15515;
wire            n15516;
wire            n15517;
wire      [7:0] n15518;
wire            n15519;
wire            n1552;
wire            n15520;
wire            n15521;
wire            n15522;
wire            n15523;
wire      [7:0] n15524;
wire            n15525;
wire            n15526;
wire            n15527;
wire            n15528;
wire            n15529;
wire            n1553;
wire      [7:0] n15530;
wire            n15531;
wire            n15532;
wire            n15533;
wire            n15534;
wire            n15535;
wire      [7:0] n15536;
wire            n15537;
wire            n15538;
wire            n15539;
wire            n1554;
wire            n15540;
wire            n15541;
wire      [7:0] n15542;
wire            n15543;
wire            n15544;
wire            n15545;
wire            n15546;
wire            n15547;
wire      [7:0] n15548;
wire            n15549;
wire            n1555;
wire            n15550;
wire            n15551;
wire            n15552;
wire            n15553;
wire      [7:0] n15554;
wire            n15555;
wire            n15556;
wire            n15557;
wire            n15558;
wire            n15559;
wire            n1556;
wire      [7:0] n15560;
wire            n15561;
wire            n15562;
wire            n15563;
wire            n15564;
wire            n15565;
wire      [7:0] n15566;
wire            n15567;
wire            n15568;
wire            n15569;
wire            n1557;
wire            n15570;
wire            n15571;
wire      [7:0] n15572;
wire            n15573;
wire            n15574;
wire            n15575;
wire            n15576;
wire            n15577;
wire      [7:0] n15578;
wire            n15579;
wire            n1558;
wire            n15580;
wire            n15581;
wire            n15582;
wire            n15583;
wire      [7:0] n15584;
wire            n15585;
wire            n15586;
wire            n15587;
wire            n15588;
wire            n15589;
wire            n1559;
wire      [7:0] n15590;
wire            n15591;
wire            n15592;
wire            n15593;
wire            n15594;
wire            n15595;
wire      [7:0] n15596;
wire            n15597;
wire            n15598;
wire            n15599;
wire            n156;
wire            n1560;
wire            n15600;
wire            n15601;
wire      [7:0] n15602;
wire            n15603;
wire            n15604;
wire            n15605;
wire            n15606;
wire            n15607;
wire      [7:0] n15608;
wire            n15609;
wire            n1561;
wire            n15610;
wire            n15611;
wire            n15612;
wire            n15613;
wire      [7:0] n15614;
wire            n15615;
wire            n15616;
wire            n15617;
wire            n15618;
wire            n15619;
wire            n1562;
wire      [7:0] n15620;
wire            n15621;
wire            n15622;
wire            n15623;
wire            n15624;
wire            n15625;
wire      [7:0] n15626;
wire            n15627;
wire            n15628;
wire            n15629;
wire            n1563;
wire            n15630;
wire            n15631;
wire      [7:0] n15632;
wire            n15633;
wire            n15634;
wire            n15635;
wire            n15636;
wire            n15637;
wire      [7:0] n15638;
wire            n15639;
wire            n1564;
wire            n15640;
wire            n15641;
wire            n15642;
wire            n15643;
wire      [7:0] n15644;
wire            n15645;
wire            n15646;
wire            n15647;
wire            n15648;
wire            n15649;
wire            n1565;
wire      [7:0] n15650;
wire            n15651;
wire            n15652;
wire            n15653;
wire            n15654;
wire            n15655;
wire      [7:0] n15656;
wire            n15657;
wire            n15658;
wire            n15659;
wire            n1566;
wire            n15660;
wire            n15661;
wire      [7:0] n15662;
wire            n15663;
wire            n15664;
wire            n15665;
wire            n15666;
wire            n15667;
wire      [7:0] n15668;
wire            n15669;
wire            n1567;
wire            n15670;
wire            n15671;
wire            n15672;
wire            n15673;
wire      [7:0] n15674;
wire            n15675;
wire            n15676;
wire            n15677;
wire            n15678;
wire            n15679;
wire            n1568;
wire      [7:0] n15680;
wire            n15681;
wire            n15682;
wire            n15683;
wire            n15684;
wire            n15685;
wire      [7:0] n15686;
wire            n15687;
wire            n15688;
wire            n15689;
wire            n1569;
wire            n15690;
wire            n15691;
wire      [7:0] n15692;
wire            n15693;
wire            n15694;
wire            n15695;
wire            n15696;
wire            n15697;
wire      [7:0] n15698;
wire            n15699;
wire            n1570;
wire            n15700;
wire            n15701;
wire            n15702;
wire            n15703;
wire      [7:0] n15704;
wire            n15705;
wire            n15706;
wire            n15707;
wire            n15708;
wire            n15709;
wire            n1571;
wire      [7:0] n15710;
wire            n15711;
wire            n15712;
wire            n15713;
wire            n15714;
wire            n15715;
wire      [7:0] n15716;
wire            n15717;
wire            n15718;
wire            n15719;
wire            n1572;
wire            n15720;
wire            n15721;
wire      [7:0] n15722;
wire            n15723;
wire            n15724;
wire            n15725;
wire            n15726;
wire            n15727;
wire      [7:0] n15728;
wire            n15729;
wire            n1573;
wire            n15730;
wire            n15731;
wire            n15732;
wire            n15733;
wire      [7:0] n15734;
wire            n15735;
wire            n15736;
wire            n15737;
wire            n15738;
wire            n15739;
wire            n1574;
wire      [7:0] n15740;
wire            n15741;
wire            n15742;
wire            n15743;
wire            n15744;
wire            n15745;
wire      [7:0] n15746;
wire            n15747;
wire            n15748;
wire            n15749;
wire            n1575;
wire            n15750;
wire            n15751;
wire      [7:0] n15752;
wire            n15753;
wire            n15754;
wire            n15755;
wire            n15756;
wire            n15757;
wire      [7:0] n15758;
wire            n15759;
wire            n1576;
wire            n15760;
wire            n15761;
wire            n15762;
wire            n15763;
wire      [7:0] n15764;
wire            n15765;
wire            n15766;
wire            n15767;
wire            n15768;
wire            n15769;
wire            n1577;
wire      [7:0] n15770;
wire            n15771;
wire            n15772;
wire            n15773;
wire            n15774;
wire            n15775;
wire      [7:0] n15776;
wire            n15777;
wire            n15778;
wire            n15779;
wire            n1578;
wire            n15780;
wire            n15781;
wire      [7:0] n15782;
wire            n15783;
wire            n15784;
wire            n15785;
wire            n15786;
wire            n15787;
wire      [7:0] n15788;
wire            n15789;
wire            n1579;
wire            n15790;
wire            n15791;
wire            n15792;
wire            n15793;
wire      [7:0] n15794;
wire            n15795;
wire            n15796;
wire            n15797;
wire            n15798;
wire            n15799;
wire            n158;
wire            n1580;
wire      [7:0] n15800;
wire            n15801;
wire            n15802;
wire            n15803;
wire            n15804;
wire            n15805;
wire      [7:0] n15806;
wire            n15807;
wire            n15808;
wire            n15809;
wire            n1581;
wire            n15810;
wire            n15811;
wire      [7:0] n15812;
wire            n15813;
wire            n15814;
wire            n15815;
wire            n15816;
wire            n15817;
wire      [7:0] n15818;
wire            n15819;
wire            n1582;
wire            n15820;
wire            n15821;
wire            n15822;
wire            n15823;
wire      [7:0] n15824;
wire            n15825;
wire            n15826;
wire            n15827;
wire            n15828;
wire            n15829;
wire            n1583;
wire      [7:0] n15830;
wire            n15831;
wire            n15832;
wire            n15833;
wire            n15834;
wire            n15835;
wire      [7:0] n15836;
wire            n15837;
wire            n15838;
wire            n15839;
wire            n1584;
wire            n15840;
wire            n15841;
wire      [7:0] n15842;
wire            n15843;
wire            n15844;
wire            n15845;
wire            n15846;
wire            n15847;
wire      [7:0] n15848;
wire            n15849;
wire            n1585;
wire            n15850;
wire            n15851;
wire            n15852;
wire            n15853;
wire      [7:0] n15854;
wire            n15855;
wire            n15856;
wire            n15857;
wire            n15858;
wire            n15859;
wire            n1586;
wire      [7:0] n15860;
wire            n15861;
wire            n15862;
wire            n15863;
wire            n15864;
wire            n15865;
wire      [7:0] n15866;
wire            n15867;
wire            n15868;
wire            n15869;
wire            n1587;
wire            n15870;
wire            n15871;
wire      [7:0] n15872;
wire            n15873;
wire            n15874;
wire            n15875;
wire            n15876;
wire            n15877;
wire      [7:0] n15878;
wire            n15879;
wire            n1588;
wire            n15880;
wire            n15881;
wire            n15882;
wire            n15883;
wire      [7:0] n15884;
wire            n15885;
wire            n15886;
wire            n15887;
wire            n15888;
wire            n15889;
wire            n1589;
wire      [7:0] n15890;
wire            n15891;
wire            n15892;
wire            n15893;
wire            n15894;
wire            n15895;
wire      [7:0] n15896;
wire            n15897;
wire            n15898;
wire            n15899;
wire            n1590;
wire            n15900;
wire            n15901;
wire      [7:0] n15902;
wire            n15903;
wire            n15904;
wire            n15905;
wire            n15906;
wire            n15907;
wire      [7:0] n15908;
wire            n15909;
wire            n1591;
wire            n15910;
wire            n15911;
wire            n15912;
wire            n15913;
wire      [7:0] n15914;
wire            n15915;
wire            n15916;
wire            n15917;
wire            n15918;
wire            n15919;
wire            n1592;
wire      [7:0] n15920;
wire            n15921;
wire            n15922;
wire            n15923;
wire            n15924;
wire            n15925;
wire      [7:0] n15926;
wire            n15927;
wire            n15928;
wire            n15929;
wire            n1593;
wire            n15930;
wire            n15931;
wire      [7:0] n15932;
wire            n15933;
wire            n15934;
wire            n15935;
wire            n15936;
wire            n15937;
wire      [7:0] n15938;
wire            n15939;
wire            n1594;
wire            n15940;
wire            n15941;
wire            n15942;
wire            n15943;
wire      [7:0] n15944;
wire            n15945;
wire            n15946;
wire            n15947;
wire            n15948;
wire            n15949;
wire            n1595;
wire      [7:0] n15950;
wire            n15951;
wire            n15952;
wire            n15953;
wire            n15954;
wire            n15955;
wire      [7:0] n15956;
wire            n15957;
wire            n15958;
wire            n15959;
wire            n1596;
wire            n15960;
wire            n15961;
wire      [7:0] n15962;
wire            n15963;
wire            n15964;
wire            n15965;
wire            n15966;
wire            n15967;
wire      [7:0] n15968;
wire            n15969;
wire            n1597;
wire            n15970;
wire            n15971;
wire            n15972;
wire            n15973;
wire      [7:0] n15974;
wire            n15975;
wire            n15976;
wire            n15977;
wire            n15978;
wire            n15979;
wire            n1598;
wire      [7:0] n15980;
wire            n15981;
wire            n15982;
wire            n15983;
wire            n15984;
wire            n15985;
wire      [7:0] n15986;
wire            n15987;
wire            n15988;
wire            n15989;
wire            n1599;
wire            n15990;
wire            n15991;
wire      [7:0] n15992;
wire            n15993;
wire            n15994;
wire            n15995;
wire            n15996;
wire            n15997;
wire      [7:0] n15998;
wire            n15999;
wire            n160;
wire            n1600;
wire            n16000;
wire            n16001;
wire            n16002;
wire            n16003;
wire      [7:0] n16004;
wire            n16005;
wire            n16006;
wire            n16007;
wire            n16008;
wire            n16009;
wire            n1601;
wire      [7:0] n16010;
wire            n16011;
wire            n16012;
wire            n16013;
wire            n16014;
wire            n16015;
wire      [7:0] n16016;
wire            n16017;
wire            n16018;
wire            n16019;
wire            n1602;
wire            n16020;
wire            n16021;
wire      [7:0] n16022;
wire            n16023;
wire            n16024;
wire            n16025;
wire            n16026;
wire            n16027;
wire      [7:0] n16028;
wire            n16029;
wire            n1603;
wire            n16030;
wire            n16031;
wire            n16032;
wire            n16033;
wire      [7:0] n16034;
wire            n16035;
wire            n16036;
wire            n16037;
wire            n16038;
wire            n16039;
wire            n1604;
wire      [7:0] n16040;
wire            n16041;
wire            n16042;
wire            n16043;
wire            n16044;
wire            n16045;
wire      [7:0] n16046;
wire            n16047;
wire            n16048;
wire            n16049;
wire            n1605;
wire            n16050;
wire            n16051;
wire      [7:0] n16052;
wire            n16053;
wire            n16054;
wire            n16055;
wire            n16056;
wire            n16057;
wire      [7:0] n16058;
wire            n16059;
wire            n1606;
wire            n16060;
wire            n16061;
wire            n16062;
wire            n16063;
wire      [7:0] n16064;
wire            n16065;
wire            n16066;
wire            n16067;
wire            n16068;
wire            n16069;
wire            n1607;
wire      [7:0] n16070;
wire            n16071;
wire            n16072;
wire            n16073;
wire            n16074;
wire            n16075;
wire      [7:0] n16076;
wire            n16077;
wire            n16078;
wire            n16079;
wire            n1608;
wire            n16080;
wire            n16081;
wire      [7:0] n16082;
wire            n16083;
wire            n16084;
wire            n16085;
wire            n16086;
wire            n16087;
wire      [7:0] n16088;
wire            n16089;
wire            n1609;
wire            n16090;
wire            n16091;
wire            n16092;
wire            n16093;
wire      [7:0] n16094;
wire            n16095;
wire            n16096;
wire            n16097;
wire            n16098;
wire            n16099;
wire      [7:0] n1610;
wire      [7:0] n16100;
wire            n16101;
wire            n16102;
wire            n16103;
wire            n16104;
wire            n16105;
wire      [7:0] n16106;
wire            n16107;
wire            n16108;
wire            n16109;
wire      [7:0] n1611;
wire            n16110;
wire            n16111;
wire      [7:0] n16112;
wire            n16113;
wire            n16114;
wire            n16115;
wire            n16116;
wire            n16117;
wire      [7:0] n16118;
wire            n16119;
wire      [7:0] n1612;
wire            n16120;
wire            n16121;
wire            n16122;
wire            n16123;
wire      [7:0] n16124;
wire            n16125;
wire            n16126;
wire            n16127;
wire            n16128;
wire            n16129;
wire      [7:0] n1613;
wire      [7:0] n16130;
wire            n16131;
wire            n16132;
wire            n16133;
wire            n16134;
wire            n16135;
wire      [7:0] n16136;
wire            n16137;
wire            n16138;
wire            n16139;
wire      [7:0] n1614;
wire            n16140;
wire            n16141;
wire      [7:0] n16142;
wire            n16143;
wire            n16144;
wire            n16145;
wire            n16146;
wire            n16147;
wire      [7:0] n16148;
wire            n16149;
wire      [7:0] n1615;
wire            n16150;
wire            n16151;
wire            n16152;
wire            n16153;
wire      [7:0] n16154;
wire            n16155;
wire            n16156;
wire            n16157;
wire            n16158;
wire            n16159;
wire      [7:0] n1616;
wire      [7:0] n16160;
wire            n16161;
wire            n16162;
wire            n16163;
wire            n16164;
wire            n16165;
wire      [7:0] n16166;
wire            n16167;
wire            n16168;
wire            n16169;
wire      [7:0] n1617;
wire            n16170;
wire            n16171;
wire      [7:0] n16172;
wire            n16173;
wire            n16174;
wire            n16175;
wire            n16176;
wire            n16177;
wire      [7:0] n16178;
wire            n16179;
wire      [7:0] n1618;
wire            n16180;
wire            n16181;
wire            n16182;
wire            n16183;
wire      [7:0] n16184;
wire            n16185;
wire            n16186;
wire            n16187;
wire            n16188;
wire            n16189;
wire      [7:0] n1619;
wire      [7:0] n16190;
wire            n16191;
wire            n16192;
wire            n16193;
wire            n16194;
wire            n16195;
wire      [7:0] n16196;
wire            n16197;
wire            n16198;
wire            n16199;
wire            n162;
wire      [7:0] n1620;
wire            n16200;
wire            n16201;
wire      [7:0] n16202;
wire            n16203;
wire            n16204;
wire            n16205;
wire            n16206;
wire            n16207;
wire      [7:0] n16208;
wire            n16209;
wire      [7:0] n1621;
wire            n16210;
wire            n16211;
wire            n16212;
wire            n16213;
wire      [7:0] n16214;
wire            n16215;
wire            n16216;
wire            n16217;
wire            n16218;
wire            n16219;
wire      [7:0] n1622;
wire      [7:0] n16220;
wire            n16221;
wire            n16222;
wire            n16223;
wire            n16224;
wire            n16225;
wire      [7:0] n16226;
wire            n16227;
wire            n16228;
wire            n16229;
wire      [7:0] n1623;
wire            n16230;
wire            n16231;
wire      [7:0] n16232;
wire            n16233;
wire            n16234;
wire            n16235;
wire            n16236;
wire            n16237;
wire      [7:0] n16238;
wire            n16239;
wire      [7:0] n1624;
wire            n16240;
wire            n16241;
wire            n16242;
wire            n16243;
wire      [7:0] n16244;
wire            n16245;
wire            n16246;
wire            n16247;
wire            n16248;
wire            n16249;
wire      [7:0] n1625;
wire      [7:0] n16250;
wire            n16251;
wire            n16252;
wire            n16253;
wire            n16254;
wire            n16255;
wire      [7:0] n16256;
wire            n16257;
wire            n16258;
wire            n16259;
wire      [7:0] n1626;
wire            n16260;
wire            n16261;
wire      [7:0] n16262;
wire            n16263;
wire            n16264;
wire            n16265;
wire            n16266;
wire            n16267;
wire      [7:0] n16268;
wire            n16269;
wire      [7:0] n1627;
wire            n16270;
wire            n16271;
wire            n16272;
wire            n16273;
wire      [7:0] n16274;
wire            n16275;
wire            n16276;
wire            n16277;
wire            n16278;
wire            n16279;
wire      [7:0] n1628;
wire      [7:0] n16280;
wire            n16281;
wire            n16282;
wire            n16283;
wire            n16284;
wire            n16285;
wire      [7:0] n16286;
wire            n16287;
wire            n16288;
wire            n16289;
wire      [7:0] n1629;
wire            n16290;
wire            n16291;
wire      [7:0] n16292;
wire            n16293;
wire            n16294;
wire            n16295;
wire            n16296;
wire            n16297;
wire      [7:0] n16298;
wire            n16299;
wire      [7:0] n1630;
wire            n16300;
wire            n16301;
wire            n16302;
wire            n16303;
wire      [7:0] n16304;
wire            n16305;
wire            n16306;
wire            n16307;
wire            n16308;
wire            n16309;
wire      [7:0] n1631;
wire      [7:0] n16310;
wire            n16311;
wire            n16312;
wire            n16313;
wire            n16314;
wire            n16315;
wire      [7:0] n16316;
wire            n16317;
wire            n16318;
wire            n16319;
wire      [7:0] n1632;
wire            n16320;
wire            n16321;
wire      [7:0] n16322;
wire            n16323;
wire            n16324;
wire            n16325;
wire            n16326;
wire            n16327;
wire      [7:0] n16328;
wire            n16329;
wire      [7:0] n1633;
wire            n16330;
wire            n16331;
wire            n16332;
wire            n16333;
wire      [7:0] n16334;
wire            n16335;
wire            n16336;
wire            n16337;
wire            n16338;
wire            n16339;
wire      [7:0] n1634;
wire      [7:0] n16340;
wire            n16341;
wire            n16342;
wire            n16343;
wire            n16344;
wire            n16345;
wire      [7:0] n16346;
wire            n16347;
wire            n16348;
wire            n16349;
wire      [7:0] n1635;
wire            n16350;
wire            n16351;
wire      [7:0] n16352;
wire            n16353;
wire            n16354;
wire            n16355;
wire            n16356;
wire            n16357;
wire      [7:0] n16358;
wire            n16359;
wire      [7:0] n1636;
wire            n16360;
wire            n16361;
wire            n16362;
wire            n16363;
wire      [7:0] n16364;
wire            n16365;
wire            n16366;
wire            n16367;
wire            n16368;
wire            n16369;
wire      [7:0] n1637;
wire      [7:0] n16370;
wire            n16371;
wire            n16372;
wire            n16373;
wire            n16374;
wire            n16375;
wire      [7:0] n16376;
wire            n16377;
wire            n16378;
wire            n16379;
wire      [7:0] n1638;
wire            n16380;
wire            n16381;
wire      [7:0] n16382;
wire            n16383;
wire            n16384;
wire            n16385;
wire            n16386;
wire            n16387;
wire      [7:0] n16388;
wire            n16389;
wire      [7:0] n1639;
wire            n16390;
wire            n16391;
wire            n16392;
wire            n16393;
wire      [7:0] n16394;
wire            n16395;
wire            n16396;
wire            n16397;
wire            n16398;
wire            n16399;
wire            n164;
wire      [7:0] n1640;
wire      [7:0] n16400;
wire            n16401;
wire            n16402;
wire            n16403;
wire            n16404;
wire            n16405;
wire      [7:0] n16406;
wire            n16407;
wire            n16408;
wire            n16409;
wire      [7:0] n1641;
wire            n16410;
wire            n16411;
wire      [7:0] n16412;
wire            n16413;
wire            n16414;
wire            n16415;
wire            n16416;
wire            n16417;
wire      [7:0] n16418;
wire            n16419;
wire      [7:0] n1642;
wire            n16420;
wire            n16421;
wire            n16422;
wire            n16423;
wire      [7:0] n16424;
wire            n16425;
wire            n16426;
wire            n16427;
wire            n16428;
wire            n16429;
wire      [7:0] n1643;
wire      [7:0] n16430;
wire            n16431;
wire            n16432;
wire            n16433;
wire            n16434;
wire            n16435;
wire      [7:0] n16436;
wire            n16437;
wire            n16438;
wire            n16439;
wire      [7:0] n1644;
wire            n16440;
wire            n16441;
wire      [7:0] n16442;
wire            n16443;
wire            n16444;
wire            n16445;
wire            n16446;
wire            n16447;
wire      [7:0] n16448;
wire            n16449;
wire      [7:0] n1645;
wire            n16450;
wire            n16451;
wire            n16452;
wire            n16453;
wire      [7:0] n16454;
wire            n16455;
wire            n16456;
wire            n16457;
wire            n16458;
wire            n16459;
wire      [7:0] n1646;
wire      [7:0] n16460;
wire            n16461;
wire            n16462;
wire            n16463;
wire            n16464;
wire            n16465;
wire      [7:0] n16466;
wire            n16467;
wire            n16468;
wire            n16469;
wire      [7:0] n1647;
wire            n16470;
wire            n16471;
wire      [7:0] n16472;
wire            n16473;
wire            n16474;
wire            n16475;
wire            n16476;
wire            n16477;
wire      [7:0] n16478;
wire            n16479;
wire      [7:0] n1648;
wire            n16480;
wire            n16481;
wire            n16482;
wire            n16483;
wire      [7:0] n16484;
wire            n16485;
wire            n16486;
wire            n16487;
wire            n16488;
wire            n16489;
wire      [7:0] n1649;
wire      [7:0] n16490;
wire            n16491;
wire            n16492;
wire            n16493;
wire            n16494;
wire            n16495;
wire      [7:0] n16496;
wire            n16497;
wire            n16498;
wire            n16499;
wire      [7:0] n1650;
wire            n16500;
wire            n16501;
wire      [7:0] n16502;
wire            n16503;
wire            n16504;
wire            n16505;
wire            n16506;
wire            n16507;
wire      [7:0] n16508;
wire            n16509;
wire      [7:0] n1651;
wire            n16510;
wire            n16511;
wire            n16512;
wire            n16513;
wire      [7:0] n16514;
wire            n16515;
wire            n16516;
wire            n16517;
wire            n16518;
wire            n16519;
wire      [7:0] n1652;
wire      [7:0] n16520;
wire            n16521;
wire            n16522;
wire            n16523;
wire            n16524;
wire            n16525;
wire      [7:0] n16526;
wire            n16527;
wire            n16528;
wire            n16529;
wire      [7:0] n1653;
wire            n16530;
wire            n16531;
wire      [7:0] n16532;
wire            n16533;
wire            n16534;
wire            n16535;
wire            n16536;
wire            n16537;
wire      [7:0] n16538;
wire            n16539;
wire      [7:0] n1654;
wire            n16540;
wire            n16541;
wire            n16542;
wire            n16543;
wire      [7:0] n16544;
wire            n16545;
wire            n16546;
wire            n16547;
wire            n16548;
wire            n16549;
wire      [7:0] n1655;
wire      [7:0] n16550;
wire            n16551;
wire            n16552;
wire            n16553;
wire            n16554;
wire            n16555;
wire      [7:0] n16556;
wire            n16557;
wire            n16558;
wire            n16559;
wire      [7:0] n1656;
wire            n16560;
wire            n16561;
wire      [7:0] n16562;
wire            n16563;
wire            n16564;
wire            n16565;
wire            n16566;
wire            n16567;
wire      [7:0] n16568;
wire            n16569;
wire      [7:0] n1657;
wire            n16570;
wire            n16571;
wire            n16572;
wire            n16573;
wire      [7:0] n16574;
wire            n16575;
wire            n16576;
wire            n16577;
wire            n16578;
wire            n16579;
wire      [7:0] n1658;
wire      [7:0] n16580;
wire            n16581;
wire            n16582;
wire            n16583;
wire            n16584;
wire            n16585;
wire      [7:0] n16586;
wire            n16587;
wire            n16588;
wire            n16589;
wire      [7:0] n1659;
wire            n16590;
wire            n16591;
wire      [7:0] n16592;
wire            n16593;
wire            n16594;
wire            n16595;
wire            n16596;
wire            n16597;
wire      [7:0] n16598;
wire            n16599;
wire            n166;
wire      [7:0] n1660;
wire            n16600;
wire            n16601;
wire            n16602;
wire            n16603;
wire      [7:0] n16604;
wire            n16605;
wire            n16606;
wire            n16607;
wire            n16608;
wire            n16609;
wire      [7:0] n1661;
wire      [7:0] n16610;
wire            n16611;
wire            n16612;
wire            n16613;
wire            n16614;
wire            n16615;
wire      [7:0] n16616;
wire            n16617;
wire            n16618;
wire            n16619;
wire      [7:0] n1662;
wire            n16620;
wire            n16621;
wire      [7:0] n16622;
wire            n16623;
wire            n16624;
wire            n16625;
wire            n16626;
wire            n16627;
wire      [7:0] n16628;
wire            n16629;
wire      [7:0] n1663;
wire            n16630;
wire            n16631;
wire            n16632;
wire            n16633;
wire      [7:0] n16634;
wire            n16635;
wire            n16636;
wire            n16637;
wire            n16638;
wire            n16639;
wire      [7:0] n1664;
wire      [7:0] n16640;
wire            n16641;
wire            n16642;
wire            n16643;
wire            n16644;
wire            n16645;
wire      [7:0] n16646;
wire            n16647;
wire            n16648;
wire            n16649;
wire      [7:0] n1665;
wire            n16650;
wire            n16651;
wire      [7:0] n16652;
wire            n16653;
wire            n16654;
wire            n16655;
wire            n16656;
wire            n16657;
wire      [7:0] n16658;
wire            n16659;
wire      [7:0] n1666;
wire            n16660;
wire            n16661;
wire            n16662;
wire            n16663;
wire      [7:0] n16664;
wire            n16665;
wire            n16666;
wire            n16667;
wire            n16668;
wire            n16669;
wire      [7:0] n1667;
wire      [7:0] n16670;
wire            n16671;
wire            n16672;
wire            n16673;
wire            n16674;
wire            n16675;
wire      [7:0] n16676;
wire            n16677;
wire            n16678;
wire            n16679;
wire      [7:0] n1668;
wire            n16680;
wire            n16681;
wire      [7:0] n16682;
wire            n16683;
wire            n16684;
wire            n16685;
wire            n16686;
wire            n16687;
wire      [7:0] n16688;
wire            n16689;
wire      [7:0] n1669;
wire            n16690;
wire            n16691;
wire            n16692;
wire            n16693;
wire      [7:0] n16694;
wire            n16695;
wire            n16696;
wire            n16697;
wire            n16698;
wire            n16699;
wire      [7:0] n1670;
wire      [7:0] n16700;
wire            n16701;
wire            n16702;
wire            n16703;
wire            n16704;
wire            n16705;
wire      [7:0] n16706;
wire            n16707;
wire            n16708;
wire            n16709;
wire      [7:0] n1671;
wire            n16710;
wire            n16711;
wire      [7:0] n16712;
wire            n16713;
wire            n16714;
wire            n16715;
wire            n16716;
wire            n16717;
wire      [7:0] n16718;
wire            n16719;
wire      [7:0] n1672;
wire            n16720;
wire            n16721;
wire            n16722;
wire            n16723;
wire      [7:0] n16724;
wire            n16725;
wire            n16726;
wire            n16727;
wire            n16728;
wire            n16729;
wire      [7:0] n1673;
wire      [7:0] n16730;
wire            n16731;
wire            n16732;
wire            n16733;
wire            n16734;
wire            n16735;
wire      [7:0] n16736;
wire            n16737;
wire            n16738;
wire            n16739;
wire      [7:0] n1674;
wire            n16740;
wire            n16741;
wire      [7:0] n16742;
wire            n16743;
wire            n16744;
wire            n16745;
wire            n16746;
wire            n16747;
wire      [7:0] n16748;
wire            n16749;
wire      [7:0] n1675;
wire            n16750;
wire            n16751;
wire            n16752;
wire            n16753;
wire      [7:0] n16754;
wire            n16755;
wire            n16756;
wire            n16757;
wire            n16758;
wire            n16759;
wire      [7:0] n1676;
wire      [7:0] n16760;
wire            n16761;
wire            n16762;
wire            n16763;
wire            n16764;
wire            n16765;
wire      [7:0] n16766;
wire            n16767;
wire            n16768;
wire            n16769;
wire      [7:0] n1677;
wire            n16770;
wire            n16771;
wire      [7:0] n16772;
wire            n16773;
wire            n16774;
wire            n16775;
wire            n16776;
wire            n16777;
wire      [7:0] n16778;
wire            n16779;
wire      [7:0] n1678;
wire            n16780;
wire            n16781;
wire            n16782;
wire            n16783;
wire      [7:0] n16784;
wire            n16785;
wire            n16786;
wire            n16787;
wire            n16788;
wire            n16789;
wire      [7:0] n1679;
wire      [7:0] n16790;
wire            n16791;
wire            n16792;
wire            n16793;
wire            n16794;
wire            n16795;
wire      [7:0] n16796;
wire            n16797;
wire            n16798;
wire            n16799;
wire            n168;
wire      [7:0] n1680;
wire            n16800;
wire            n16801;
wire      [7:0] n16802;
wire            n16803;
wire            n16804;
wire            n16805;
wire            n16806;
wire            n16807;
wire      [7:0] n16808;
wire            n16809;
wire      [7:0] n1681;
wire            n16810;
wire            n16811;
wire            n16812;
wire            n16813;
wire      [7:0] n16814;
wire            n16815;
wire            n16816;
wire            n16817;
wire            n16818;
wire            n16819;
wire      [7:0] n1682;
wire      [7:0] n16820;
wire            n16821;
wire            n16822;
wire            n16823;
wire            n16824;
wire            n16825;
wire      [7:0] n16826;
wire            n16827;
wire            n16828;
wire            n16829;
wire      [7:0] n1683;
wire            n16830;
wire            n16831;
wire      [7:0] n16832;
wire            n16833;
wire            n16834;
wire            n16835;
wire            n16836;
wire            n16837;
wire      [7:0] n16838;
wire            n16839;
wire      [7:0] n1684;
wire            n16840;
wire            n16841;
wire            n16842;
wire            n16843;
wire      [7:0] n16844;
wire            n16845;
wire            n16846;
wire            n16847;
wire            n16848;
wire            n16849;
wire      [7:0] n1685;
wire      [7:0] n16850;
wire            n16851;
wire            n16852;
wire            n16853;
wire            n16854;
wire            n16855;
wire      [7:0] n16856;
wire            n16857;
wire            n16858;
wire            n16859;
wire      [7:0] n1686;
wire            n16860;
wire            n16861;
wire      [7:0] n16862;
wire            n16863;
wire            n16864;
wire            n16865;
wire            n16866;
wire            n16867;
wire      [7:0] n16868;
wire            n16869;
wire      [7:0] n1687;
wire            n16870;
wire            n16871;
wire            n16872;
wire            n16873;
wire      [7:0] n16874;
wire            n16875;
wire            n16876;
wire            n16877;
wire            n16878;
wire            n16879;
wire      [7:0] n1688;
wire      [7:0] n16880;
wire            n16881;
wire            n16882;
wire            n16883;
wire            n16884;
wire            n16885;
wire      [7:0] n16886;
wire            n16887;
wire            n16888;
wire            n16889;
wire      [7:0] n1689;
wire            n16890;
wire            n16891;
wire      [7:0] n16892;
wire            n16893;
wire            n16894;
wire            n16895;
wire            n16896;
wire            n16897;
wire      [7:0] n16898;
wire            n16899;
wire      [7:0] n1690;
wire            n16900;
wire            n16901;
wire            n16902;
wire            n16903;
wire      [7:0] n16904;
wire            n16905;
wire            n16906;
wire            n16907;
wire            n16908;
wire            n16909;
wire      [7:0] n1691;
wire      [7:0] n16910;
wire            n16911;
wire            n16912;
wire            n16913;
wire            n16914;
wire            n16915;
wire      [7:0] n16916;
wire            n16917;
wire            n16918;
wire            n16919;
wire      [7:0] n1692;
wire            n16920;
wire            n16921;
wire      [7:0] n16922;
wire            n16923;
wire            n16924;
wire            n16925;
wire            n16926;
wire            n16927;
wire      [7:0] n16928;
wire            n16929;
wire      [7:0] n1693;
wire            n16930;
wire            n16931;
wire            n16932;
wire            n16933;
wire      [7:0] n16934;
wire            n16935;
wire            n16936;
wire            n16937;
wire            n16938;
wire            n16939;
wire      [7:0] n1694;
wire      [7:0] n16940;
wire            n16941;
wire            n16942;
wire            n16943;
wire            n16944;
wire            n16945;
wire      [7:0] n16946;
wire            n16947;
wire            n16948;
wire            n16949;
wire      [7:0] n1695;
wire            n16950;
wire            n16951;
wire      [7:0] n16952;
wire            n16953;
wire            n16954;
wire            n16955;
wire            n16956;
wire            n16957;
wire      [7:0] n16958;
wire            n16959;
wire      [7:0] n1696;
wire            n16960;
wire            n16961;
wire            n16962;
wire            n16963;
wire      [7:0] n16964;
wire            n16965;
wire            n16966;
wire            n16967;
wire            n16968;
wire            n16969;
wire      [7:0] n1697;
wire      [7:0] n16970;
wire            n16971;
wire            n16972;
wire            n16973;
wire            n16974;
wire            n16975;
wire      [7:0] n16976;
wire            n16977;
wire            n16978;
wire            n16979;
wire      [7:0] n1698;
wire            n16980;
wire            n16981;
wire      [7:0] n16982;
wire            n16983;
wire            n16984;
wire            n16985;
wire            n16986;
wire            n16987;
wire      [7:0] n16988;
wire            n16989;
wire      [7:0] n1699;
wire            n16990;
wire            n16991;
wire            n16992;
wire            n16993;
wire      [7:0] n16994;
wire            n16995;
wire            n16996;
wire            n16997;
wire            n16998;
wire            n16999;
wire            n17;
wire            n170;
wire      [7:0] n1700;
wire      [7:0] n17000;
wire            n17001;
wire            n17002;
wire            n17003;
wire            n17004;
wire            n17005;
wire      [7:0] n17006;
wire            n17007;
wire            n17008;
wire            n17009;
wire      [7:0] n1701;
wire            n17010;
wire            n17011;
wire      [7:0] n17012;
wire            n17013;
wire            n17014;
wire            n17015;
wire            n17016;
wire            n17017;
wire      [7:0] n17018;
wire            n17019;
wire      [7:0] n1702;
wire            n17020;
wire            n17021;
wire            n17022;
wire            n17023;
wire      [7:0] n17024;
wire            n17025;
wire            n17026;
wire            n17027;
wire            n17028;
wire            n17029;
wire      [7:0] n1703;
wire      [7:0] n17030;
wire            n17031;
wire            n17032;
wire            n17033;
wire            n17034;
wire            n17035;
wire      [7:0] n17036;
wire            n17037;
wire            n17038;
wire            n17039;
wire      [7:0] n1704;
wire            n17040;
wire            n17041;
wire      [7:0] n17042;
wire            n17043;
wire            n17044;
wire            n17045;
wire            n17046;
wire            n17047;
wire      [7:0] n17048;
wire            n17049;
wire      [7:0] n1705;
wire            n17050;
wire            n17051;
wire            n17052;
wire            n17053;
wire      [7:0] n17054;
wire            n17055;
wire            n17056;
wire            n17057;
wire            n17058;
wire            n17059;
wire      [7:0] n1706;
wire      [7:0] n17060;
wire            n17061;
wire            n17062;
wire            n17063;
wire            n17064;
wire            n17065;
wire      [7:0] n17066;
wire            n17067;
wire            n17068;
wire            n17069;
wire      [7:0] n1707;
wire            n17070;
wire            n17071;
wire      [7:0] n17072;
wire            n17073;
wire            n17074;
wire            n17075;
wire            n17076;
wire            n17077;
wire      [7:0] n17078;
wire            n17079;
wire      [7:0] n1708;
wire            n17080;
wire            n17081;
wire            n17082;
wire            n17083;
wire      [7:0] n17084;
wire            n17085;
wire            n17086;
wire            n17087;
wire            n17088;
wire            n17089;
wire      [7:0] n1709;
wire      [7:0] n17090;
wire            n17091;
wire            n17092;
wire            n17093;
wire            n17094;
wire            n17095;
wire      [7:0] n17096;
wire            n17097;
wire            n17098;
wire            n17099;
wire      [7:0] n1710;
wire            n17100;
wire            n17101;
wire      [7:0] n17102;
wire            n17103;
wire            n17104;
wire            n17105;
wire            n17106;
wire            n17107;
wire      [7:0] n17108;
wire            n17109;
wire      [7:0] n1711;
wire            n17110;
wire            n17111;
wire            n17112;
wire            n17113;
wire      [7:0] n17114;
wire            n17115;
wire            n17116;
wire            n17117;
wire            n17118;
wire            n17119;
wire      [7:0] n1712;
wire      [7:0] n17120;
wire            n17121;
wire            n17122;
wire            n17123;
wire            n17124;
wire            n17125;
wire      [7:0] n17126;
wire            n17127;
wire            n17128;
wire            n17129;
wire      [7:0] n1713;
wire            n17130;
wire            n17131;
wire      [7:0] n17132;
wire            n17133;
wire            n17134;
wire            n17135;
wire            n17136;
wire            n17137;
wire      [7:0] n17138;
wire            n17139;
wire      [7:0] n1714;
wire            n17140;
wire            n17141;
wire            n17142;
wire            n17143;
wire      [7:0] n17144;
wire            n17145;
wire            n17146;
wire            n17147;
wire            n17148;
wire            n17149;
wire      [7:0] n1715;
wire      [7:0] n17150;
wire            n17151;
wire            n17152;
wire            n17153;
wire            n17154;
wire            n17155;
wire      [7:0] n17156;
wire            n17157;
wire            n17158;
wire            n17159;
wire      [7:0] n1716;
wire            n17160;
wire            n17161;
wire      [7:0] n17162;
wire            n17163;
wire            n17164;
wire            n17165;
wire            n17166;
wire            n17167;
wire      [7:0] n17168;
wire            n17169;
wire      [7:0] n1717;
wire            n17170;
wire            n17171;
wire            n17172;
wire            n17173;
wire      [7:0] n17174;
wire            n17175;
wire            n17176;
wire            n17177;
wire            n17178;
wire            n17179;
wire      [7:0] n1718;
wire      [7:0] n17180;
wire            n17181;
wire            n17182;
wire            n17183;
wire            n17184;
wire            n17185;
wire      [7:0] n17186;
wire            n17187;
wire            n17188;
wire            n17189;
wire      [7:0] n1719;
wire            n17190;
wire            n17191;
wire      [7:0] n17192;
wire            n17193;
wire            n17194;
wire            n17195;
wire            n17196;
wire            n17197;
wire      [7:0] n17198;
wire            n17199;
wire            n172;
wire      [7:0] n1720;
wire            n17200;
wire            n17201;
wire            n17202;
wire            n17203;
wire      [7:0] n17204;
wire            n17205;
wire            n17206;
wire            n17207;
wire            n17208;
wire            n17209;
wire      [7:0] n1721;
wire      [7:0] n17210;
wire            n17211;
wire            n17212;
wire            n17213;
wire            n17214;
wire            n17215;
wire      [7:0] n17216;
wire            n17217;
wire            n17218;
wire            n17219;
wire      [7:0] n1722;
wire            n17220;
wire            n17221;
wire      [7:0] n17222;
wire            n17223;
wire            n17224;
wire            n17225;
wire            n17226;
wire            n17227;
wire      [7:0] n17228;
wire            n17229;
wire      [7:0] n1723;
wire            n17230;
wire            n17231;
wire            n17232;
wire            n17233;
wire      [7:0] n17234;
wire            n17235;
wire            n17236;
wire            n17237;
wire            n17238;
wire            n17239;
wire      [7:0] n1724;
wire      [7:0] n17240;
wire            n17241;
wire            n17242;
wire            n17243;
wire            n17244;
wire            n17245;
wire      [7:0] n17246;
wire            n17247;
wire            n17248;
wire            n17249;
wire      [7:0] n1725;
wire            n17250;
wire            n17251;
wire      [7:0] n17252;
wire            n17253;
wire            n17254;
wire            n17255;
wire            n17256;
wire            n17257;
wire      [7:0] n17258;
wire            n17259;
wire      [7:0] n1726;
wire            n17260;
wire            n17261;
wire            n17262;
wire            n17263;
wire      [7:0] n17264;
wire            n17265;
wire            n17266;
wire            n17267;
wire            n17268;
wire            n17269;
wire      [7:0] n1727;
wire      [7:0] n17270;
wire            n17271;
wire            n17272;
wire            n17273;
wire            n17274;
wire            n17275;
wire      [7:0] n17276;
wire            n17277;
wire            n17278;
wire            n17279;
wire      [7:0] n1728;
wire            n17280;
wire            n17281;
wire      [7:0] n17282;
wire            n17283;
wire            n17284;
wire            n17285;
wire            n17286;
wire            n17287;
wire      [7:0] n17288;
wire            n17289;
wire      [7:0] n1729;
wire            n17290;
wire            n17291;
wire            n17292;
wire            n17293;
wire      [7:0] n17294;
wire            n17295;
wire            n17296;
wire            n17297;
wire            n17298;
wire            n17299;
wire      [7:0] n1730;
wire      [7:0] n17300;
wire            n17301;
wire            n17302;
wire            n17303;
wire            n17304;
wire            n17305;
wire      [7:0] n17306;
wire            n17307;
wire            n17308;
wire            n17309;
wire      [7:0] n1731;
wire            n17310;
wire            n17311;
wire      [7:0] n17312;
wire            n17313;
wire            n17314;
wire            n17315;
wire            n17316;
wire            n17317;
wire      [7:0] n17318;
wire            n17319;
wire      [7:0] n1732;
wire            n17320;
wire            n17321;
wire            n17322;
wire            n17323;
wire      [7:0] n17324;
wire            n17325;
wire            n17326;
wire            n17327;
wire            n17328;
wire            n17329;
wire      [7:0] n1733;
wire      [7:0] n17330;
wire            n17331;
wire            n17332;
wire            n17333;
wire            n17334;
wire            n17335;
wire      [7:0] n17336;
wire            n17337;
wire            n17338;
wire            n17339;
wire      [7:0] n1734;
wire            n17340;
wire            n17341;
wire      [7:0] n17342;
wire            n17343;
wire            n17344;
wire            n17345;
wire            n17346;
wire            n17347;
wire      [7:0] n17348;
wire            n17349;
wire      [7:0] n1735;
wire            n17350;
wire            n17351;
wire            n17352;
wire            n17353;
wire      [7:0] n17354;
wire            n17355;
wire            n17356;
wire            n17357;
wire            n17358;
wire            n17359;
wire      [7:0] n1736;
wire      [7:0] n17360;
wire            n17361;
wire            n17362;
wire            n17363;
wire            n17364;
wire            n17365;
wire      [7:0] n17366;
wire            n17367;
wire            n17368;
wire            n17369;
wire      [7:0] n1737;
wire            n17370;
wire            n17371;
wire      [7:0] n17372;
wire            n17373;
wire            n17374;
wire            n17375;
wire            n17376;
wire            n17377;
wire      [7:0] n17378;
wire            n17379;
wire      [7:0] n1738;
wire            n17380;
wire            n17381;
wire            n17382;
wire            n17383;
wire      [7:0] n17384;
wire            n17385;
wire            n17386;
wire            n17387;
wire            n17388;
wire            n17389;
wire      [7:0] n1739;
wire      [7:0] n17390;
wire            n17391;
wire            n17392;
wire            n17393;
wire            n17394;
wire            n17395;
wire      [7:0] n17396;
wire            n17397;
wire            n17398;
wire            n17399;
wire            n174;
wire      [7:0] n1740;
wire            n17400;
wire            n17401;
wire      [7:0] n17402;
wire            n17403;
wire            n17404;
wire            n17405;
wire            n17406;
wire            n17407;
wire      [7:0] n17408;
wire            n17409;
wire      [7:0] n1741;
wire            n17410;
wire            n17411;
wire            n17412;
wire            n17413;
wire      [7:0] n17414;
wire            n17415;
wire            n17416;
wire            n17417;
wire            n17418;
wire            n17419;
wire      [7:0] n1742;
wire      [7:0] n17420;
wire            n17421;
wire            n17422;
wire            n17423;
wire            n17424;
wire            n17425;
wire      [7:0] n17426;
wire            n17427;
wire            n17428;
wire            n17429;
wire      [7:0] n1743;
wire            n17430;
wire            n17431;
wire      [7:0] n17432;
wire            n17433;
wire            n17434;
wire            n17435;
wire            n17436;
wire            n17437;
wire      [7:0] n17438;
wire            n17439;
wire      [7:0] n1744;
wire            n17440;
wire            n17441;
wire            n17442;
wire            n17443;
wire      [7:0] n17444;
wire            n17445;
wire            n17446;
wire            n17447;
wire            n17448;
wire            n17449;
wire      [7:0] n1745;
wire      [7:0] n17450;
wire            n17451;
wire            n17452;
wire            n17453;
wire            n17454;
wire            n17455;
wire      [7:0] n17456;
wire            n17457;
wire            n17458;
wire            n17459;
wire      [7:0] n1746;
wire            n17460;
wire            n17461;
wire      [7:0] n17462;
wire            n17463;
wire            n17464;
wire            n17465;
wire            n17466;
wire            n17467;
wire      [7:0] n17468;
wire            n17469;
wire      [7:0] n1747;
wire            n17470;
wire            n17471;
wire            n17472;
wire            n17473;
wire      [7:0] n17474;
wire            n17475;
wire            n17476;
wire            n17477;
wire            n17478;
wire            n17479;
wire      [7:0] n1748;
wire      [7:0] n17480;
wire            n17481;
wire            n17482;
wire            n17483;
wire            n17484;
wire            n17485;
wire      [7:0] n17486;
wire            n17487;
wire            n17488;
wire            n17489;
wire      [7:0] n1749;
wire            n17490;
wire            n17491;
wire      [7:0] n17492;
wire            n17493;
wire            n17494;
wire            n17495;
wire            n17496;
wire            n17497;
wire      [7:0] n17498;
wire            n17499;
wire      [7:0] n1750;
wire            n17500;
wire            n17501;
wire            n17502;
wire            n17503;
wire      [7:0] n17504;
wire            n17505;
wire            n17506;
wire            n17507;
wire            n17508;
wire            n17509;
wire      [7:0] n1751;
wire      [7:0] n17510;
wire            n17511;
wire            n17512;
wire            n17513;
wire            n17514;
wire            n17515;
wire      [7:0] n17516;
wire            n17517;
wire            n17518;
wire            n17519;
wire      [7:0] n1752;
wire            n17520;
wire            n17521;
wire      [7:0] n17522;
wire            n17523;
wire            n17524;
wire            n17525;
wire            n17526;
wire            n17527;
wire      [7:0] n17528;
wire            n17529;
wire      [7:0] n1753;
wire            n17530;
wire            n17531;
wire            n17532;
wire            n17533;
wire      [7:0] n17534;
wire            n17535;
wire            n17536;
wire            n17537;
wire            n17538;
wire            n17539;
wire      [7:0] n1754;
wire      [7:0] n17540;
wire            n17541;
wire            n17542;
wire            n17543;
wire            n17544;
wire            n17545;
wire      [7:0] n17546;
wire            n17547;
wire            n17548;
wire            n17549;
wire      [7:0] n1755;
wire            n17550;
wire            n17551;
wire      [7:0] n17552;
wire            n17553;
wire            n17554;
wire            n17555;
wire            n17556;
wire            n17557;
wire      [7:0] n17558;
wire            n17559;
wire      [7:0] n1756;
wire            n17560;
wire            n17561;
wire            n17562;
wire            n17563;
wire      [7:0] n17564;
wire            n17565;
wire            n17566;
wire            n17567;
wire            n17568;
wire            n17569;
wire      [7:0] n1757;
wire      [7:0] n17570;
wire            n17571;
wire            n17572;
wire            n17573;
wire            n17574;
wire            n17575;
wire      [7:0] n17576;
wire            n17577;
wire            n17578;
wire            n17579;
wire      [7:0] n1758;
wire            n17580;
wire            n17581;
wire      [7:0] n17582;
wire            n17583;
wire            n17584;
wire            n17585;
wire            n17586;
wire            n17587;
wire      [7:0] n17588;
wire            n17589;
wire      [7:0] n1759;
wire            n17590;
wire            n17591;
wire            n17592;
wire            n17593;
wire      [7:0] n17594;
wire            n17595;
wire            n17596;
wire            n17597;
wire            n17598;
wire            n17599;
wire            n176;
wire      [7:0] n1760;
wire      [7:0] n17600;
wire            n17601;
wire            n17602;
wire            n17603;
wire            n17604;
wire            n17605;
wire      [7:0] n17606;
wire            n17607;
wire            n17608;
wire            n17609;
wire      [7:0] n1761;
wire            n17610;
wire            n17611;
wire      [7:0] n17612;
wire            n17613;
wire            n17614;
wire            n17615;
wire            n17616;
wire            n17617;
wire      [7:0] n17618;
wire            n17619;
wire      [7:0] n1762;
wire            n17620;
wire            n17621;
wire            n17622;
wire            n17623;
wire      [7:0] n17624;
wire            n17625;
wire            n17626;
wire            n17627;
wire            n17628;
wire            n17629;
wire      [7:0] n1763;
wire      [7:0] n17630;
wire            n17631;
wire            n17632;
wire            n17633;
wire            n17634;
wire            n17635;
wire      [7:0] n17636;
wire            n17637;
wire            n17638;
wire            n17639;
wire      [7:0] n1764;
wire            n17640;
wire            n17641;
wire      [7:0] n17642;
wire            n17643;
wire            n17644;
wire            n17645;
wire            n17646;
wire            n17647;
wire      [7:0] n17648;
wire            n17649;
wire      [7:0] n1765;
wire            n17650;
wire            n17651;
wire            n17652;
wire            n17653;
wire      [7:0] n17654;
wire            n17655;
wire            n17656;
wire            n17657;
wire            n17658;
wire            n17659;
wire      [7:0] n1766;
wire      [7:0] n17660;
wire            n17661;
wire            n17662;
wire            n17663;
wire            n17664;
wire            n17665;
wire      [7:0] n17666;
wire            n17667;
wire            n17668;
wire            n17669;
wire      [7:0] n1767;
wire            n17670;
wire            n17671;
wire      [7:0] n17672;
wire            n17673;
wire            n17674;
wire            n17675;
wire            n17676;
wire            n17677;
wire      [7:0] n17678;
wire            n17679;
wire      [7:0] n1768;
wire            n17680;
wire            n17681;
wire            n17682;
wire            n17683;
wire      [7:0] n17684;
wire            n17685;
wire            n17686;
wire            n17687;
wire            n17688;
wire            n17689;
wire      [7:0] n1769;
wire      [7:0] n17690;
wire            n17691;
wire            n17692;
wire            n17693;
wire            n17694;
wire            n17695;
wire      [7:0] n17696;
wire            n17697;
wire            n17698;
wire            n17699;
wire      [7:0] n1770;
wire            n17700;
wire            n17701;
wire      [7:0] n17702;
wire            n17703;
wire            n17704;
wire            n17705;
wire            n17706;
wire            n17707;
wire      [7:0] n17708;
wire            n17709;
wire      [7:0] n1771;
wire            n17710;
wire            n17711;
wire            n17712;
wire            n17713;
wire      [7:0] n17714;
wire            n17715;
wire            n17716;
wire            n17717;
wire            n17718;
wire            n17719;
wire      [7:0] n1772;
wire      [7:0] n17720;
wire            n17721;
wire            n17722;
wire            n17723;
wire            n17724;
wire            n17725;
wire      [7:0] n17726;
wire            n17727;
wire            n17728;
wire            n17729;
wire      [7:0] n1773;
wire            n17730;
wire            n17731;
wire      [7:0] n17732;
wire            n17733;
wire            n17734;
wire            n17735;
wire            n17736;
wire            n17737;
wire      [7:0] n17738;
wire            n17739;
wire      [7:0] n1774;
wire            n17740;
wire            n17741;
wire            n17742;
wire            n17743;
wire      [7:0] n17744;
wire            n17745;
wire            n17746;
wire            n17747;
wire            n17748;
wire            n17749;
wire      [7:0] n1775;
wire      [7:0] n17750;
wire            n17751;
wire            n17752;
wire            n17753;
wire            n17754;
wire            n17755;
wire      [7:0] n17756;
wire            n17757;
wire            n17758;
wire            n17759;
wire      [7:0] n1776;
wire            n17760;
wire            n17761;
wire      [7:0] n17762;
wire            n17763;
wire            n17764;
wire            n17765;
wire            n17766;
wire            n17767;
wire      [7:0] n17768;
wire            n17769;
wire      [7:0] n1777;
wire            n17770;
wire            n17771;
wire            n17772;
wire            n17773;
wire      [7:0] n17774;
wire            n17775;
wire            n17776;
wire            n17777;
wire            n17778;
wire            n17779;
wire      [7:0] n1778;
wire      [7:0] n17780;
wire            n17781;
wire            n17782;
wire            n17783;
wire            n17784;
wire            n17785;
wire      [7:0] n17786;
wire            n17787;
wire            n17788;
wire            n17789;
wire      [7:0] n1779;
wire            n17790;
wire            n17791;
wire      [7:0] n17792;
wire            n17793;
wire            n17794;
wire            n17795;
wire            n17796;
wire            n17797;
wire      [7:0] n17798;
wire            n17799;
wire            n178;
wire      [7:0] n1780;
wire            n17800;
wire            n17801;
wire            n17802;
wire            n17803;
wire      [7:0] n17804;
wire            n17805;
wire            n17806;
wire            n17807;
wire            n17808;
wire            n17809;
wire      [7:0] n1781;
wire      [7:0] n17810;
wire            n17811;
wire            n17812;
wire            n17813;
wire            n17814;
wire            n17815;
wire      [7:0] n17816;
wire            n17817;
wire            n17818;
wire            n17819;
wire      [7:0] n1782;
wire            n17820;
wire            n17821;
wire      [7:0] n17822;
wire            n17823;
wire            n17824;
wire            n17825;
wire            n17826;
wire            n17827;
wire      [7:0] n17828;
wire            n17829;
wire      [7:0] n1783;
wire            n17830;
wire            n17831;
wire            n17832;
wire            n17833;
wire      [7:0] n17834;
wire            n17835;
wire            n17836;
wire            n17837;
wire            n17838;
wire            n17839;
wire      [7:0] n1784;
wire      [7:0] n17840;
wire            n17841;
wire            n17842;
wire            n17843;
wire            n17844;
wire            n17845;
wire      [7:0] n17846;
wire            n17847;
wire            n17848;
wire            n17849;
wire      [7:0] n1785;
wire            n17850;
wire            n17851;
wire      [7:0] n17852;
wire            n17853;
wire            n17854;
wire            n17855;
wire            n17856;
wire            n17857;
wire      [7:0] n17858;
wire            n17859;
wire      [7:0] n1786;
wire            n17860;
wire            n17861;
wire            n17862;
wire            n17863;
wire      [7:0] n17864;
wire            n17865;
wire            n17866;
wire            n17867;
wire            n17868;
wire            n17869;
wire      [7:0] n1787;
wire      [7:0] n17870;
wire            n17871;
wire            n17872;
wire            n17873;
wire            n17874;
wire            n17875;
wire      [7:0] n17876;
wire            n17877;
wire            n17878;
wire            n17879;
wire      [7:0] n1788;
wire            n17880;
wire            n17881;
wire      [7:0] n17882;
wire            n17883;
wire            n17884;
wire            n17885;
wire            n17886;
wire            n17887;
wire      [7:0] n17888;
wire            n17889;
wire      [7:0] n1789;
wire            n17890;
wire            n17891;
wire            n17892;
wire            n17893;
wire      [7:0] n17894;
wire            n17895;
wire            n17896;
wire            n17897;
wire            n17898;
wire            n17899;
wire      [7:0] n1790;
wire      [7:0] n17900;
wire            n17901;
wire            n17902;
wire            n17903;
wire            n17904;
wire            n17905;
wire      [7:0] n17906;
wire            n17907;
wire            n17908;
wire            n17909;
wire      [7:0] n1791;
wire            n17910;
wire            n17911;
wire      [7:0] n17912;
wire            n17913;
wire            n17914;
wire            n17915;
wire            n17916;
wire            n17917;
wire      [7:0] n17918;
wire            n17919;
wire      [7:0] n1792;
wire            n17920;
wire            n17921;
wire            n17922;
wire            n17923;
wire      [7:0] n17924;
wire            n17925;
wire            n17926;
wire            n17927;
wire            n17928;
wire            n17929;
wire      [7:0] n1793;
wire      [7:0] n17930;
wire            n17931;
wire            n17932;
wire            n17933;
wire            n17934;
wire            n17935;
wire      [7:0] n17936;
wire            n17937;
wire            n17938;
wire            n17939;
wire      [7:0] n1794;
wire            n17940;
wire            n17941;
wire      [7:0] n17942;
wire            n17943;
wire            n17944;
wire            n17945;
wire            n17946;
wire            n17947;
wire      [7:0] n17948;
wire            n17949;
wire      [7:0] n1795;
wire            n17950;
wire            n17951;
wire            n17952;
wire            n17953;
wire      [7:0] n17954;
wire            n17955;
wire            n17956;
wire            n17957;
wire            n17958;
wire            n17959;
wire      [7:0] n1796;
wire      [7:0] n17960;
wire            n17961;
wire            n17962;
wire            n17963;
wire            n17964;
wire            n17965;
wire      [7:0] n17966;
wire            n17967;
wire            n17968;
wire            n17969;
wire      [7:0] n1797;
wire            n17970;
wire            n17971;
wire      [7:0] n17972;
wire            n17973;
wire            n17974;
wire            n17975;
wire            n17976;
wire            n17977;
wire      [7:0] n17978;
wire            n17979;
wire      [7:0] n1798;
wire            n17980;
wire            n17981;
wire            n17982;
wire            n17983;
wire      [7:0] n17984;
wire            n17985;
wire            n17986;
wire            n17987;
wire            n17988;
wire            n17989;
wire      [7:0] n1799;
wire      [7:0] n17990;
wire            n17991;
wire            n17992;
wire            n17993;
wire            n17994;
wire            n17995;
wire      [7:0] n17996;
wire            n17997;
wire            n17998;
wire            n17999;
wire            n180;
wire      [7:0] n1800;
wire            n18000;
wire            n18001;
wire      [7:0] n18002;
wire            n18003;
wire            n18004;
wire            n18005;
wire            n18006;
wire            n18007;
wire      [7:0] n18008;
wire            n18009;
wire      [7:0] n1801;
wire            n18010;
wire            n18011;
wire            n18012;
wire            n18013;
wire      [7:0] n18014;
wire            n18015;
wire            n18016;
wire            n18017;
wire            n18018;
wire            n18019;
wire      [7:0] n1802;
wire      [7:0] n18020;
wire            n18021;
wire            n18022;
wire            n18023;
wire            n18024;
wire            n18025;
wire      [7:0] n18026;
wire            n18027;
wire            n18028;
wire            n18029;
wire      [7:0] n1803;
wire            n18030;
wire            n18031;
wire      [7:0] n18032;
wire            n18033;
wire            n18034;
wire            n18035;
wire            n18036;
wire            n18037;
wire      [7:0] n18038;
wire            n18039;
wire      [7:0] n1804;
wire            n18040;
wire            n18041;
wire            n18042;
wire            n18043;
wire      [7:0] n18044;
wire            n18045;
wire            n18046;
wire            n18047;
wire            n18048;
wire            n18049;
wire      [7:0] n1805;
wire      [7:0] n18050;
wire            n18051;
wire            n18052;
wire            n18053;
wire            n18054;
wire            n18055;
wire      [7:0] n18056;
wire            n18057;
wire            n18058;
wire            n18059;
wire      [7:0] n1806;
wire            n18060;
wire            n18061;
wire      [7:0] n18062;
wire            n18063;
wire            n18064;
wire            n18065;
wire            n18066;
wire            n18067;
wire      [7:0] n18068;
wire            n18069;
wire      [7:0] n1807;
wire            n18070;
wire            n18071;
wire            n18072;
wire            n18073;
wire      [7:0] n18074;
wire            n18075;
wire            n18076;
wire            n18077;
wire            n18078;
wire            n18079;
wire      [7:0] n1808;
wire      [7:0] n18080;
wire            n18081;
wire            n18082;
wire            n18083;
wire            n18084;
wire            n18085;
wire      [7:0] n18086;
wire            n18087;
wire            n18088;
wire            n18089;
wire      [7:0] n1809;
wire            n18090;
wire            n18091;
wire      [7:0] n18092;
wire            n18093;
wire            n18094;
wire            n18095;
wire            n18096;
wire            n18097;
wire      [7:0] n18098;
wire            n18099;
wire      [7:0] n1810;
wire            n18100;
wire            n18101;
wire            n18102;
wire            n18103;
wire      [7:0] n18104;
wire            n18105;
wire            n18106;
wire            n18107;
wire            n18108;
wire            n18109;
wire      [7:0] n1811;
wire      [7:0] n18110;
wire            n18111;
wire            n18112;
wire            n18113;
wire            n18114;
wire            n18115;
wire      [7:0] n18116;
wire            n18117;
wire            n18118;
wire            n18119;
wire      [7:0] n1812;
wire            n18120;
wire            n18121;
wire      [7:0] n18122;
wire            n18123;
wire            n18124;
wire            n18125;
wire            n18126;
wire            n18127;
wire      [7:0] n18128;
wire            n18129;
wire      [7:0] n1813;
wire            n18130;
wire            n18131;
wire            n18132;
wire            n18133;
wire      [7:0] n18134;
wire            n18135;
wire            n18136;
wire            n18137;
wire            n18138;
wire            n18139;
wire      [7:0] n1814;
wire      [7:0] n18140;
wire            n18141;
wire            n18142;
wire            n18143;
wire            n18144;
wire            n18145;
wire      [7:0] n18146;
wire            n18147;
wire            n18148;
wire            n18149;
wire      [7:0] n1815;
wire            n18150;
wire            n18151;
wire      [7:0] n18152;
wire            n18153;
wire            n18154;
wire            n18155;
wire            n18156;
wire            n18157;
wire      [7:0] n18158;
wire            n18159;
wire      [7:0] n1816;
wire            n18160;
wire            n18161;
wire            n18162;
wire            n18163;
wire      [7:0] n18164;
wire            n18165;
wire            n18166;
wire            n18167;
wire            n18168;
wire            n18169;
wire      [7:0] n1817;
wire      [7:0] n18170;
wire            n18171;
wire            n18172;
wire            n18173;
wire            n18174;
wire            n18175;
wire      [7:0] n18176;
wire            n18177;
wire            n18178;
wire            n18179;
wire      [7:0] n1818;
wire            n18180;
wire            n18181;
wire      [7:0] n18182;
wire            n18183;
wire            n18184;
wire            n18185;
wire            n18186;
wire            n18187;
wire      [7:0] n18188;
wire            n18189;
wire      [7:0] n1819;
wire            n18190;
wire            n18191;
wire            n18192;
wire            n18193;
wire      [7:0] n18194;
wire            n18195;
wire            n18196;
wire            n18197;
wire            n18198;
wire            n18199;
wire            n182;
wire      [7:0] n1820;
wire      [7:0] n18200;
wire            n18201;
wire            n18202;
wire            n18203;
wire            n18204;
wire            n18205;
wire      [7:0] n18206;
wire            n18207;
wire            n18208;
wire            n18209;
wire      [7:0] n1821;
wire            n18210;
wire            n18211;
wire      [7:0] n18212;
wire            n18213;
wire            n18214;
wire            n18215;
wire            n18216;
wire            n18217;
wire      [7:0] n18218;
wire            n18219;
wire      [7:0] n1822;
wire            n18220;
wire            n18221;
wire            n18222;
wire            n18223;
wire      [7:0] n18224;
wire            n18225;
wire            n18226;
wire            n18227;
wire            n18228;
wire            n18229;
wire      [7:0] n1823;
wire      [7:0] n18230;
wire            n18231;
wire            n18232;
wire            n18233;
wire            n18234;
wire            n18235;
wire      [7:0] n18236;
wire            n18237;
wire            n18238;
wire            n18239;
wire      [7:0] n1824;
wire            n18240;
wire            n18241;
wire      [7:0] n18242;
wire            n18243;
wire            n18244;
wire            n18245;
wire            n18246;
wire            n18247;
wire      [7:0] n18248;
wire            n18249;
wire      [7:0] n1825;
wire            n18250;
wire            n18251;
wire            n18252;
wire            n18253;
wire      [7:0] n18254;
wire            n18255;
wire            n18256;
wire            n18257;
wire            n18258;
wire            n18259;
wire      [7:0] n1826;
wire      [7:0] n18260;
wire            n18261;
wire            n18262;
wire            n18263;
wire            n18264;
wire            n18265;
wire      [7:0] n18266;
wire            n18267;
wire            n18268;
wire            n18269;
wire      [7:0] n1827;
wire            n18270;
wire            n18271;
wire      [7:0] n18272;
wire            n18273;
wire            n18274;
wire            n18275;
wire            n18276;
wire            n18277;
wire      [7:0] n18278;
wire            n18279;
wire      [7:0] n1828;
wire            n18280;
wire            n18281;
wire            n18282;
wire            n18283;
wire      [7:0] n18284;
wire            n18285;
wire            n18286;
wire            n18287;
wire            n18288;
wire            n18289;
wire      [7:0] n1829;
wire      [7:0] n18290;
wire            n18291;
wire            n18292;
wire            n18293;
wire            n18294;
wire            n18295;
wire      [7:0] n18296;
wire            n18297;
wire            n18298;
wire            n18299;
wire      [7:0] n1830;
wire            n18300;
wire            n18301;
wire      [7:0] n18302;
wire            n18303;
wire            n18304;
wire            n18305;
wire            n18306;
wire            n18307;
wire      [7:0] n18308;
wire            n18309;
wire      [7:0] n1831;
wire            n18310;
wire            n18311;
wire            n18312;
wire            n18313;
wire      [7:0] n18314;
wire            n18315;
wire            n18316;
wire            n18317;
wire            n18318;
wire            n18319;
wire      [7:0] n1832;
wire      [7:0] n18320;
wire            n18321;
wire            n18322;
wire            n18323;
wire            n18324;
wire            n18325;
wire      [7:0] n18326;
wire            n18327;
wire            n18328;
wire            n18329;
wire      [7:0] n1833;
wire            n18330;
wire            n18331;
wire      [7:0] n18332;
wire            n18333;
wire            n18334;
wire            n18335;
wire            n18336;
wire            n18337;
wire      [7:0] n18338;
wire            n18339;
wire      [7:0] n1834;
wire            n18340;
wire            n18341;
wire            n18342;
wire            n18343;
wire      [7:0] n18344;
wire            n18345;
wire            n18346;
wire            n18347;
wire            n18348;
wire            n18349;
wire      [7:0] n1835;
wire      [7:0] n18350;
wire            n18351;
wire            n18352;
wire            n18353;
wire            n18354;
wire            n18355;
wire      [7:0] n18356;
wire            n18357;
wire            n18358;
wire            n18359;
wire      [7:0] n1836;
wire            n18360;
wire            n18361;
wire      [7:0] n18362;
wire            n18363;
wire            n18364;
wire            n18365;
wire            n18366;
wire            n18367;
wire      [7:0] n18368;
wire            n18369;
wire      [7:0] n1837;
wire            n18370;
wire            n18371;
wire            n18372;
wire            n18373;
wire      [7:0] n18374;
wire            n18375;
wire            n18376;
wire            n18377;
wire            n18378;
wire            n18379;
wire      [7:0] n1838;
wire      [7:0] n18380;
wire            n18381;
wire            n18382;
wire            n18383;
wire            n18384;
wire            n18385;
wire      [7:0] n18386;
wire            n18387;
wire            n18388;
wire            n18389;
wire      [7:0] n1839;
wire            n18390;
wire            n18391;
wire      [7:0] n18392;
wire            n18393;
wire            n18394;
wire            n18395;
wire            n18396;
wire            n18397;
wire      [7:0] n18398;
wire            n18399;
wire            n184;
wire      [7:0] n1840;
wire            n18400;
wire            n18401;
wire            n18402;
wire            n18403;
wire      [7:0] n18404;
wire            n18405;
wire            n18406;
wire            n18407;
wire            n18408;
wire            n18409;
wire      [7:0] n1841;
wire      [7:0] n18410;
wire            n18411;
wire            n18412;
wire            n18413;
wire            n18414;
wire            n18415;
wire      [7:0] n18416;
wire            n18417;
wire            n18418;
wire            n18419;
wire      [7:0] n1842;
wire            n18420;
wire            n18421;
wire      [7:0] n18422;
wire            n18423;
wire            n18424;
wire            n18425;
wire            n18426;
wire            n18427;
wire      [7:0] n18428;
wire            n18429;
wire      [7:0] n1843;
wire            n18430;
wire            n18431;
wire            n18432;
wire            n18433;
wire      [7:0] n18434;
wire            n18435;
wire            n18436;
wire            n18437;
wire            n18438;
wire            n18439;
wire      [7:0] n1844;
wire      [7:0] n18440;
wire            n18441;
wire            n18442;
wire            n18443;
wire            n18444;
wire            n18445;
wire      [7:0] n18446;
wire            n18447;
wire            n18448;
wire            n18449;
wire      [7:0] n1845;
wire            n18450;
wire            n18451;
wire      [7:0] n18452;
wire            n18453;
wire            n18454;
wire            n18455;
wire            n18456;
wire            n18457;
wire      [7:0] n18458;
wire            n18459;
wire      [7:0] n1846;
wire            n18460;
wire            n18461;
wire            n18462;
wire            n18463;
wire      [7:0] n18464;
wire            n18465;
wire            n18466;
wire            n18467;
wire            n18468;
wire            n18469;
wire      [7:0] n1847;
wire      [7:0] n18470;
wire            n18471;
wire            n18472;
wire            n18473;
wire            n18474;
wire            n18475;
wire      [7:0] n18476;
wire            n18477;
wire            n18478;
wire            n18479;
wire      [7:0] n1848;
wire            n18480;
wire            n18481;
wire      [7:0] n18482;
wire            n18483;
wire            n18484;
wire            n18485;
wire            n18486;
wire            n18487;
wire      [7:0] n18488;
wire            n18489;
wire      [7:0] n1849;
wire            n18490;
wire            n18491;
wire            n18492;
wire            n18493;
wire      [7:0] n18494;
wire            n18495;
wire            n18496;
wire            n18497;
wire            n18498;
wire            n18499;
wire      [7:0] n1850;
wire      [7:0] n18500;
wire            n18501;
wire            n18502;
wire            n18503;
wire            n18504;
wire            n18505;
wire      [7:0] n18506;
wire            n18507;
wire            n18508;
wire            n18509;
wire      [7:0] n1851;
wire            n18510;
wire            n18511;
wire      [7:0] n18512;
wire            n18513;
wire            n18514;
wire            n18515;
wire            n18516;
wire            n18517;
wire      [7:0] n18518;
wire            n18519;
wire      [7:0] n1852;
wire            n18520;
wire            n18521;
wire            n18522;
wire            n18523;
wire      [7:0] n18524;
wire            n18525;
wire            n18526;
wire            n18527;
wire            n18528;
wire            n18529;
wire      [7:0] n1853;
wire      [7:0] n18530;
wire            n18531;
wire            n18532;
wire            n18533;
wire            n18534;
wire            n18535;
wire      [7:0] n18536;
wire            n18537;
wire            n18538;
wire            n18539;
wire      [7:0] n1854;
wire            n18540;
wire            n18541;
wire      [7:0] n18542;
wire            n18543;
wire            n18544;
wire            n18545;
wire            n18546;
wire            n18547;
wire      [7:0] n18548;
wire            n18549;
wire      [7:0] n1855;
wire            n18550;
wire            n18551;
wire            n18552;
wire            n18553;
wire      [7:0] n18554;
wire            n18555;
wire            n18556;
wire            n18557;
wire            n18558;
wire            n18559;
wire      [7:0] n1856;
wire      [7:0] n18560;
wire            n18561;
wire            n18562;
wire            n18563;
wire            n18564;
wire            n18565;
wire      [7:0] n18566;
wire            n18567;
wire            n18568;
wire            n18569;
wire      [7:0] n1857;
wire            n18570;
wire            n18571;
wire      [7:0] n18572;
wire            n18573;
wire            n18574;
wire            n18575;
wire            n18576;
wire            n18577;
wire      [7:0] n18578;
wire            n18579;
wire      [7:0] n1858;
wire            n18580;
wire            n18581;
wire            n18582;
wire            n18583;
wire      [7:0] n18584;
wire            n18585;
wire            n18586;
wire            n18587;
wire            n18588;
wire            n18589;
wire      [7:0] n1859;
wire      [7:0] n18590;
wire            n18591;
wire            n18592;
wire            n18593;
wire            n18594;
wire            n18595;
wire      [7:0] n18596;
wire            n18597;
wire            n18598;
wire            n18599;
wire            n186;
wire      [7:0] n1860;
wire            n18600;
wire            n18601;
wire      [7:0] n18602;
wire            n18603;
wire            n18604;
wire            n18605;
wire            n18606;
wire            n18607;
wire      [7:0] n18608;
wire            n18609;
wire      [7:0] n1861;
wire            n18610;
wire            n18611;
wire            n18612;
wire            n18613;
wire      [7:0] n18614;
wire            n18615;
wire            n18616;
wire            n18617;
wire            n18618;
wire            n18619;
wire      [7:0] n1862;
wire      [7:0] n18620;
wire            n18621;
wire            n18622;
wire            n18623;
wire            n18624;
wire            n18625;
wire      [7:0] n18626;
wire            n18627;
wire            n18628;
wire            n18629;
wire      [7:0] n1863;
wire            n18630;
wire            n18631;
wire      [7:0] n18632;
wire            n18633;
wire            n18634;
wire            n18635;
wire            n18636;
wire            n18637;
wire      [7:0] n18638;
wire            n18639;
wire      [7:0] n1864;
wire            n18640;
wire            n18641;
wire            n18642;
wire            n18643;
wire      [7:0] n18644;
wire            n18645;
wire            n18646;
wire            n18647;
wire            n18648;
wire            n18649;
wire            n1865;
wire      [7:0] n18650;
wire            n18651;
wire            n18652;
wire            n18653;
wire            n18654;
wire            n18655;
wire      [7:0] n18656;
wire            n18657;
wire            n18658;
wire            n18659;
wire            n1866;
wire            n18660;
wire            n18661;
wire      [7:0] n18662;
wire            n18663;
wire            n18664;
wire            n18665;
wire            n18666;
wire            n18667;
wire      [7:0] n18668;
wire            n18669;
wire      [3:0] n1867;
wire            n18670;
wire            n18671;
wire            n18672;
wire            n18673;
wire      [7:0] n18674;
wire            n18675;
wire            n18676;
wire            n18677;
wire            n18678;
wire            n18679;
wire      [4:0] n1868;
wire      [7:0] n18680;
wire            n18681;
wire            n18682;
wire            n18683;
wire            n18684;
wire            n18685;
wire      [7:0] n18686;
wire            n18687;
wire            n18688;
wire            n18689;
wire      [7:0] n1869;
wire            n18690;
wire            n18691;
wire      [7:0] n18692;
wire            n18693;
wire            n18694;
wire            n18695;
wire            n18696;
wire            n18697;
wire      [7:0] n18698;
wire            n18699;
wire      [3:0] n1870;
wire            n18700;
wire            n18701;
wire            n18702;
wire            n18703;
wire      [7:0] n18704;
wire            n18705;
wire            n18706;
wire            n18707;
wire            n18708;
wire            n18709;
wire      [7:0] n1871;
wire      [7:0] n18710;
wire            n18711;
wire            n18712;
wire            n18713;
wire            n18714;
wire            n18715;
wire      [7:0] n18716;
wire            n18717;
wire            n18718;
wire            n18719;
wire      [7:0] n1872;
wire            n18720;
wire            n18721;
wire      [7:0] n18722;
wire            n18723;
wire            n18724;
wire            n18725;
wire            n18726;
wire            n18727;
wire      [7:0] n18728;
wire            n18729;
wire      [7:0] n1873;
wire            n18730;
wire            n18731;
wire            n18732;
wire            n18733;
wire      [7:0] n18734;
wire            n18735;
wire            n18736;
wire            n18737;
wire            n18738;
wire            n18739;
wire      [7:0] n1874;
wire      [7:0] n18740;
wire            n18741;
wire            n18742;
wire            n18743;
wire            n18744;
wire            n18745;
wire      [7:0] n18746;
wire            n18747;
wire            n18748;
wire            n18749;
wire            n1875;
wire            n18750;
wire            n18751;
wire      [7:0] n18752;
wire            n18753;
wire            n18754;
wire            n18755;
wire            n18756;
wire            n18757;
wire      [7:0] n18758;
wire            n18759;
wire            n1876;
wire            n18760;
wire            n18761;
wire            n18762;
wire            n18763;
wire      [7:0] n18764;
wire            n18765;
wire            n18766;
wire            n18767;
wire            n18768;
wire            n18769;
wire            n1877;
wire      [7:0] n18770;
wire            n18771;
wire            n18772;
wire            n18773;
wire            n18774;
wire            n18775;
wire      [7:0] n18776;
wire            n18777;
wire            n18778;
wire            n18779;
wire            n1878;
wire            n18780;
wire            n18781;
wire      [7:0] n18782;
wire            n18783;
wire            n18784;
wire            n18785;
wire            n18786;
wire            n18787;
wire      [7:0] n18788;
wire            n18789;
wire            n1879;
wire            n18790;
wire            n18791;
wire            n18792;
wire            n18793;
wire      [7:0] n18794;
wire            n18795;
wire            n18796;
wire            n18797;
wire            n18798;
wire            n18799;
wire            n188;
wire            n1880;
wire      [7:0] n18800;
wire            n18801;
wire            n18802;
wire            n18803;
wire            n18804;
wire            n18805;
wire      [7:0] n18806;
wire            n18807;
wire            n18808;
wire            n18809;
wire            n1881;
wire            n18810;
wire            n18811;
wire      [7:0] n18812;
wire            n18813;
wire            n18814;
wire            n18815;
wire            n18816;
wire            n18817;
wire      [7:0] n18818;
wire            n18819;
wire            n1882;
wire            n18820;
wire            n18821;
wire            n18822;
wire            n18823;
wire      [7:0] n18824;
wire            n18825;
wire            n18826;
wire            n18827;
wire            n18828;
wire            n18829;
wire            n1883;
wire      [7:0] n18830;
wire            n18831;
wire            n18832;
wire            n18833;
wire            n18834;
wire            n18835;
wire      [7:0] n18836;
wire            n18837;
wire            n18838;
wire            n18839;
wire            n1884;
wire            n18840;
wire            n18841;
wire      [7:0] n18842;
wire            n18843;
wire            n18844;
wire            n18845;
wire            n18846;
wire            n18847;
wire      [7:0] n18848;
wire            n18849;
wire            n1885;
wire            n18850;
wire            n18851;
wire            n18852;
wire            n18853;
wire      [7:0] n18854;
wire            n18855;
wire            n18856;
wire            n18857;
wire            n18858;
wire            n18859;
wire            n1886;
wire      [7:0] n18860;
wire            n18861;
wire            n18862;
wire            n18863;
wire            n18864;
wire            n18865;
wire      [7:0] n18866;
wire            n18867;
wire            n18868;
wire            n18869;
wire            n1887;
wire            n18870;
wire            n18871;
wire      [7:0] n18872;
wire            n18873;
wire            n18874;
wire            n18875;
wire            n18876;
wire            n18877;
wire      [7:0] n18878;
wire            n18879;
wire            n1888;
wire            n18880;
wire            n18881;
wire            n18882;
wire            n18883;
wire      [7:0] n18884;
wire            n18885;
wire            n18886;
wire            n18887;
wire            n18888;
wire            n18889;
wire            n1889;
wire      [7:0] n18890;
wire            n18891;
wire            n18892;
wire            n18893;
wire            n18894;
wire            n18895;
wire      [7:0] n18896;
wire            n18897;
wire            n18898;
wire            n18899;
wire            n1890;
wire            n18900;
wire            n18901;
wire      [7:0] n18902;
wire            n18903;
wire            n18904;
wire            n18905;
wire            n18906;
wire            n18907;
wire      [7:0] n18908;
wire            n18909;
wire            n1891;
wire            n18910;
wire            n18911;
wire            n18912;
wire            n18913;
wire      [7:0] n18914;
wire            n18915;
wire            n18916;
wire            n18917;
wire            n18918;
wire            n18919;
wire            n1892;
wire      [7:0] n18920;
wire            n18921;
wire            n18922;
wire            n18923;
wire            n18924;
wire            n18925;
wire      [7:0] n18926;
wire            n18927;
wire            n18928;
wire            n18929;
wire            n1893;
wire            n18930;
wire            n18931;
wire      [7:0] n18932;
wire            n18933;
wire            n18934;
wire            n18935;
wire            n18936;
wire            n18937;
wire      [7:0] n18938;
wire            n18939;
wire            n1894;
wire            n18940;
wire            n18941;
wire            n18942;
wire            n18943;
wire      [7:0] n18944;
wire            n18945;
wire            n18946;
wire            n18947;
wire            n18948;
wire            n18949;
wire            n1895;
wire      [7:0] n18950;
wire            n18951;
wire            n18952;
wire            n18953;
wire            n18954;
wire            n18955;
wire      [7:0] n18956;
wire            n18957;
wire            n18958;
wire            n18959;
wire            n1896;
wire            n18960;
wire            n18961;
wire      [7:0] n18962;
wire            n18963;
wire            n18964;
wire            n18965;
wire            n18966;
wire            n18967;
wire      [7:0] n18968;
wire            n18969;
wire            n1897;
wire            n18970;
wire            n18971;
wire            n18972;
wire            n18973;
wire      [7:0] n18974;
wire            n18975;
wire            n18976;
wire            n18977;
wire            n18978;
wire            n18979;
wire            n1898;
wire      [7:0] n18980;
wire            n18981;
wire            n18982;
wire            n18983;
wire            n18984;
wire            n18985;
wire      [7:0] n18986;
wire            n18987;
wire            n18988;
wire            n18989;
wire            n1899;
wire            n18990;
wire            n18991;
wire      [7:0] n18992;
wire            n18993;
wire            n18994;
wire            n18995;
wire            n18996;
wire            n18997;
wire      [7:0] n18998;
wire            n18999;
wire            n19;
wire            n190;
wire            n1900;
wire            n19000;
wire            n19001;
wire            n19002;
wire            n19003;
wire      [7:0] n19004;
wire            n19005;
wire            n19006;
wire            n19007;
wire            n19008;
wire            n19009;
wire            n1901;
wire      [7:0] n19010;
wire            n19011;
wire            n19012;
wire            n19013;
wire            n19014;
wire            n19015;
wire      [7:0] n19016;
wire            n19017;
wire            n19018;
wire            n19019;
wire            n1902;
wire            n19020;
wire            n19021;
wire      [7:0] n19022;
wire            n19023;
wire            n19024;
wire            n19025;
wire            n19026;
wire            n19027;
wire      [7:0] n19028;
wire            n19029;
wire            n1903;
wire            n19030;
wire            n19031;
wire            n19032;
wire            n19033;
wire      [7:0] n19034;
wire            n19035;
wire            n19036;
wire            n19037;
wire            n19038;
wire            n19039;
wire            n1904;
wire      [7:0] n19040;
wire            n19041;
wire            n19042;
wire            n19043;
wire            n19044;
wire            n19045;
wire      [7:0] n19046;
wire            n19047;
wire            n19048;
wire            n19049;
wire            n1905;
wire            n19050;
wire            n19051;
wire      [7:0] n19052;
wire            n19053;
wire            n19054;
wire            n19055;
wire            n19056;
wire            n19057;
wire      [7:0] n19058;
wire            n19059;
wire            n1906;
wire            n19060;
wire            n19061;
wire            n19062;
wire            n19063;
wire      [7:0] n19064;
wire            n19065;
wire            n19066;
wire            n19067;
wire            n19068;
wire            n19069;
wire            n1907;
wire      [7:0] n19070;
wire            n19071;
wire            n19072;
wire            n19073;
wire            n19074;
wire            n19075;
wire      [7:0] n19076;
wire            n19077;
wire            n19078;
wire            n19079;
wire            n1908;
wire            n19080;
wire            n19081;
wire      [7:0] n19082;
wire            n19083;
wire            n19084;
wire            n19085;
wire            n19086;
wire            n19087;
wire      [7:0] n19088;
wire            n19089;
wire            n1909;
wire            n19090;
wire            n19091;
wire            n19092;
wire            n19093;
wire      [7:0] n19094;
wire            n19095;
wire            n19096;
wire            n19097;
wire            n19098;
wire            n19099;
wire            n1910;
wire      [7:0] n19100;
wire            n19101;
wire            n19102;
wire            n19103;
wire            n19104;
wire            n19105;
wire      [7:0] n19106;
wire            n19107;
wire            n19108;
wire            n19109;
wire            n1911;
wire            n19110;
wire            n19111;
wire      [7:0] n19112;
wire            n19113;
wire            n19114;
wire            n19115;
wire            n19116;
wire            n19117;
wire      [7:0] n19118;
wire            n19119;
wire            n1912;
wire            n19120;
wire            n19121;
wire            n19122;
wire            n19123;
wire      [7:0] n19124;
wire            n19125;
wire            n19126;
wire            n19127;
wire            n19128;
wire            n19129;
wire            n1913;
wire      [7:0] n19130;
wire            n19131;
wire            n19132;
wire            n19133;
wire            n19134;
wire            n19135;
wire      [7:0] n19136;
wire            n19137;
wire            n19138;
wire            n19139;
wire            n1914;
wire            n19140;
wire            n19141;
wire      [7:0] n19142;
wire            n19143;
wire            n19144;
wire            n19145;
wire            n19146;
wire            n19147;
wire      [7:0] n19148;
wire            n19149;
wire            n1915;
wire            n19150;
wire            n19151;
wire            n19152;
wire            n19153;
wire      [7:0] n19154;
wire            n19155;
wire            n19156;
wire            n19157;
wire            n19158;
wire            n19159;
wire            n1916;
wire      [7:0] n19160;
wire            n19161;
wire            n19162;
wire            n19163;
wire            n19164;
wire            n19165;
wire      [7:0] n19166;
wire            n19167;
wire            n19168;
wire            n19169;
wire            n1917;
wire            n19170;
wire            n19171;
wire      [7:0] n19172;
wire            n19173;
wire            n19174;
wire            n19175;
wire            n19176;
wire            n19177;
wire      [7:0] n19178;
wire            n19179;
wire            n1918;
wire            n19180;
wire            n19181;
wire            n19182;
wire            n19183;
wire      [7:0] n19184;
wire            n19185;
wire            n19186;
wire            n19187;
wire            n19188;
wire            n19189;
wire            n1919;
wire      [7:0] n19190;
wire            n19191;
wire            n19192;
wire            n19193;
wire            n19194;
wire            n19195;
wire      [7:0] n19196;
wire            n19197;
wire            n19198;
wire            n19199;
wire            n192;
wire            n1920;
wire            n19200;
wire            n19201;
wire      [7:0] n19202;
wire            n19203;
wire            n19204;
wire            n19205;
wire            n19206;
wire            n19207;
wire      [7:0] n19208;
wire            n19209;
wire            n1921;
wire            n19210;
wire            n19211;
wire            n19212;
wire            n19213;
wire      [7:0] n19214;
wire            n19215;
wire            n19216;
wire            n19217;
wire            n19218;
wire            n19219;
wire            n1922;
wire      [7:0] n19220;
wire            n19221;
wire            n19222;
wire            n19223;
wire            n19224;
wire            n19225;
wire      [7:0] n19226;
wire            n19227;
wire            n19228;
wire            n19229;
wire            n1923;
wire            n19230;
wire            n19231;
wire      [7:0] n19232;
wire            n19233;
wire            n19234;
wire            n19235;
wire            n19236;
wire            n19237;
wire      [7:0] n19238;
wire            n19239;
wire            n1924;
wire            n19240;
wire            n19241;
wire            n19242;
wire            n19243;
wire      [7:0] n19244;
wire            n19245;
wire            n19246;
wire            n19247;
wire            n19248;
wire            n19249;
wire            n1925;
wire      [7:0] n19250;
wire            n19251;
wire            n19252;
wire            n19253;
wire            n19254;
wire            n19255;
wire      [7:0] n19256;
wire            n19257;
wire            n19258;
wire            n19259;
wire            n1926;
wire            n19260;
wire            n19261;
wire      [7:0] n19262;
wire            n19263;
wire            n19264;
wire            n19265;
wire            n19266;
wire            n19267;
wire      [7:0] n19268;
wire            n19269;
wire            n1927;
wire            n19270;
wire            n19271;
wire            n19272;
wire            n19273;
wire      [7:0] n19274;
wire            n19275;
wire            n19276;
wire            n19277;
wire            n19278;
wire            n19279;
wire            n1928;
wire      [7:0] n19280;
wire            n19281;
wire            n19282;
wire            n19283;
wire            n19284;
wire            n19285;
wire      [7:0] n19286;
wire            n19287;
wire            n19288;
wire            n19289;
wire            n1929;
wire            n19290;
wire            n19291;
wire      [7:0] n19292;
wire            n19293;
wire            n19294;
wire            n19295;
wire            n19296;
wire            n19297;
wire      [7:0] n19298;
wire            n19299;
wire            n1930;
wire            n19300;
wire            n19301;
wire            n19302;
wire            n19303;
wire      [7:0] n19304;
wire            n19305;
wire            n19306;
wire            n19307;
wire            n19308;
wire            n19309;
wire            n1931;
wire      [7:0] n19310;
wire            n19311;
wire            n19312;
wire            n19313;
wire            n19314;
wire            n19315;
wire      [7:0] n19316;
wire            n19317;
wire            n19318;
wire            n19319;
wire            n1932;
wire            n19320;
wire            n19321;
wire      [7:0] n19322;
wire            n19323;
wire            n19324;
wire            n19325;
wire            n19326;
wire            n19327;
wire      [7:0] n19328;
wire            n19329;
wire            n1933;
wire            n19330;
wire            n19331;
wire            n19332;
wire            n19333;
wire      [7:0] n19334;
wire            n19335;
wire            n19336;
wire            n19337;
wire            n19338;
wire            n19339;
wire            n1934;
wire      [7:0] n19340;
wire            n19341;
wire            n19342;
wire            n19343;
wire            n19344;
wire            n19345;
wire      [7:0] n19346;
wire            n19347;
wire            n19348;
wire            n19349;
wire            n1935;
wire            n19350;
wire            n19351;
wire      [7:0] n19352;
wire            n19353;
wire            n19354;
wire            n19355;
wire            n19356;
wire            n19357;
wire      [7:0] n19358;
wire            n19359;
wire            n1936;
wire            n19360;
wire            n19361;
wire            n19362;
wire            n19363;
wire      [7:0] n19364;
wire            n19365;
wire            n19366;
wire            n19367;
wire            n19368;
wire            n19369;
wire            n1937;
wire      [7:0] n19370;
wire            n19371;
wire            n19372;
wire            n19373;
wire            n19374;
wire            n19375;
wire      [7:0] n19376;
wire            n19377;
wire            n19378;
wire            n19379;
wire            n1938;
wire            n19380;
wire            n19381;
wire      [7:0] n19382;
wire            n19383;
wire            n19384;
wire            n19385;
wire            n19386;
wire            n19387;
wire      [7:0] n19388;
wire            n19389;
wire            n1939;
wire            n19390;
wire            n19391;
wire            n19392;
wire            n19393;
wire      [7:0] n19394;
wire            n19395;
wire            n19396;
wire            n19397;
wire            n19398;
wire            n19399;
wire            n194;
wire            n1940;
wire      [7:0] n19400;
wire            n19401;
wire            n19402;
wire            n19403;
wire            n19404;
wire            n19405;
wire      [7:0] n19406;
wire            n19407;
wire            n19408;
wire            n19409;
wire            n1941;
wire            n19410;
wire            n19411;
wire      [7:0] n19412;
wire            n19413;
wire            n19414;
wire            n19415;
wire            n19416;
wire            n19417;
wire      [7:0] n19418;
wire            n19419;
wire            n1942;
wire            n19420;
wire            n19421;
wire            n19422;
wire            n19423;
wire      [7:0] n19424;
wire            n19425;
wire            n19426;
wire            n19427;
wire            n19428;
wire            n19429;
wire            n1943;
wire      [7:0] n19430;
wire            n19431;
wire            n19432;
wire            n19433;
wire            n19434;
wire            n19435;
wire      [7:0] n19436;
wire            n19437;
wire            n19438;
wire            n19439;
wire            n1944;
wire            n19440;
wire            n19441;
wire      [7:0] n19442;
wire            n19443;
wire            n19444;
wire            n19445;
wire            n19446;
wire            n19447;
wire      [7:0] n19448;
wire            n19449;
wire            n1945;
wire            n19450;
wire            n19451;
wire            n19452;
wire            n19453;
wire      [7:0] n19454;
wire            n19455;
wire            n19456;
wire            n19457;
wire            n19458;
wire            n19459;
wire            n1946;
wire      [7:0] n19460;
wire            n19461;
wire            n19462;
wire            n19463;
wire            n19464;
wire            n19465;
wire      [7:0] n19466;
wire            n19467;
wire            n19468;
wire            n19469;
wire            n1947;
wire            n19470;
wire            n19471;
wire      [7:0] n19472;
wire            n19473;
wire            n19474;
wire            n19475;
wire            n19476;
wire            n19477;
wire      [7:0] n19478;
wire            n19479;
wire            n1948;
wire            n19480;
wire            n19481;
wire            n19482;
wire            n19483;
wire      [7:0] n19484;
wire            n19485;
wire            n19486;
wire            n19487;
wire            n19488;
wire            n19489;
wire            n1949;
wire      [7:0] n19490;
wire            n19491;
wire            n19492;
wire            n19493;
wire            n19494;
wire            n19495;
wire      [7:0] n19496;
wire            n19497;
wire            n19498;
wire            n19499;
wire            n1950;
wire            n19500;
wire            n19501;
wire      [7:0] n19502;
wire            n19503;
wire            n19504;
wire            n19505;
wire            n19506;
wire            n19507;
wire      [7:0] n19508;
wire            n19509;
wire            n1951;
wire            n19510;
wire            n19511;
wire            n19512;
wire            n19513;
wire      [7:0] n19514;
wire            n19515;
wire            n19516;
wire            n19517;
wire            n19518;
wire            n19519;
wire            n1952;
wire      [7:0] n19520;
wire            n19521;
wire            n19522;
wire            n19523;
wire            n19524;
wire            n19525;
wire      [7:0] n19526;
wire            n19527;
wire            n19528;
wire            n19529;
wire            n1953;
wire            n19530;
wire            n19531;
wire      [7:0] n19532;
wire            n19533;
wire            n19534;
wire            n19535;
wire            n19536;
wire            n19537;
wire      [7:0] n19538;
wire            n19539;
wire            n1954;
wire            n19540;
wire            n19541;
wire            n19542;
wire            n19543;
wire      [7:0] n19544;
wire            n19545;
wire            n19546;
wire            n19547;
wire            n19548;
wire            n19549;
wire            n1955;
wire      [7:0] n19550;
wire            n19551;
wire            n19552;
wire            n19553;
wire            n19554;
wire            n19555;
wire      [7:0] n19556;
wire            n19557;
wire            n19558;
wire            n19559;
wire            n1956;
wire            n19560;
wire            n19561;
wire      [7:0] n19562;
wire            n19563;
wire            n19564;
wire            n19565;
wire            n19566;
wire            n19567;
wire      [7:0] n19568;
wire            n19569;
wire            n1957;
wire            n19570;
wire            n19571;
wire            n19572;
wire            n19573;
wire      [7:0] n19574;
wire            n19575;
wire            n19576;
wire            n19577;
wire            n19578;
wire            n19579;
wire            n1958;
wire      [7:0] n19580;
wire            n19581;
wire            n19582;
wire            n19583;
wire            n19584;
wire            n19585;
wire      [7:0] n19586;
wire            n19587;
wire            n19588;
wire            n19589;
wire            n1959;
wire            n19590;
wire            n19591;
wire      [7:0] n19592;
wire            n19593;
wire            n19594;
wire            n19595;
wire            n19596;
wire            n19597;
wire      [7:0] n19598;
wire            n19599;
wire            n196;
wire            n1960;
wire            n19600;
wire            n19601;
wire            n19602;
wire            n19603;
wire      [7:0] n19604;
wire            n19605;
wire            n19606;
wire            n19607;
wire            n19608;
wire            n19609;
wire            n1961;
wire      [7:0] n19610;
wire            n19611;
wire            n19612;
wire            n19613;
wire            n19614;
wire            n19615;
wire      [7:0] n19616;
wire            n19617;
wire            n19618;
wire            n19619;
wire            n1962;
wire            n19620;
wire            n19621;
wire      [7:0] n19622;
wire            n19623;
wire            n19624;
wire            n19625;
wire            n19626;
wire            n19627;
wire      [7:0] n19628;
wire            n19629;
wire            n1963;
wire            n19630;
wire            n19631;
wire            n19632;
wire            n19633;
wire      [7:0] n19634;
wire            n19635;
wire            n19636;
wire            n19637;
wire            n19638;
wire            n19639;
wire            n1964;
wire      [7:0] n19640;
wire            n19641;
wire            n19642;
wire            n19643;
wire            n19644;
wire            n19645;
wire      [7:0] n19646;
wire            n19647;
wire            n19648;
wire            n19649;
wire            n1965;
wire            n19650;
wire            n19651;
wire      [7:0] n19652;
wire            n19653;
wire            n19654;
wire            n19655;
wire            n19656;
wire            n19657;
wire      [7:0] n19658;
wire            n19659;
wire            n1966;
wire            n19660;
wire            n19661;
wire            n19662;
wire            n19663;
wire      [7:0] n19664;
wire            n19665;
wire            n19666;
wire            n19667;
wire            n19668;
wire            n19669;
wire            n1967;
wire      [7:0] n19670;
wire            n19671;
wire            n19672;
wire            n19673;
wire            n19674;
wire            n19675;
wire      [7:0] n19676;
wire            n19677;
wire            n19678;
wire            n19679;
wire            n1968;
wire            n19680;
wire            n19681;
wire      [7:0] n19682;
wire            n19683;
wire            n19684;
wire            n19685;
wire            n19686;
wire            n19687;
wire      [7:0] n19688;
wire            n19689;
wire            n1969;
wire            n19690;
wire            n19691;
wire            n19692;
wire            n19693;
wire      [7:0] n19694;
wire            n19695;
wire            n19696;
wire            n19697;
wire            n19698;
wire            n19699;
wire            n1970;
wire      [7:0] n19700;
wire            n19701;
wire            n19702;
wire            n19703;
wire            n19704;
wire            n19705;
wire      [7:0] n19706;
wire            n19707;
wire            n19708;
wire            n19709;
wire            n1971;
wire            n19710;
wire            n19711;
wire      [7:0] n19712;
wire            n19713;
wire            n19714;
wire            n19715;
wire            n19716;
wire            n19717;
wire      [7:0] n19718;
wire            n19719;
wire            n1972;
wire            n19720;
wire            n19721;
wire            n19722;
wire            n19723;
wire      [7:0] n19724;
wire            n19725;
wire            n19726;
wire            n19727;
wire            n19728;
wire            n19729;
wire            n1973;
wire      [7:0] n19730;
wire            n19731;
wire            n19732;
wire            n19733;
wire            n19734;
wire            n19735;
wire      [7:0] n19736;
wire            n19737;
wire            n19738;
wire            n19739;
wire            n1974;
wire            n19740;
wire            n19741;
wire      [7:0] n19742;
wire            n19743;
wire            n19744;
wire            n19745;
wire            n19746;
wire            n19747;
wire      [7:0] n19748;
wire            n19749;
wire            n1975;
wire            n19750;
wire            n19751;
wire            n19752;
wire            n19753;
wire      [7:0] n19754;
wire            n19755;
wire            n19756;
wire            n19757;
wire            n19758;
wire            n19759;
wire            n1976;
wire      [7:0] n19760;
wire            n19761;
wire            n19762;
wire            n19763;
wire            n19764;
wire            n19765;
wire      [7:0] n19766;
wire            n19767;
wire            n19768;
wire            n19769;
wire            n1977;
wire            n19770;
wire            n19771;
wire      [7:0] n19772;
wire            n19773;
wire            n19774;
wire            n19775;
wire            n19776;
wire            n19777;
wire      [7:0] n19778;
wire            n19779;
wire            n1978;
wire            n19780;
wire            n19781;
wire            n19782;
wire            n19783;
wire      [7:0] n19784;
wire            n19785;
wire            n19786;
wire            n19787;
wire            n19788;
wire            n19789;
wire            n1979;
wire      [7:0] n19790;
wire            n19791;
wire            n19792;
wire            n19793;
wire            n19794;
wire            n19795;
wire      [7:0] n19796;
wire            n19797;
wire            n19798;
wire            n19799;
wire            n198;
wire            n1980;
wire            n19800;
wire            n19801;
wire      [7:0] n19802;
wire            n19803;
wire            n19804;
wire            n19805;
wire            n19806;
wire            n19807;
wire      [7:0] n19808;
wire            n19809;
wire            n1981;
wire            n19810;
wire            n19811;
wire            n19812;
wire            n19813;
wire      [7:0] n19814;
wire            n19815;
wire            n19816;
wire            n19817;
wire            n19818;
wire            n19819;
wire            n1982;
wire      [7:0] n19820;
wire            n19821;
wire            n19822;
wire            n19823;
wire            n19824;
wire            n19825;
wire      [7:0] n19826;
wire            n19827;
wire            n19828;
wire            n19829;
wire            n1983;
wire            n19830;
wire            n19831;
wire      [7:0] n19832;
wire            n19833;
wire            n19834;
wire            n19835;
wire            n19836;
wire            n19837;
wire      [7:0] n19838;
wire            n19839;
wire            n1984;
wire            n19840;
wire            n19841;
wire            n19842;
wire            n19843;
wire      [7:0] n19844;
wire            n19845;
wire            n19846;
wire            n19847;
wire            n19848;
wire            n19849;
wire            n1985;
wire      [7:0] n19850;
wire            n19851;
wire            n19852;
wire            n19853;
wire            n19854;
wire            n19855;
wire      [7:0] n19856;
wire            n19857;
wire            n19858;
wire            n19859;
wire            n1986;
wire            n19860;
wire            n19861;
wire      [7:0] n19862;
wire            n19863;
wire            n19864;
wire            n19865;
wire            n19866;
wire            n19867;
wire      [7:0] n19868;
wire            n19869;
wire            n1987;
wire            n19870;
wire            n19871;
wire            n19872;
wire            n19873;
wire      [7:0] n19874;
wire            n19875;
wire            n19876;
wire            n19877;
wire            n19878;
wire            n19879;
wire            n1988;
wire      [7:0] n19880;
wire            n19881;
wire            n19882;
wire            n19883;
wire            n19884;
wire            n19885;
wire      [7:0] n19886;
wire            n19887;
wire            n19888;
wire            n19889;
wire            n1989;
wire            n19890;
wire            n19891;
wire      [7:0] n19892;
wire            n19893;
wire            n19894;
wire            n19895;
wire            n19896;
wire            n19897;
wire      [7:0] n19898;
wire            n19899;
wire            n1990;
wire            n19900;
wire            n19901;
wire            n19902;
wire            n19903;
wire      [7:0] n19904;
wire            n19905;
wire            n19906;
wire            n19907;
wire            n19908;
wire            n19909;
wire            n1991;
wire      [7:0] n19910;
wire            n19911;
wire            n19912;
wire            n19913;
wire            n19914;
wire            n19915;
wire      [7:0] n19916;
wire            n19917;
wire            n19918;
wire            n19919;
wire            n1992;
wire            n19920;
wire            n19921;
wire      [7:0] n19922;
wire            n19923;
wire            n19924;
wire            n19925;
wire            n19926;
wire            n19927;
wire      [7:0] n19928;
wire            n19929;
wire            n1993;
wire            n19930;
wire            n19931;
wire            n19932;
wire            n19933;
wire      [7:0] n19934;
wire            n19935;
wire            n19936;
wire            n19937;
wire            n19938;
wire            n19939;
wire            n1994;
wire      [7:0] n19940;
wire            n19941;
wire            n19942;
wire            n19943;
wire            n19944;
wire            n19945;
wire      [7:0] n19946;
wire            n19947;
wire            n19948;
wire            n19949;
wire            n1995;
wire            n19950;
wire            n19951;
wire      [7:0] n19952;
wire            n19953;
wire            n19954;
wire            n19955;
wire            n19956;
wire            n19957;
wire      [7:0] n19958;
wire            n19959;
wire            n1996;
wire            n19960;
wire            n19961;
wire            n19962;
wire            n19963;
wire      [7:0] n19964;
wire            n19965;
wire            n19966;
wire            n19967;
wire            n19968;
wire            n19969;
wire            n1997;
wire      [7:0] n19970;
wire            n19971;
wire            n19972;
wire            n19973;
wire            n19974;
wire            n19975;
wire      [7:0] n19976;
wire            n19977;
wire            n19978;
wire            n19979;
wire            n1998;
wire            n19980;
wire            n19981;
wire      [7:0] n19982;
wire            n19983;
wire            n19984;
wire            n19985;
wire            n19986;
wire            n19987;
wire      [7:0] n19988;
wire            n19989;
wire            n1999;
wire            n19990;
wire            n19991;
wire            n19992;
wire            n19993;
wire      [7:0] n19994;
wire            n19995;
wire            n19996;
wire            n19997;
wire            n19998;
wire            n19999;
wire            n200;
wire            n2000;
wire      [7:0] n20000;
wire            n20001;
wire            n20002;
wire            n20003;
wire            n20004;
wire            n20005;
wire      [7:0] n20006;
wire            n20007;
wire            n20008;
wire            n20009;
wire            n2001;
wire            n20010;
wire            n20011;
wire      [7:0] n20012;
wire            n20013;
wire            n20014;
wire            n20015;
wire            n20016;
wire            n20017;
wire      [7:0] n20018;
wire            n20019;
wire            n2002;
wire            n20020;
wire            n20021;
wire            n20022;
wire            n20023;
wire      [7:0] n20024;
wire            n20025;
wire            n20026;
wire            n20027;
wire            n20028;
wire            n20029;
wire            n2003;
wire      [7:0] n20030;
wire            n20031;
wire            n20032;
wire            n20033;
wire            n20034;
wire            n20035;
wire      [7:0] n20036;
wire            n20037;
wire            n20038;
wire            n20039;
wire            n2004;
wire            n20040;
wire            n20041;
wire      [7:0] n20042;
wire            n20043;
wire            n20044;
wire            n20045;
wire            n20046;
wire            n20047;
wire      [7:0] n20048;
wire            n20049;
wire            n2005;
wire            n20050;
wire            n20051;
wire            n20052;
wire            n20053;
wire      [7:0] n20054;
wire            n20055;
wire            n20056;
wire            n20057;
wire            n20058;
wire            n20059;
wire            n2006;
wire      [7:0] n20060;
wire            n20061;
wire            n20062;
wire            n20063;
wire            n20064;
wire            n20065;
wire      [7:0] n20066;
wire            n20067;
wire            n20068;
wire            n20069;
wire            n2007;
wire            n20070;
wire            n20071;
wire      [7:0] n20072;
wire            n20073;
wire            n20074;
wire            n20075;
wire            n20076;
wire            n20077;
wire      [7:0] n20078;
wire            n20079;
wire            n2008;
wire            n20080;
wire            n20081;
wire            n20082;
wire            n20083;
wire      [7:0] n20084;
wire            n20085;
wire            n20086;
wire            n20087;
wire            n20088;
wire            n20089;
wire            n2009;
wire      [7:0] n20090;
wire            n20091;
wire            n20092;
wire            n20093;
wire            n20094;
wire            n20095;
wire      [7:0] n20096;
wire            n20097;
wire            n20098;
wire            n20099;
wire            n2010;
wire            n20100;
wire            n20101;
wire      [7:0] n20102;
wire            n20103;
wire            n20104;
wire            n20105;
wire            n20106;
wire            n20107;
wire      [7:0] n20108;
wire            n20109;
wire            n2011;
wire            n20110;
wire            n20111;
wire            n20112;
wire            n20113;
wire      [7:0] n20114;
wire            n20115;
wire            n20116;
wire            n20117;
wire            n20118;
wire            n20119;
wire            n2012;
wire      [7:0] n20120;
wire            n20121;
wire            n20122;
wire            n20123;
wire            n20124;
wire            n20125;
wire      [7:0] n20126;
wire            n20127;
wire            n20128;
wire            n20129;
wire            n2013;
wire            n20130;
wire            n20131;
wire      [7:0] n20132;
wire            n20133;
wire            n20134;
wire            n20135;
wire            n20136;
wire            n20137;
wire      [7:0] n20138;
wire            n20139;
wire            n2014;
wire            n20140;
wire            n20141;
wire            n20142;
wire            n20143;
wire      [7:0] n20144;
wire            n20145;
wire            n20146;
wire            n20147;
wire            n20148;
wire            n20149;
wire            n2015;
wire      [7:0] n20150;
wire            n20151;
wire            n20152;
wire            n20153;
wire            n20154;
wire            n20155;
wire      [7:0] n20156;
wire            n20157;
wire            n20158;
wire            n20159;
wire            n2016;
wire            n20160;
wire            n20161;
wire      [7:0] n20162;
wire            n20163;
wire            n20164;
wire            n20165;
wire            n20166;
wire            n20167;
wire      [7:0] n20168;
wire            n20169;
wire            n2017;
wire            n20170;
wire            n20171;
wire            n20172;
wire            n20173;
wire      [7:0] n20174;
wire            n20175;
wire            n20176;
wire            n20177;
wire            n20178;
wire            n20179;
wire            n2018;
wire      [7:0] n20180;
wire            n20181;
wire            n20182;
wire            n20183;
wire            n20184;
wire            n20185;
wire      [7:0] n20186;
wire            n20187;
wire            n20188;
wire            n20189;
wire            n2019;
wire            n20190;
wire            n20191;
wire      [7:0] n20192;
wire            n20193;
wire            n20194;
wire            n20195;
wire            n20196;
wire            n20197;
wire      [7:0] n20198;
wire            n20199;
wire            n202;
wire            n2020;
wire            n20200;
wire            n20201;
wire            n20202;
wire            n20203;
wire      [7:0] n20204;
wire            n20205;
wire            n20206;
wire            n20207;
wire            n20208;
wire            n20209;
wire            n2021;
wire      [7:0] n20210;
wire            n20211;
wire            n20212;
wire            n20213;
wire            n20214;
wire            n20215;
wire      [7:0] n20216;
wire            n20217;
wire            n20218;
wire            n20219;
wire            n2022;
wire            n20220;
wire            n20221;
wire      [7:0] n20222;
wire            n20223;
wire            n20224;
wire            n20225;
wire            n20226;
wire            n20227;
wire      [7:0] n20228;
wire            n20229;
wire            n2023;
wire            n20230;
wire            n20231;
wire            n20232;
wire            n20233;
wire      [7:0] n20234;
wire            n20235;
wire            n20236;
wire            n20237;
wire            n20238;
wire            n20239;
wire            n2024;
wire      [7:0] n20240;
wire            n20241;
wire            n20242;
wire            n20243;
wire            n20244;
wire            n20245;
wire      [7:0] n20246;
wire            n20247;
wire            n20248;
wire            n20249;
wire            n2025;
wire            n20250;
wire            n20251;
wire      [7:0] n20252;
wire            n20253;
wire            n20254;
wire            n20255;
wire            n20256;
wire            n20257;
wire      [7:0] n20258;
wire            n20259;
wire            n2026;
wire            n20260;
wire            n20261;
wire            n20262;
wire            n20263;
wire      [7:0] n20264;
wire            n20265;
wire            n20266;
wire            n20267;
wire            n20268;
wire            n20269;
wire            n2027;
wire      [7:0] n20270;
wire            n20271;
wire            n20272;
wire            n20273;
wire            n20274;
wire            n20275;
wire      [7:0] n20276;
wire            n20277;
wire            n20278;
wire            n20279;
wire            n2028;
wire            n20280;
wire            n20281;
wire      [7:0] n20282;
wire            n20283;
wire            n20284;
wire            n20285;
wire            n20286;
wire            n20287;
wire      [7:0] n20288;
wire            n20289;
wire            n2029;
wire            n20290;
wire            n20291;
wire            n20292;
wire            n20293;
wire      [7:0] n20294;
wire            n20295;
wire            n20296;
wire            n20297;
wire            n20298;
wire            n20299;
wire            n2030;
wire      [7:0] n20300;
wire            n20301;
wire            n20302;
wire            n20303;
wire            n20304;
wire            n20305;
wire      [7:0] n20306;
wire            n20307;
wire            n20308;
wire            n20309;
wire            n2031;
wire            n20310;
wire            n20311;
wire      [7:0] n20312;
wire            n20313;
wire            n20314;
wire            n20315;
wire            n20316;
wire            n20317;
wire      [7:0] n20318;
wire            n20319;
wire            n2032;
wire            n20320;
wire            n20321;
wire            n20322;
wire            n20323;
wire      [7:0] n20324;
wire            n20325;
wire            n20326;
wire            n20327;
wire            n20328;
wire            n20329;
wire            n2033;
wire      [7:0] n20330;
wire            n20331;
wire            n20332;
wire            n20333;
wire            n20334;
wire            n20335;
wire      [7:0] n20336;
wire            n20337;
wire            n20338;
wire            n20339;
wire            n2034;
wire            n20340;
wire            n20341;
wire      [7:0] n20342;
wire            n20343;
wire            n20344;
wire            n20345;
wire            n20346;
wire            n20347;
wire      [7:0] n20348;
wire            n20349;
wire            n2035;
wire            n20350;
wire            n20351;
wire            n20352;
wire            n20353;
wire      [7:0] n20354;
wire            n20355;
wire            n20356;
wire            n20357;
wire            n20358;
wire            n20359;
wire            n2036;
wire      [7:0] n20360;
wire            n20361;
wire            n20362;
wire            n20363;
wire            n20364;
wire            n20365;
wire      [7:0] n20366;
wire            n20367;
wire            n20368;
wire            n20369;
wire            n2037;
wire            n20370;
wire            n20371;
wire      [7:0] n20372;
wire            n20373;
wire            n20374;
wire            n20375;
wire            n20376;
wire            n20377;
wire      [7:0] n20378;
wire            n20379;
wire            n2038;
wire            n20380;
wire            n20381;
wire            n20382;
wire            n20383;
wire      [7:0] n20384;
wire            n20385;
wire            n20386;
wire            n20387;
wire            n20388;
wire            n20389;
wire            n2039;
wire      [7:0] n20390;
wire            n20391;
wire            n20392;
wire            n20393;
wire            n20394;
wire            n20395;
wire      [7:0] n20396;
wire            n20397;
wire            n20398;
wire            n20399;
wire            n204;
wire            n2040;
wire            n20400;
wire            n20401;
wire      [7:0] n20402;
wire            n20403;
wire            n20404;
wire            n20405;
wire            n20406;
wire            n20407;
wire      [7:0] n20408;
wire            n20409;
wire            n2041;
wire            n20410;
wire            n20411;
wire            n20412;
wire            n20413;
wire      [7:0] n20414;
wire            n20415;
wire            n20416;
wire            n20417;
wire            n20418;
wire            n20419;
wire            n2042;
wire      [7:0] n20420;
wire            n20421;
wire            n20422;
wire            n20423;
wire            n20424;
wire            n20425;
wire      [7:0] n20426;
wire            n20427;
wire            n20428;
wire            n20429;
wire            n2043;
wire            n20430;
wire            n20431;
wire      [7:0] n20432;
wire            n20433;
wire            n20434;
wire            n20435;
wire            n20436;
wire            n20437;
wire      [7:0] n20438;
wire            n20439;
wire            n2044;
wire            n20440;
wire            n20441;
wire            n20442;
wire            n20443;
wire      [7:0] n20444;
wire            n20445;
wire            n20446;
wire            n20447;
wire            n20448;
wire            n20449;
wire            n2045;
wire      [7:0] n20450;
wire            n20451;
wire            n20452;
wire            n20453;
wire            n20454;
wire            n20455;
wire      [7:0] n20456;
wire            n20457;
wire            n20458;
wire            n20459;
wire            n2046;
wire            n20460;
wire            n20461;
wire      [7:0] n20462;
wire            n20463;
wire            n20464;
wire            n20465;
wire            n20466;
wire            n20467;
wire      [7:0] n20468;
wire            n20469;
wire            n2047;
wire            n20470;
wire            n20471;
wire            n20472;
wire            n20473;
wire      [7:0] n20474;
wire            n20475;
wire            n20476;
wire            n20477;
wire            n20478;
wire            n20479;
wire            n2048;
wire      [7:0] n20480;
wire            n20481;
wire            n20482;
wire            n20483;
wire            n20484;
wire            n20485;
wire      [7:0] n20486;
wire            n20487;
wire            n20488;
wire            n20489;
wire            n2049;
wire            n20490;
wire            n20491;
wire      [7:0] n20492;
wire            n20493;
wire            n20494;
wire            n20495;
wire            n20496;
wire            n20497;
wire      [7:0] n20498;
wire            n20499;
wire            n2050;
wire            n20500;
wire            n20501;
wire            n20502;
wire            n20503;
wire      [7:0] n20504;
wire            n20505;
wire            n20506;
wire            n20507;
wire            n20508;
wire            n20509;
wire            n2051;
wire      [7:0] n20510;
wire            n20511;
wire            n20512;
wire            n20513;
wire            n20514;
wire            n20515;
wire      [7:0] n20516;
wire            n20517;
wire            n20518;
wire            n20519;
wire            n2052;
wire            n20520;
wire            n20521;
wire      [7:0] n20522;
wire            n20523;
wire            n20524;
wire            n20525;
wire            n20526;
wire            n20527;
wire      [7:0] n20528;
wire            n20529;
wire            n2053;
wire            n20530;
wire            n20531;
wire            n20532;
wire            n20533;
wire      [7:0] n20534;
wire            n20535;
wire            n20536;
wire            n20537;
wire            n20538;
wire            n20539;
wire            n2054;
wire      [7:0] n20540;
wire            n20541;
wire            n20542;
wire            n20543;
wire            n20544;
wire            n20545;
wire      [7:0] n20546;
wire            n20547;
wire            n20548;
wire            n20549;
wire            n2055;
wire            n20550;
wire            n20551;
wire      [7:0] n20552;
wire            n20553;
wire            n20554;
wire            n20555;
wire            n20556;
wire            n20557;
wire      [7:0] n20558;
wire            n20559;
wire            n2056;
wire            n20560;
wire            n20561;
wire            n20562;
wire            n20563;
wire      [7:0] n20564;
wire            n20565;
wire            n20566;
wire            n20567;
wire            n20568;
wire            n20569;
wire            n2057;
wire      [7:0] n20570;
wire            n20571;
wire            n20572;
wire            n20573;
wire            n20574;
wire            n20575;
wire      [7:0] n20576;
wire            n20577;
wire            n20578;
wire            n20579;
wire            n2058;
wire            n20580;
wire            n20581;
wire      [7:0] n20582;
wire            n20583;
wire            n20584;
wire            n20585;
wire            n20586;
wire            n20587;
wire      [7:0] n20588;
wire            n20589;
wire            n2059;
wire            n20590;
wire            n20591;
wire            n20592;
wire            n20593;
wire      [7:0] n20594;
wire            n20595;
wire            n20596;
wire            n20597;
wire            n20598;
wire            n20599;
wire            n206;
wire            n2060;
wire      [7:0] n20600;
wire            n20601;
wire            n20602;
wire            n20603;
wire            n20604;
wire            n20605;
wire      [7:0] n20606;
wire            n20607;
wire            n20608;
wire            n20609;
wire            n2061;
wire            n20610;
wire            n20611;
wire      [7:0] n20612;
wire            n20613;
wire            n20614;
wire            n20615;
wire            n20616;
wire            n20617;
wire      [7:0] n20618;
wire            n20619;
wire            n2062;
wire            n20620;
wire            n20621;
wire            n20622;
wire            n20623;
wire      [7:0] n20624;
wire            n20625;
wire            n20626;
wire            n20627;
wire            n20628;
wire            n20629;
wire            n2063;
wire      [7:0] n20630;
wire            n20631;
wire            n20632;
wire            n20633;
wire            n20634;
wire            n20635;
wire      [7:0] n20636;
wire            n20637;
wire            n20638;
wire            n20639;
wire            n2064;
wire            n20640;
wire            n20641;
wire      [7:0] n20642;
wire            n20643;
wire            n20644;
wire            n20645;
wire            n20646;
wire            n20647;
wire      [7:0] n20648;
wire            n20649;
wire            n2065;
wire            n20650;
wire            n20651;
wire            n20652;
wire            n20653;
wire      [7:0] n20654;
wire            n20655;
wire            n20656;
wire            n20657;
wire            n20658;
wire            n20659;
wire            n2066;
wire      [7:0] n20660;
wire            n20661;
wire            n20662;
wire            n20663;
wire            n20664;
wire            n20665;
wire      [7:0] n20666;
wire            n20667;
wire            n20668;
wire            n20669;
wire            n2067;
wire            n20670;
wire            n20671;
wire      [7:0] n20672;
wire            n20673;
wire            n20674;
wire            n20675;
wire            n20676;
wire            n20677;
wire      [7:0] n20678;
wire            n20679;
wire            n2068;
wire            n20680;
wire            n20681;
wire            n20682;
wire            n20683;
wire      [7:0] n20684;
wire            n20685;
wire            n20686;
wire            n20687;
wire            n20688;
wire            n20689;
wire            n2069;
wire      [7:0] n20690;
wire            n20691;
wire            n20692;
wire            n20693;
wire            n20694;
wire            n20695;
wire      [7:0] n20696;
wire            n20697;
wire            n20698;
wire            n20699;
wire            n2070;
wire            n20700;
wire            n20701;
wire      [7:0] n20702;
wire            n20703;
wire            n20704;
wire            n20705;
wire            n20706;
wire            n20707;
wire      [7:0] n20708;
wire            n20709;
wire            n2071;
wire            n20710;
wire            n20711;
wire            n20712;
wire            n20713;
wire      [7:0] n20714;
wire            n20715;
wire            n20716;
wire            n20717;
wire            n20718;
wire            n20719;
wire            n2072;
wire      [7:0] n20720;
wire            n20721;
wire            n20722;
wire            n20723;
wire            n20724;
wire            n20725;
wire      [7:0] n20726;
wire            n20727;
wire            n20728;
wire            n20729;
wire            n2073;
wire            n20730;
wire            n20731;
wire      [7:0] n20732;
wire            n20733;
wire            n20734;
wire            n20735;
wire            n20736;
wire            n20737;
wire      [7:0] n20738;
wire            n20739;
wire            n2074;
wire            n20740;
wire            n20741;
wire            n20742;
wire            n20743;
wire      [7:0] n20744;
wire            n20745;
wire            n20746;
wire            n20747;
wire            n20748;
wire            n20749;
wire            n2075;
wire      [7:0] n20750;
wire            n20751;
wire            n20752;
wire            n20753;
wire            n20754;
wire            n20755;
wire      [7:0] n20756;
wire            n20757;
wire            n20758;
wire            n20759;
wire            n2076;
wire            n20760;
wire            n20761;
wire      [7:0] n20762;
wire            n20763;
wire            n20764;
wire            n20765;
wire            n20766;
wire            n20767;
wire      [7:0] n20768;
wire            n20769;
wire            n2077;
wire            n20770;
wire            n20771;
wire            n20772;
wire            n20773;
wire      [7:0] n20774;
wire            n20775;
wire            n20776;
wire            n20777;
wire            n20778;
wire            n20779;
wire            n2078;
wire      [7:0] n20780;
wire            n20781;
wire            n20782;
wire            n20783;
wire            n20784;
wire            n20785;
wire      [7:0] n20786;
wire            n20787;
wire            n20788;
wire            n20789;
wire            n2079;
wire            n20790;
wire            n20791;
wire      [7:0] n20792;
wire            n20793;
wire            n20794;
wire            n20795;
wire            n20796;
wire            n20797;
wire      [7:0] n20798;
wire            n20799;
wire            n208;
wire            n2080;
wire            n20800;
wire            n20801;
wire            n20802;
wire            n20803;
wire      [7:0] n20804;
wire            n20805;
wire            n20806;
wire            n20807;
wire            n20808;
wire            n20809;
wire            n2081;
wire      [7:0] n20810;
wire            n20811;
wire            n20812;
wire            n20813;
wire            n20814;
wire            n20815;
wire      [7:0] n20816;
wire            n20817;
wire            n20818;
wire            n20819;
wire            n2082;
wire            n20820;
wire            n20821;
wire      [7:0] n20822;
wire            n20823;
wire            n20824;
wire            n20825;
wire            n20826;
wire            n20827;
wire      [7:0] n20828;
wire            n20829;
wire            n2083;
wire            n20830;
wire            n20831;
wire            n20832;
wire            n20833;
wire      [7:0] n20834;
wire            n20835;
wire            n20836;
wire            n20837;
wire            n20838;
wire            n20839;
wire            n2084;
wire      [7:0] n20840;
wire            n20841;
wire            n20842;
wire            n20843;
wire            n20844;
wire            n20845;
wire      [7:0] n20846;
wire            n20847;
wire            n20848;
wire            n20849;
wire            n2085;
wire            n20850;
wire            n20851;
wire      [7:0] n20852;
wire            n20853;
wire            n20854;
wire            n20855;
wire            n20856;
wire            n20857;
wire      [7:0] n20858;
wire            n20859;
wire            n2086;
wire            n20860;
wire            n20861;
wire            n20862;
wire            n20863;
wire      [7:0] n20864;
wire            n20865;
wire            n20866;
wire            n20867;
wire            n20868;
wire            n20869;
wire            n2087;
wire      [7:0] n20870;
wire            n20871;
wire            n20872;
wire            n20873;
wire            n20874;
wire            n20875;
wire      [7:0] n20876;
wire            n20877;
wire            n20878;
wire            n20879;
wire            n2088;
wire            n20880;
wire            n20881;
wire      [7:0] n20882;
wire            n20883;
wire            n20884;
wire            n20885;
wire            n20886;
wire            n20887;
wire      [7:0] n20888;
wire            n20889;
wire            n2089;
wire            n20890;
wire            n20891;
wire            n20892;
wire            n20893;
wire      [7:0] n20894;
wire            n20895;
wire            n20896;
wire            n20897;
wire            n20898;
wire            n20899;
wire            n2090;
wire      [7:0] n20900;
wire            n20901;
wire            n20902;
wire            n20903;
wire            n20904;
wire            n20905;
wire      [7:0] n20906;
wire            n20907;
wire            n20908;
wire            n20909;
wire            n2091;
wire            n20910;
wire            n20911;
wire      [7:0] n20912;
wire            n20913;
wire            n20914;
wire            n20915;
wire            n20916;
wire            n20917;
wire      [7:0] n20918;
wire            n20919;
wire            n2092;
wire            n20920;
wire            n20921;
wire            n20922;
wire            n20923;
wire      [7:0] n20924;
wire            n20925;
wire            n20926;
wire            n20927;
wire            n20928;
wire            n20929;
wire            n2093;
wire      [7:0] n20930;
wire            n20931;
wire            n20932;
wire            n20933;
wire            n20934;
wire            n20935;
wire      [7:0] n20936;
wire            n20937;
wire            n20938;
wire            n20939;
wire            n2094;
wire            n20940;
wire            n20941;
wire      [7:0] n20942;
wire            n20943;
wire            n20944;
wire            n20945;
wire            n20946;
wire            n20947;
wire      [7:0] n20948;
wire            n20949;
wire            n2095;
wire            n20950;
wire            n20951;
wire            n20952;
wire            n20953;
wire      [7:0] n20954;
wire            n20955;
wire            n20956;
wire            n20957;
wire            n20958;
wire            n20959;
wire            n2096;
wire      [7:0] n20960;
wire            n20961;
wire            n20962;
wire            n20963;
wire            n20964;
wire            n20965;
wire      [7:0] n20966;
wire            n20967;
wire            n20968;
wire            n20969;
wire            n2097;
wire            n20970;
wire            n20971;
wire      [7:0] n20972;
wire            n20973;
wire            n20974;
wire            n20975;
wire            n20976;
wire            n20977;
wire      [7:0] n20978;
wire            n20979;
wire            n2098;
wire            n20980;
wire            n20981;
wire            n20982;
wire            n20983;
wire      [7:0] n20984;
wire            n20985;
wire            n20986;
wire            n20987;
wire            n20988;
wire            n20989;
wire            n2099;
wire      [7:0] n20990;
wire            n20991;
wire            n20992;
wire            n20993;
wire            n20994;
wire            n20995;
wire      [7:0] n20996;
wire            n20997;
wire            n20998;
wire            n20999;
wire            n21;
wire            n210;
wire            n2100;
wire            n21000;
wire            n21001;
wire      [7:0] n21002;
wire            n21003;
wire            n21004;
wire            n21005;
wire            n21006;
wire            n21007;
wire      [7:0] n21008;
wire            n21009;
wire            n2101;
wire            n21010;
wire            n21011;
wire            n21012;
wire            n21013;
wire      [7:0] n21014;
wire            n21015;
wire            n21016;
wire            n21017;
wire            n21018;
wire            n21019;
wire            n2102;
wire      [7:0] n21020;
wire            n21021;
wire            n21022;
wire            n21023;
wire            n21024;
wire            n21025;
wire      [7:0] n21026;
wire            n21027;
wire            n21028;
wire            n21029;
wire            n2103;
wire            n21030;
wire            n21031;
wire      [7:0] n21032;
wire            n21033;
wire            n21034;
wire            n21035;
wire            n21036;
wire            n21037;
wire      [7:0] n21038;
wire            n21039;
wire            n2104;
wire            n21040;
wire            n21041;
wire            n21042;
wire            n21043;
wire      [7:0] n21044;
wire            n21045;
wire            n21046;
wire            n21047;
wire            n21048;
wire            n21049;
wire            n2105;
wire      [7:0] n21050;
wire            n21051;
wire            n21052;
wire            n21053;
wire            n21054;
wire            n21055;
wire      [7:0] n21056;
wire            n21057;
wire            n21058;
wire            n21059;
wire            n2106;
wire            n21060;
wire            n21061;
wire      [7:0] n21062;
wire            n21063;
wire            n21064;
wire            n21065;
wire            n21066;
wire            n21067;
wire      [7:0] n21068;
wire            n21069;
wire            n2107;
wire            n21070;
wire            n21071;
wire            n21072;
wire            n21073;
wire      [7:0] n21074;
wire            n21075;
wire            n21076;
wire            n21077;
wire            n21078;
wire            n21079;
wire            n2108;
wire      [7:0] n21080;
wire            n21081;
wire            n21082;
wire            n21083;
wire            n21084;
wire            n21085;
wire      [7:0] n21086;
wire            n21087;
wire            n21088;
wire            n21089;
wire            n2109;
wire            n21090;
wire            n21091;
wire      [7:0] n21092;
wire            n21093;
wire            n21094;
wire            n21095;
wire            n21096;
wire            n21097;
wire      [7:0] n21098;
wire            n21099;
wire            n2110;
wire            n21100;
wire            n21101;
wire            n21102;
wire            n21103;
wire      [7:0] n21104;
wire            n21105;
wire            n21106;
wire            n21107;
wire            n21108;
wire            n21109;
wire            n2111;
wire      [7:0] n21110;
wire            n21111;
wire            n21112;
wire            n21113;
wire            n21114;
wire            n21115;
wire      [7:0] n21116;
wire            n21117;
wire            n21118;
wire            n21119;
wire            n2112;
wire            n21120;
wire            n21121;
wire      [7:0] n21122;
wire            n21123;
wire            n21124;
wire            n21125;
wire            n21126;
wire            n21127;
wire      [7:0] n21128;
wire            n21129;
wire            n2113;
wire            n21130;
wire            n21131;
wire            n21132;
wire            n21133;
wire      [7:0] n21134;
wire            n21135;
wire            n21136;
wire            n21137;
wire            n21138;
wire            n21139;
wire            n2114;
wire      [7:0] n21140;
wire            n21141;
wire            n21142;
wire            n21143;
wire            n21144;
wire            n21145;
wire      [7:0] n21146;
wire            n21147;
wire            n21148;
wire            n21149;
wire            n2115;
wire            n21150;
wire            n21151;
wire      [7:0] n21152;
wire            n21153;
wire            n21154;
wire            n21155;
wire            n21156;
wire            n21157;
wire      [7:0] n21158;
wire            n21159;
wire            n2116;
wire            n21160;
wire            n21161;
wire            n21162;
wire            n21163;
wire      [7:0] n21164;
wire            n21165;
wire            n21166;
wire            n21167;
wire            n21168;
wire            n21169;
wire            n2117;
wire      [7:0] n21170;
wire            n21171;
wire            n21172;
wire            n21173;
wire            n21174;
wire            n21175;
wire      [7:0] n21176;
wire            n21177;
wire            n21178;
wire            n21179;
wire            n2118;
wire            n21180;
wire            n21181;
wire      [7:0] n21182;
wire            n21183;
wire            n21184;
wire            n21185;
wire            n21186;
wire            n21187;
wire      [7:0] n21188;
wire            n21189;
wire            n2119;
wire            n21190;
wire            n21191;
wire            n21192;
wire            n21193;
wire      [7:0] n21194;
wire            n21195;
wire            n21196;
wire            n21197;
wire            n21198;
wire            n21199;
wire            n212;
wire            n2120;
wire      [7:0] n21200;
wire            n21201;
wire            n21202;
wire            n21203;
wire            n21204;
wire            n21205;
wire      [7:0] n21206;
wire            n21207;
wire            n21208;
wire            n21209;
wire            n2121;
wire            n21210;
wire            n21211;
wire      [7:0] n21212;
wire            n21213;
wire            n21214;
wire            n21215;
wire            n21216;
wire            n21217;
wire      [7:0] n21218;
wire            n21219;
wire            n2122;
wire            n21220;
wire            n21221;
wire            n21222;
wire            n21223;
wire      [7:0] n21224;
wire            n21225;
wire            n21226;
wire            n21227;
wire            n21228;
wire            n21229;
wire            n2123;
wire      [7:0] n21230;
wire            n21231;
wire            n21232;
wire            n21233;
wire            n21234;
wire            n21235;
wire      [7:0] n21236;
wire            n21237;
wire            n21238;
wire            n21239;
wire            n2124;
wire            n21240;
wire            n21241;
wire      [7:0] n21242;
wire            n21243;
wire            n21244;
wire            n21245;
wire            n21246;
wire            n21247;
wire      [7:0] n21248;
wire            n21249;
wire            n2125;
wire            n21250;
wire            n21251;
wire            n21252;
wire            n21253;
wire      [7:0] n21254;
wire            n21255;
wire            n21256;
wire            n21257;
wire            n21258;
wire            n21259;
wire            n2126;
wire      [7:0] n21260;
wire            n21261;
wire            n21262;
wire            n21263;
wire            n21264;
wire            n21265;
wire      [7:0] n21266;
wire            n21267;
wire            n21268;
wire            n21269;
wire            n2127;
wire            n21270;
wire            n21271;
wire      [7:0] n21272;
wire            n21273;
wire            n21274;
wire            n21275;
wire            n21276;
wire            n21277;
wire      [7:0] n21278;
wire            n21279;
wire            n2128;
wire            n21280;
wire            n21281;
wire            n21282;
wire            n21283;
wire      [7:0] n21284;
wire            n21285;
wire            n21286;
wire            n21287;
wire            n21288;
wire            n21289;
wire            n2129;
wire      [7:0] n21290;
wire            n21291;
wire            n21292;
wire            n21293;
wire            n21294;
wire            n21295;
wire      [7:0] n21296;
wire            n21297;
wire            n21298;
wire            n21299;
wire      [7:0] n2130;
wire            n21300;
wire            n21301;
wire      [7:0] n21302;
wire            n21303;
wire            n21304;
wire            n21305;
wire            n21306;
wire            n21307;
wire      [7:0] n21308;
wire            n21309;
wire      [7:0] n2131;
wire            n21310;
wire            n21311;
wire            n21312;
wire            n21313;
wire      [7:0] n21314;
wire            n21315;
wire            n21316;
wire            n21317;
wire            n21318;
wire            n21319;
wire      [7:0] n2132;
wire      [7:0] n21320;
wire            n21321;
wire            n21322;
wire            n21323;
wire            n21324;
wire            n21325;
wire      [7:0] n21326;
wire            n21327;
wire            n21328;
wire            n21329;
wire      [7:0] n2133;
wire            n21330;
wire            n21331;
wire      [7:0] n21332;
wire            n21333;
wire            n21334;
wire            n21335;
wire            n21336;
wire            n21337;
wire      [7:0] n21338;
wire            n21339;
wire      [7:0] n2134;
wire            n21340;
wire            n21341;
wire            n21342;
wire            n21343;
wire      [7:0] n21344;
wire            n21345;
wire            n21346;
wire            n21347;
wire            n21348;
wire            n21349;
wire      [7:0] n2135;
wire      [7:0] n21350;
wire            n21351;
wire            n21352;
wire            n21353;
wire            n21354;
wire            n21355;
wire      [7:0] n21356;
wire            n21357;
wire            n21358;
wire            n21359;
wire      [7:0] n2136;
wire            n21360;
wire            n21361;
wire      [7:0] n21362;
wire            n21363;
wire            n21364;
wire            n21365;
wire            n21366;
wire            n21367;
wire      [7:0] n21368;
wire            n21369;
wire      [7:0] n2137;
wire            n21370;
wire            n21371;
wire            n21372;
wire            n21373;
wire      [7:0] n21374;
wire            n21375;
wire            n21376;
wire            n21377;
wire            n21378;
wire            n21379;
wire      [7:0] n2138;
wire      [7:0] n21380;
wire            n21381;
wire            n21382;
wire            n21383;
wire            n21384;
wire            n21385;
wire      [7:0] n21386;
wire            n21387;
wire            n21388;
wire            n21389;
wire      [7:0] n2139;
wire            n21390;
wire            n21391;
wire      [7:0] n21392;
wire            n21393;
wire            n21394;
wire            n21395;
wire            n21396;
wire            n21397;
wire      [7:0] n21398;
wire            n21399;
wire            n214;
wire      [7:0] n2140;
wire            n21400;
wire            n21401;
wire            n21402;
wire            n21403;
wire      [7:0] n21404;
wire            n21405;
wire            n21406;
wire            n21407;
wire            n21408;
wire            n21409;
wire      [7:0] n2141;
wire      [7:0] n21410;
wire            n21411;
wire            n21412;
wire            n21413;
wire            n21414;
wire            n21415;
wire      [7:0] n21416;
wire            n21417;
wire            n21418;
wire            n21419;
wire      [7:0] n2142;
wire            n21420;
wire            n21421;
wire      [7:0] n21422;
wire            n21423;
wire            n21424;
wire            n21425;
wire            n21426;
wire            n21427;
wire      [7:0] n21428;
wire            n21429;
wire      [7:0] n2143;
wire            n21430;
wire            n21431;
wire            n21432;
wire            n21433;
wire      [7:0] n21434;
wire            n21435;
wire            n21436;
wire            n21437;
wire            n21438;
wire            n21439;
wire      [7:0] n2144;
wire      [7:0] n21440;
wire            n21441;
wire            n21442;
wire            n21443;
wire            n21444;
wire            n21445;
wire      [7:0] n21446;
wire            n21447;
wire            n21448;
wire            n21449;
wire      [7:0] n2145;
wire            n21450;
wire            n21451;
wire      [7:0] n21452;
wire            n21453;
wire            n21454;
wire            n21455;
wire            n21456;
wire            n21457;
wire      [7:0] n21458;
wire            n21459;
wire      [7:0] n2146;
wire            n21460;
wire            n21461;
wire            n21462;
wire            n21463;
wire      [7:0] n21464;
wire            n21465;
wire            n21466;
wire            n21467;
wire            n21468;
wire            n21469;
wire      [7:0] n2147;
wire      [7:0] n21470;
wire            n21471;
wire            n21472;
wire            n21473;
wire            n21474;
wire            n21475;
wire      [7:0] n21476;
wire            n21477;
wire            n21478;
wire            n21479;
wire      [7:0] n2148;
wire            n21480;
wire            n21481;
wire      [7:0] n21482;
wire            n21483;
wire            n21484;
wire            n21485;
wire            n21486;
wire            n21487;
wire      [7:0] n21488;
wire            n21489;
wire      [7:0] n2149;
wire            n21490;
wire            n21491;
wire            n21492;
wire            n21493;
wire      [7:0] n21494;
wire            n21495;
wire            n21496;
wire            n21497;
wire            n21498;
wire            n21499;
wire      [7:0] n2150;
wire      [7:0] n21500;
wire            n21501;
wire            n21502;
wire            n21503;
wire            n21504;
wire            n21505;
wire      [7:0] n21506;
wire            n21507;
wire            n21508;
wire            n21509;
wire      [7:0] n2151;
wire            n21510;
wire            n21511;
wire      [7:0] n21512;
wire            n21513;
wire            n21514;
wire            n21515;
wire            n21516;
wire            n21517;
wire      [7:0] n21518;
wire            n21519;
wire      [7:0] n2152;
wire            n21520;
wire            n21521;
wire            n21522;
wire            n21523;
wire      [7:0] n21524;
wire            n21525;
wire            n21526;
wire            n21527;
wire            n21528;
wire            n21529;
wire      [7:0] n2153;
wire      [7:0] n21530;
wire            n21531;
wire            n21532;
wire            n21533;
wire            n21534;
wire            n21535;
wire      [7:0] n21536;
wire            n21537;
wire            n21538;
wire            n21539;
wire      [7:0] n2154;
wire            n21540;
wire            n21541;
wire      [7:0] n21542;
wire            n21543;
wire            n21544;
wire            n21545;
wire            n21546;
wire            n21547;
wire      [7:0] n21548;
wire            n21549;
wire      [7:0] n2155;
wire            n21550;
wire            n21551;
wire            n21552;
wire            n21553;
wire      [7:0] n21554;
wire            n21555;
wire            n21556;
wire            n21557;
wire            n21558;
wire            n21559;
wire      [7:0] n2156;
wire      [7:0] n21560;
wire            n21561;
wire            n21562;
wire            n21563;
wire            n21564;
wire            n21565;
wire      [7:0] n21566;
wire            n21567;
wire            n21568;
wire            n21569;
wire      [7:0] n2157;
wire            n21570;
wire            n21571;
wire      [7:0] n21572;
wire            n21573;
wire            n21574;
wire            n21575;
wire            n21576;
wire            n21577;
wire      [7:0] n21578;
wire            n21579;
wire      [7:0] n2158;
wire            n21580;
wire            n21581;
wire            n21582;
wire            n21583;
wire      [7:0] n21584;
wire            n21585;
wire            n21586;
wire            n21587;
wire            n21588;
wire            n21589;
wire      [7:0] n2159;
wire      [7:0] n21590;
wire            n21591;
wire            n21592;
wire            n21593;
wire            n21594;
wire            n21595;
wire      [7:0] n21596;
wire            n21597;
wire            n21598;
wire            n21599;
wire            n216;
wire      [7:0] n2160;
wire            n21600;
wire            n21601;
wire      [7:0] n21602;
wire            n21603;
wire            n21604;
wire            n21605;
wire            n21606;
wire            n21607;
wire      [7:0] n21608;
wire            n21609;
wire      [7:0] n2161;
wire            n21610;
wire            n21611;
wire            n21612;
wire            n21613;
wire      [7:0] n21614;
wire            n21615;
wire            n21616;
wire            n21617;
wire            n21618;
wire            n21619;
wire      [7:0] n2162;
wire      [7:0] n21620;
wire            n21621;
wire            n21622;
wire            n21623;
wire            n21624;
wire            n21625;
wire      [7:0] n21626;
wire            n21627;
wire            n21628;
wire            n21629;
wire      [7:0] n2163;
wire            n21630;
wire            n21631;
wire      [7:0] n21632;
wire            n21633;
wire            n21634;
wire            n21635;
wire            n21636;
wire            n21637;
wire      [7:0] n21638;
wire            n21639;
wire      [7:0] n2164;
wire            n21640;
wire            n21641;
wire            n21642;
wire            n21643;
wire      [7:0] n21644;
wire            n21645;
wire            n21646;
wire            n21647;
wire            n21648;
wire            n21649;
wire      [7:0] n2165;
wire      [7:0] n21650;
wire            n21651;
wire            n21652;
wire            n21653;
wire            n21654;
wire            n21655;
wire      [7:0] n21656;
wire            n21657;
wire            n21658;
wire            n21659;
wire      [7:0] n2166;
wire            n21660;
wire            n21661;
wire      [7:0] n21662;
wire            n21663;
wire            n21664;
wire            n21665;
wire            n21666;
wire            n21667;
wire      [7:0] n21668;
wire            n21669;
wire      [7:0] n2167;
wire            n21670;
wire            n21671;
wire            n21672;
wire            n21673;
wire      [7:0] n21674;
wire            n21675;
wire            n21676;
wire            n21677;
wire            n21678;
wire            n21679;
wire      [7:0] n2168;
wire      [7:0] n21680;
wire            n21681;
wire            n21682;
wire            n21683;
wire            n21684;
wire            n21685;
wire      [7:0] n21686;
wire            n21687;
wire            n21688;
wire            n21689;
wire      [7:0] n2169;
wire            n21690;
wire            n21691;
wire      [7:0] n21692;
wire            n21693;
wire            n21694;
wire            n21695;
wire            n21696;
wire            n21697;
wire      [7:0] n21698;
wire            n21699;
wire      [7:0] n2170;
wire            n21700;
wire            n21701;
wire            n21702;
wire            n21703;
wire      [7:0] n21704;
wire            n21705;
wire            n21706;
wire            n21707;
wire            n21708;
wire            n21709;
wire      [7:0] n2171;
wire      [7:0] n21710;
wire            n21711;
wire            n21712;
wire            n21713;
wire            n21714;
wire            n21715;
wire      [7:0] n21716;
wire            n21717;
wire            n21718;
wire            n21719;
wire      [7:0] n2172;
wire            n21720;
wire            n21721;
wire      [7:0] n21722;
wire            n21723;
wire            n21724;
wire            n21725;
wire            n21726;
wire            n21727;
wire      [7:0] n21728;
wire            n21729;
wire      [7:0] n2173;
wire            n21730;
wire            n21731;
wire            n21732;
wire            n21733;
wire      [7:0] n21734;
wire            n21735;
wire            n21736;
wire            n21737;
wire            n21738;
wire            n21739;
wire      [7:0] n2174;
wire      [7:0] n21740;
wire            n21741;
wire            n21742;
wire            n21743;
wire            n21744;
wire            n21745;
wire      [7:0] n21746;
wire            n21747;
wire            n21748;
wire            n21749;
wire      [7:0] n2175;
wire            n21750;
wire            n21751;
wire      [7:0] n21752;
wire            n21753;
wire            n21754;
wire            n21755;
wire            n21756;
wire            n21757;
wire      [7:0] n21758;
wire            n21759;
wire      [7:0] n2176;
wire            n21760;
wire            n21761;
wire            n21762;
wire            n21763;
wire      [7:0] n21764;
wire            n21765;
wire            n21766;
wire            n21767;
wire            n21768;
wire            n21769;
wire      [7:0] n2177;
wire      [7:0] n21770;
wire            n21771;
wire            n21772;
wire            n21773;
wire            n21774;
wire            n21775;
wire      [7:0] n21776;
wire            n21777;
wire            n21778;
wire            n21779;
wire      [7:0] n2178;
wire            n21780;
wire            n21781;
wire      [7:0] n21782;
wire            n21783;
wire            n21784;
wire            n21785;
wire            n21786;
wire            n21787;
wire      [7:0] n21788;
wire            n21789;
wire      [7:0] n2179;
wire            n21790;
wire            n21791;
wire            n21792;
wire            n21793;
wire      [7:0] n21794;
wire            n21795;
wire            n21796;
wire            n21797;
wire            n21798;
wire            n21799;
wire            n218;
wire      [7:0] n2180;
wire      [7:0] n21800;
wire            n21801;
wire            n21802;
wire            n21803;
wire            n21804;
wire            n21805;
wire      [7:0] n21806;
wire            n21807;
wire            n21808;
wire            n21809;
wire      [7:0] n2181;
wire            n21810;
wire            n21811;
wire      [7:0] n21812;
wire            n21813;
wire            n21814;
wire            n21815;
wire            n21816;
wire            n21817;
wire      [7:0] n21818;
wire            n21819;
wire      [7:0] n2182;
wire            n21820;
wire            n21821;
wire            n21822;
wire            n21823;
wire      [7:0] n21824;
wire            n21825;
wire            n21826;
wire            n21827;
wire            n21828;
wire            n21829;
wire      [7:0] n2183;
wire      [7:0] n21830;
wire            n21831;
wire            n21832;
wire            n21833;
wire            n21834;
wire            n21835;
wire      [7:0] n21836;
wire            n21837;
wire            n21838;
wire            n21839;
wire      [7:0] n2184;
wire            n21840;
wire            n21841;
wire      [7:0] n21842;
wire            n21843;
wire            n21844;
wire            n21845;
wire            n21846;
wire            n21847;
wire      [7:0] n21848;
wire            n21849;
wire      [7:0] n2185;
wire            n21850;
wire            n21851;
wire            n21852;
wire            n21853;
wire      [7:0] n21854;
wire            n21855;
wire            n21856;
wire            n21857;
wire            n21858;
wire            n21859;
wire      [7:0] n2186;
wire      [7:0] n21860;
wire            n21861;
wire            n21862;
wire            n21863;
wire            n21864;
wire            n21865;
wire      [7:0] n21866;
wire            n21867;
wire            n21868;
wire            n21869;
wire      [7:0] n2187;
wire            n21870;
wire            n21871;
wire      [7:0] n21872;
wire            n21873;
wire            n21874;
wire            n21875;
wire            n21876;
wire            n21877;
wire      [7:0] n21878;
wire            n21879;
wire      [7:0] n2188;
wire            n21880;
wire            n21881;
wire            n21882;
wire            n21883;
wire      [7:0] n21884;
wire            n21885;
wire            n21886;
wire            n21887;
wire            n21888;
wire            n21889;
wire      [7:0] n2189;
wire      [7:0] n21890;
wire            n21891;
wire            n21892;
wire            n21893;
wire            n21894;
wire            n21895;
wire      [7:0] n21896;
wire            n21897;
wire            n21898;
wire            n21899;
wire      [7:0] n2190;
wire            n21900;
wire            n21901;
wire      [7:0] n21902;
wire            n21903;
wire            n21904;
wire            n21905;
wire            n21906;
wire            n21907;
wire      [7:0] n21908;
wire            n21909;
wire      [7:0] n2191;
wire            n21910;
wire            n21911;
wire            n21912;
wire            n21913;
wire      [7:0] n21914;
wire            n21915;
wire            n21916;
wire            n21917;
wire            n21918;
wire            n21919;
wire      [7:0] n2192;
wire      [7:0] n21920;
wire            n21921;
wire            n21922;
wire            n21923;
wire            n21924;
wire            n21925;
wire      [7:0] n21926;
wire            n21927;
wire            n21928;
wire            n21929;
wire      [7:0] n2193;
wire            n21930;
wire            n21931;
wire      [7:0] n21932;
wire            n21933;
wire            n21934;
wire            n21935;
wire            n21936;
wire            n21937;
wire      [7:0] n21938;
wire            n21939;
wire      [7:0] n2194;
wire            n21940;
wire            n21941;
wire            n21942;
wire            n21943;
wire      [7:0] n21944;
wire            n21945;
wire            n21946;
wire            n21947;
wire            n21948;
wire            n21949;
wire      [7:0] n2195;
wire      [7:0] n21950;
wire            n21951;
wire            n21952;
wire            n21953;
wire            n21954;
wire            n21955;
wire      [7:0] n21956;
wire            n21957;
wire            n21958;
wire            n21959;
wire      [7:0] n2196;
wire            n21960;
wire            n21961;
wire      [7:0] n21962;
wire            n21963;
wire            n21964;
wire            n21965;
wire            n21966;
wire            n21967;
wire      [7:0] n21968;
wire            n21969;
wire      [7:0] n2197;
wire            n21970;
wire            n21971;
wire            n21972;
wire            n21973;
wire      [7:0] n21974;
wire            n21975;
wire            n21976;
wire            n21977;
wire            n21978;
wire            n21979;
wire      [7:0] n2198;
wire      [7:0] n21980;
wire            n21981;
wire            n21982;
wire            n21983;
wire            n21984;
wire            n21985;
wire      [7:0] n21986;
wire            n21987;
wire            n21988;
wire            n21989;
wire      [7:0] n2199;
wire            n21990;
wire            n21991;
wire      [7:0] n21992;
wire            n21993;
wire            n21994;
wire            n21995;
wire            n21996;
wire            n21997;
wire      [7:0] n21998;
wire            n21999;
wire            n220;
wire      [7:0] n2200;
wire            n22000;
wire            n22001;
wire            n22002;
wire            n22003;
wire      [7:0] n22004;
wire            n22005;
wire            n22006;
wire            n22007;
wire            n22008;
wire            n22009;
wire      [7:0] n2201;
wire      [7:0] n22010;
wire            n22011;
wire            n22012;
wire            n22013;
wire            n22014;
wire            n22015;
wire      [7:0] n22016;
wire            n22017;
wire            n22018;
wire            n22019;
wire      [7:0] n2202;
wire            n22020;
wire            n22021;
wire      [7:0] n22022;
wire            n22023;
wire            n22024;
wire            n22025;
wire            n22026;
wire            n22027;
wire      [7:0] n22028;
wire            n22029;
wire      [7:0] n2203;
wire            n22030;
wire            n22031;
wire            n22032;
wire            n22033;
wire      [7:0] n22034;
wire            n22035;
wire            n22036;
wire            n22037;
wire            n22038;
wire            n22039;
wire      [7:0] n2204;
wire      [7:0] n22040;
wire            n22041;
wire            n22042;
wire            n22043;
wire            n22044;
wire            n22045;
wire      [7:0] n22046;
wire            n22047;
wire            n22048;
wire            n22049;
wire      [7:0] n2205;
wire            n22050;
wire            n22051;
wire      [7:0] n22052;
wire            n22053;
wire            n22054;
wire            n22055;
wire            n22056;
wire            n22057;
wire      [7:0] n22058;
wire            n22059;
wire      [7:0] n2206;
wire            n22060;
wire            n22061;
wire            n22062;
wire            n22063;
wire      [7:0] n22064;
wire            n22065;
wire            n22066;
wire            n22067;
wire            n22068;
wire            n22069;
wire      [7:0] n2207;
wire      [7:0] n22070;
wire            n22071;
wire            n22072;
wire            n22073;
wire            n22074;
wire            n22075;
wire      [7:0] n22076;
wire            n22077;
wire            n22078;
wire            n22079;
wire      [7:0] n2208;
wire            n22080;
wire            n22081;
wire      [7:0] n22082;
wire            n22083;
wire            n22084;
wire            n22085;
wire            n22086;
wire            n22087;
wire      [7:0] n22088;
wire            n22089;
wire      [7:0] n2209;
wire            n22090;
wire            n22091;
wire            n22092;
wire            n22093;
wire      [7:0] n22094;
wire            n22095;
wire            n22096;
wire            n22097;
wire            n22098;
wire            n22099;
wire      [7:0] n2210;
wire      [7:0] n22100;
wire            n22101;
wire            n22102;
wire            n22103;
wire            n22104;
wire            n22105;
wire      [7:0] n22106;
wire            n22107;
wire            n22108;
wire            n22109;
wire      [7:0] n2211;
wire            n22110;
wire            n22111;
wire      [7:0] n22112;
wire            n22113;
wire            n22114;
wire            n22115;
wire            n22116;
wire            n22117;
wire      [7:0] n22118;
wire            n22119;
wire      [7:0] n2212;
wire            n22120;
wire            n22121;
wire            n22122;
wire            n22123;
wire      [7:0] n22124;
wire            n22125;
wire            n22126;
wire            n22127;
wire            n22128;
wire            n22129;
wire      [7:0] n2213;
wire      [7:0] n22130;
wire            n22131;
wire            n22132;
wire            n22133;
wire            n22134;
wire            n22135;
wire      [7:0] n22136;
wire            n22137;
wire            n22138;
wire            n22139;
wire      [7:0] n2214;
wire            n22140;
wire            n22141;
wire      [7:0] n22142;
wire            n22143;
wire            n22144;
wire            n22145;
wire            n22146;
wire            n22147;
wire      [7:0] n22148;
wire            n22149;
wire      [7:0] n2215;
wire            n22150;
wire            n22151;
wire            n22152;
wire            n22153;
wire      [7:0] n22154;
wire            n22155;
wire            n22156;
wire            n22157;
wire            n22158;
wire            n22159;
wire      [7:0] n2216;
wire      [7:0] n22160;
wire            n22161;
wire            n22162;
wire            n22163;
wire            n22164;
wire            n22165;
wire      [7:0] n22166;
wire            n22167;
wire            n22168;
wire            n22169;
wire      [7:0] n2217;
wire            n22170;
wire            n22171;
wire      [7:0] n22172;
wire            n22173;
wire            n22174;
wire            n22175;
wire            n22176;
wire            n22177;
wire      [7:0] n22178;
wire            n22179;
wire      [7:0] n2218;
wire            n22180;
wire            n22181;
wire            n22182;
wire            n22183;
wire      [7:0] n22184;
wire            n22185;
wire            n22186;
wire            n22187;
wire            n22188;
wire            n22189;
wire      [7:0] n2219;
wire      [7:0] n22190;
wire            n22191;
wire            n22192;
wire            n22193;
wire            n22194;
wire            n22195;
wire      [7:0] n22196;
wire            n22197;
wire            n22198;
wire            n22199;
wire            n222;
wire      [7:0] n2220;
wire            n22200;
wire            n22201;
wire      [7:0] n22202;
wire            n22203;
wire            n22204;
wire            n22205;
wire            n22206;
wire            n22207;
wire      [7:0] n22208;
wire            n22209;
wire      [7:0] n2221;
wire            n22210;
wire            n22211;
wire            n22212;
wire            n22213;
wire      [7:0] n22214;
wire            n22215;
wire            n22216;
wire            n22217;
wire            n22218;
wire            n22219;
wire      [7:0] n2222;
wire      [7:0] n22220;
wire            n22221;
wire            n22222;
wire            n22223;
wire            n22224;
wire            n22225;
wire      [7:0] n22226;
wire            n22227;
wire            n22228;
wire            n22229;
wire      [7:0] n2223;
wire            n22230;
wire            n22231;
wire      [7:0] n22232;
wire            n22233;
wire            n22234;
wire            n22235;
wire            n22236;
wire            n22237;
wire      [7:0] n22238;
wire            n22239;
wire      [7:0] n2224;
wire            n22240;
wire            n22241;
wire            n22242;
wire            n22243;
wire      [7:0] n22244;
wire            n22245;
wire            n22246;
wire            n22247;
wire            n22248;
wire            n22249;
wire      [7:0] n2225;
wire      [7:0] n22250;
wire            n22251;
wire            n22252;
wire            n22253;
wire            n22254;
wire            n22255;
wire      [7:0] n22256;
wire            n22257;
wire            n22258;
wire            n22259;
wire      [7:0] n2226;
wire            n22260;
wire            n22261;
wire      [7:0] n22262;
wire            n22263;
wire            n22264;
wire            n22265;
wire            n22266;
wire            n22267;
wire      [7:0] n22268;
wire            n22269;
wire      [7:0] n2227;
wire            n22270;
wire            n22271;
wire            n22272;
wire            n22273;
wire      [7:0] n22274;
wire            n22275;
wire            n22276;
wire            n22277;
wire            n22278;
wire            n22279;
wire      [7:0] n2228;
wire      [7:0] n22280;
wire            n22281;
wire            n22282;
wire            n22283;
wire            n22284;
wire            n22285;
wire      [7:0] n22286;
wire            n22287;
wire            n22288;
wire            n22289;
wire      [7:0] n2229;
wire            n22290;
wire            n22291;
wire      [7:0] n22292;
wire            n22293;
wire            n22294;
wire            n22295;
wire            n22296;
wire            n22297;
wire      [7:0] n22298;
wire            n22299;
wire      [7:0] n2230;
wire            n22300;
wire            n22301;
wire            n22302;
wire            n22303;
wire      [7:0] n22304;
wire            n22305;
wire            n22306;
wire            n22307;
wire            n22308;
wire            n22309;
wire      [7:0] n2231;
wire      [7:0] n22310;
wire            n22311;
wire            n22312;
wire            n22313;
wire            n22314;
wire            n22315;
wire      [7:0] n22316;
wire            n22317;
wire            n22318;
wire            n22319;
wire      [7:0] n2232;
wire            n22320;
wire            n22321;
wire      [7:0] n22322;
wire            n22323;
wire            n22324;
wire            n22325;
wire            n22326;
wire            n22327;
wire      [7:0] n22328;
wire            n22329;
wire      [7:0] n2233;
wire            n22330;
wire            n22331;
wire            n22332;
wire            n22333;
wire      [7:0] n22334;
wire            n22335;
wire            n22336;
wire            n22337;
wire            n22338;
wire            n22339;
wire      [7:0] n2234;
wire      [7:0] n22340;
wire            n22341;
wire            n22342;
wire            n22343;
wire            n22344;
wire            n22345;
wire      [7:0] n22346;
wire            n22347;
wire            n22348;
wire            n22349;
wire      [7:0] n2235;
wire            n22350;
wire            n22351;
wire      [7:0] n22352;
wire            n22353;
wire            n22354;
wire            n22355;
wire            n22356;
wire            n22357;
wire      [7:0] n22358;
wire            n22359;
wire      [7:0] n2236;
wire            n22360;
wire            n22361;
wire            n22362;
wire            n22363;
wire      [7:0] n22364;
wire            n22365;
wire            n22366;
wire            n22367;
wire            n22368;
wire            n22369;
wire      [7:0] n2237;
wire      [7:0] n22370;
wire            n22371;
wire            n22372;
wire            n22373;
wire            n22374;
wire            n22375;
wire      [7:0] n22376;
wire            n22377;
wire            n22378;
wire            n22379;
wire      [7:0] n2238;
wire            n22380;
wire            n22381;
wire      [7:0] n22382;
wire            n22383;
wire            n22384;
wire            n22385;
wire            n22386;
wire            n22387;
wire      [7:0] n22388;
wire            n22389;
wire      [7:0] n2239;
wire            n22390;
wire            n22391;
wire            n22392;
wire            n22393;
wire      [7:0] n22394;
wire            n22395;
wire            n22396;
wire            n22397;
wire            n22398;
wire            n22399;
wire            n224;
wire      [7:0] n2240;
wire      [7:0] n22400;
wire            n22401;
wire            n22402;
wire            n22403;
wire            n22404;
wire            n22405;
wire      [7:0] n22406;
wire            n22407;
wire            n22408;
wire            n22409;
wire      [7:0] n2241;
wire            n22410;
wire            n22411;
wire      [7:0] n22412;
wire            n22413;
wire            n22414;
wire            n22415;
wire            n22416;
wire            n22417;
wire      [7:0] n22418;
wire            n22419;
wire      [7:0] n2242;
wire            n22420;
wire            n22421;
wire            n22422;
wire            n22423;
wire      [7:0] n22424;
wire            n22425;
wire            n22426;
wire            n22427;
wire            n22428;
wire            n22429;
wire      [7:0] n2243;
wire      [7:0] n22430;
wire            n22431;
wire            n22432;
wire            n22433;
wire            n22434;
wire            n22435;
wire      [7:0] n22436;
wire            n22437;
wire            n22438;
wire            n22439;
wire      [7:0] n2244;
wire            n22440;
wire            n22441;
wire      [7:0] n22442;
wire            n22443;
wire            n22444;
wire            n22445;
wire            n22446;
wire            n22447;
wire      [7:0] n22448;
wire            n22449;
wire      [7:0] n2245;
wire            n22450;
wire            n22451;
wire            n22452;
wire            n22453;
wire      [7:0] n22454;
wire            n22455;
wire            n22456;
wire            n22457;
wire            n22458;
wire            n22459;
wire      [7:0] n2246;
wire      [7:0] n22460;
wire            n22461;
wire            n22462;
wire            n22463;
wire            n22464;
wire            n22465;
wire      [7:0] n22466;
wire            n22467;
wire            n22468;
wire            n22469;
wire      [7:0] n2247;
wire            n22470;
wire            n22471;
wire      [7:0] n22472;
wire            n22473;
wire            n22474;
wire            n22475;
wire            n22476;
wire            n22477;
wire      [7:0] n22478;
wire            n22479;
wire      [7:0] n2248;
wire            n22480;
wire            n22481;
wire            n22482;
wire            n22483;
wire      [7:0] n22484;
wire            n22485;
wire            n22486;
wire            n22487;
wire            n22488;
wire            n22489;
wire      [7:0] n2249;
wire      [7:0] n22490;
wire            n22491;
wire            n22492;
wire            n22493;
wire            n22494;
wire            n22495;
wire      [7:0] n22496;
wire            n22497;
wire            n22498;
wire            n22499;
wire      [7:0] n2250;
wire            n22500;
wire            n22501;
wire      [7:0] n22502;
wire            n22503;
wire            n22504;
wire            n22505;
wire            n22506;
wire            n22507;
wire      [7:0] n22508;
wire            n22509;
wire      [7:0] n2251;
wire            n22510;
wire            n22511;
wire            n22512;
wire            n22513;
wire      [7:0] n22514;
wire            n22515;
wire            n22516;
wire            n22517;
wire            n22518;
wire            n22519;
wire      [7:0] n2252;
wire      [7:0] n22520;
wire            n22521;
wire            n22522;
wire            n22523;
wire            n22524;
wire            n22525;
wire      [7:0] n22526;
wire            n22527;
wire            n22528;
wire            n22529;
wire      [7:0] n2253;
wire            n22530;
wire            n22531;
wire      [7:0] n22532;
wire            n22533;
wire            n22534;
wire            n22535;
wire            n22536;
wire            n22537;
wire      [7:0] n22538;
wire            n22539;
wire      [7:0] n2254;
wire            n22540;
wire            n22541;
wire            n22542;
wire            n22543;
wire      [7:0] n22544;
wire            n22545;
wire            n22546;
wire            n22547;
wire            n22548;
wire            n22549;
wire      [7:0] n2255;
wire      [7:0] n22550;
wire            n22551;
wire            n22552;
wire            n22553;
wire            n22554;
wire            n22555;
wire      [7:0] n22556;
wire            n22557;
wire            n22558;
wire            n22559;
wire      [7:0] n2256;
wire            n22560;
wire            n22561;
wire      [7:0] n22562;
wire            n22563;
wire            n22564;
wire            n22565;
wire            n22566;
wire            n22567;
wire      [7:0] n22568;
wire            n22569;
wire      [7:0] n2257;
wire            n22570;
wire            n22571;
wire            n22572;
wire            n22573;
wire      [7:0] n22574;
wire            n22575;
wire            n22576;
wire            n22577;
wire            n22578;
wire            n22579;
wire      [7:0] n2258;
wire      [7:0] n22580;
wire            n22581;
wire            n22582;
wire            n22583;
wire            n22584;
wire            n22585;
wire      [7:0] n22586;
wire            n22587;
wire            n22588;
wire            n22589;
wire      [7:0] n2259;
wire            n22590;
wire            n22591;
wire      [7:0] n22592;
wire            n22593;
wire            n22594;
wire            n22595;
wire            n22596;
wire            n22597;
wire      [7:0] n22598;
wire            n22599;
wire            n226;
wire      [7:0] n2260;
wire            n22600;
wire            n22601;
wire            n22602;
wire            n22603;
wire      [7:0] n22604;
wire            n22605;
wire            n22606;
wire            n22607;
wire            n22608;
wire            n22609;
wire      [7:0] n2261;
wire      [7:0] n22610;
wire            n22611;
wire            n22612;
wire            n22613;
wire            n22614;
wire            n22615;
wire      [7:0] n22616;
wire            n22617;
wire            n22618;
wire            n22619;
wire      [7:0] n2262;
wire            n22620;
wire            n22621;
wire      [7:0] n22622;
wire            n22623;
wire            n22624;
wire            n22625;
wire            n22626;
wire            n22627;
wire      [7:0] n22628;
wire            n22629;
wire      [7:0] n2263;
wire            n22630;
wire            n22631;
wire            n22632;
wire            n22633;
wire      [7:0] n22634;
wire            n22635;
wire            n22636;
wire            n22637;
wire            n22638;
wire            n22639;
wire      [7:0] n2264;
wire      [7:0] n22640;
wire            n22641;
wire            n22642;
wire            n22643;
wire            n22644;
wire            n22645;
wire      [7:0] n22646;
wire            n22647;
wire            n22648;
wire            n22649;
wire      [7:0] n2265;
wire            n22650;
wire            n22651;
wire      [7:0] n22652;
wire            n22653;
wire            n22654;
wire            n22655;
wire            n22656;
wire            n22657;
wire      [7:0] n22658;
wire            n22659;
wire      [7:0] n2266;
wire            n22660;
wire            n22661;
wire            n22662;
wire            n22663;
wire      [7:0] n22664;
wire            n22665;
wire            n22666;
wire            n22667;
wire            n22668;
wire            n22669;
wire      [7:0] n2267;
wire      [7:0] n22670;
wire            n22671;
wire            n22672;
wire            n22673;
wire            n22674;
wire            n22675;
wire      [7:0] n22676;
wire            n22677;
wire            n22678;
wire            n22679;
wire      [7:0] n2268;
wire            n22680;
wire            n22681;
wire      [7:0] n22682;
wire            n22683;
wire            n22684;
wire            n22685;
wire            n22686;
wire            n22687;
wire      [7:0] n22688;
wire            n22689;
wire      [7:0] n2269;
wire            n22690;
wire            n22691;
wire            n22692;
wire            n22693;
wire      [7:0] n22694;
wire            n22695;
wire            n22696;
wire            n22697;
wire            n22698;
wire            n22699;
wire      [7:0] n2270;
wire      [7:0] n22700;
wire            n22701;
wire            n22702;
wire            n22703;
wire            n22704;
wire            n22705;
wire      [7:0] n22706;
wire            n22707;
wire            n22708;
wire            n22709;
wire      [7:0] n2271;
wire            n22710;
wire            n22711;
wire      [7:0] n22712;
wire            n22713;
wire            n22714;
wire            n22715;
wire            n22716;
wire            n22717;
wire      [7:0] n22718;
wire            n22719;
wire      [7:0] n2272;
wire            n22720;
wire            n22721;
wire            n22722;
wire            n22723;
wire      [7:0] n22724;
wire            n22725;
wire            n22726;
wire            n22727;
wire            n22728;
wire            n22729;
wire      [7:0] n2273;
wire      [7:0] n22730;
wire            n22731;
wire            n22732;
wire            n22733;
wire            n22734;
wire            n22735;
wire      [7:0] n22736;
wire            n22737;
wire            n22738;
wire            n22739;
wire      [7:0] n2274;
wire            n22740;
wire            n22741;
wire      [7:0] n22742;
wire            n22743;
wire            n22744;
wire            n22745;
wire            n22746;
wire            n22747;
wire      [7:0] n22748;
wire            n22749;
wire      [7:0] n2275;
wire            n22750;
wire            n22751;
wire            n22752;
wire            n22753;
wire      [7:0] n22754;
wire            n22755;
wire            n22756;
wire            n22757;
wire            n22758;
wire            n22759;
wire      [7:0] n2276;
wire      [7:0] n22760;
wire            n22761;
wire            n22762;
wire            n22763;
wire            n22764;
wire            n22765;
wire      [7:0] n22766;
wire            n22767;
wire            n22768;
wire            n22769;
wire      [7:0] n2277;
wire            n22770;
wire            n22771;
wire      [7:0] n22772;
wire            n22773;
wire            n22774;
wire            n22775;
wire            n22776;
wire            n22777;
wire      [7:0] n22778;
wire            n22779;
wire      [7:0] n2278;
wire            n22780;
wire            n22781;
wire            n22782;
wire            n22783;
wire      [7:0] n22784;
wire            n22785;
wire            n22786;
wire            n22787;
wire            n22788;
wire            n22789;
wire      [7:0] n2279;
wire      [7:0] n22790;
wire            n22791;
wire            n22792;
wire            n22793;
wire            n22794;
wire            n22795;
wire      [7:0] n22796;
wire            n22797;
wire            n22798;
wire            n22799;
wire            n228;
wire      [7:0] n2280;
wire            n22800;
wire            n22801;
wire      [7:0] n22802;
wire            n22803;
wire            n22804;
wire            n22805;
wire            n22806;
wire            n22807;
wire      [7:0] n22808;
wire            n22809;
wire      [7:0] n2281;
wire            n22810;
wire            n22811;
wire            n22812;
wire            n22813;
wire      [7:0] n22814;
wire            n22815;
wire            n22816;
wire            n22817;
wire            n22818;
wire            n22819;
wire      [7:0] n2282;
wire      [7:0] n22820;
wire            n22821;
wire            n22822;
wire            n22823;
wire            n22824;
wire            n22825;
wire      [7:0] n22826;
wire            n22827;
wire            n22828;
wire            n22829;
wire      [7:0] n2283;
wire            n22830;
wire            n22831;
wire      [7:0] n22832;
wire            n22833;
wire            n22834;
wire            n22835;
wire            n22836;
wire            n22837;
wire      [7:0] n22838;
wire            n22839;
wire      [7:0] n2284;
wire            n22840;
wire            n22841;
wire            n22842;
wire            n22843;
wire      [7:0] n22844;
wire            n22845;
wire            n22846;
wire            n22847;
wire            n22848;
wire            n22849;
wire      [7:0] n2285;
wire      [7:0] n22850;
wire            n22851;
wire            n22852;
wire            n22853;
wire            n22854;
wire            n22855;
wire      [7:0] n22856;
wire            n22857;
wire            n22858;
wire            n22859;
wire      [7:0] n2286;
wire            n22860;
wire            n22861;
wire      [7:0] n22862;
wire            n22863;
wire            n22864;
wire            n22865;
wire            n22866;
wire            n22867;
wire      [7:0] n22868;
wire            n22869;
wire      [7:0] n2287;
wire            n22870;
wire            n22871;
wire            n22872;
wire            n22873;
wire      [7:0] n22874;
wire            n22875;
wire            n22876;
wire            n22877;
wire            n22878;
wire            n22879;
wire      [7:0] n2288;
wire      [7:0] n22880;
wire            n22881;
wire            n22882;
wire            n22883;
wire            n22884;
wire            n22885;
wire      [7:0] n22886;
wire            n22887;
wire            n22888;
wire            n22889;
wire      [7:0] n2289;
wire            n22890;
wire            n22891;
wire      [7:0] n22892;
wire            n22893;
wire            n22894;
wire            n22895;
wire            n22896;
wire            n22897;
wire      [7:0] n22898;
wire            n22899;
wire      [7:0] n2290;
wire            n22900;
wire            n22901;
wire            n22902;
wire            n22903;
wire      [7:0] n22904;
wire            n22905;
wire            n22906;
wire            n22907;
wire            n22908;
wire            n22909;
wire      [7:0] n2291;
wire      [7:0] n22910;
wire            n22911;
wire            n22912;
wire            n22913;
wire            n22914;
wire            n22915;
wire      [7:0] n22916;
wire            n22917;
wire            n22918;
wire            n22919;
wire      [7:0] n2292;
wire            n22920;
wire            n22921;
wire      [7:0] n22922;
wire            n22923;
wire            n22924;
wire            n22925;
wire            n22926;
wire            n22927;
wire      [7:0] n22928;
wire            n22929;
wire      [7:0] n2293;
wire            n22930;
wire            n22931;
wire            n22932;
wire            n22933;
wire      [7:0] n22934;
wire            n22935;
wire            n22936;
wire            n22937;
wire            n22938;
wire            n22939;
wire      [7:0] n2294;
wire      [7:0] n22940;
wire            n22941;
wire            n22942;
wire            n22943;
wire            n22944;
wire            n22945;
wire      [7:0] n22946;
wire            n22947;
wire            n22948;
wire            n22949;
wire      [7:0] n2295;
wire            n22950;
wire            n22951;
wire      [7:0] n22952;
wire            n22953;
wire            n22954;
wire            n22955;
wire            n22956;
wire            n22957;
wire      [7:0] n22958;
wire            n22959;
wire      [7:0] n2296;
wire            n22960;
wire            n22961;
wire            n22962;
wire            n22963;
wire      [7:0] n22964;
wire            n22965;
wire            n22966;
wire            n22967;
wire            n22968;
wire            n22969;
wire      [7:0] n2297;
wire      [7:0] n22970;
wire            n22971;
wire            n22972;
wire            n22973;
wire            n22974;
wire            n22975;
wire      [7:0] n22976;
wire            n22977;
wire            n22978;
wire            n22979;
wire      [7:0] n2298;
wire            n22980;
wire            n22981;
wire      [7:0] n22982;
wire            n22983;
wire            n22984;
wire            n22985;
wire            n22986;
wire            n22987;
wire      [7:0] n22988;
wire            n22989;
wire      [7:0] n2299;
wire            n22990;
wire            n22991;
wire            n22992;
wire            n22993;
wire      [7:0] n22994;
wire            n22995;
wire            n22996;
wire            n22997;
wire            n22998;
wire            n22999;
wire            n23;
wire            n230;
wire      [7:0] n2300;
wire      [7:0] n23000;
wire            n23001;
wire            n23002;
wire            n23003;
wire            n23004;
wire            n23005;
wire      [7:0] n23006;
wire            n23007;
wire            n23008;
wire            n23009;
wire      [7:0] n2301;
wire            n23010;
wire            n23011;
wire      [7:0] n23012;
wire            n23013;
wire            n23014;
wire            n23015;
wire            n23016;
wire            n23017;
wire      [7:0] n23018;
wire            n23019;
wire      [7:0] n2302;
wire            n23020;
wire            n23021;
wire            n23022;
wire            n23023;
wire      [7:0] n23024;
wire            n23025;
wire            n23026;
wire            n23027;
wire            n23028;
wire            n23029;
wire      [7:0] n2303;
wire      [7:0] n23030;
wire            n23031;
wire            n23032;
wire            n23033;
wire            n23034;
wire            n23035;
wire      [7:0] n23036;
wire            n23037;
wire            n23038;
wire            n23039;
wire      [7:0] n2304;
wire            n23040;
wire            n23041;
wire      [7:0] n23042;
wire            n23043;
wire            n23044;
wire            n23045;
wire            n23046;
wire            n23047;
wire      [7:0] n23048;
wire            n23049;
wire      [7:0] n2305;
wire            n23050;
wire            n23051;
wire            n23052;
wire            n23053;
wire      [7:0] n23054;
wire            n23055;
wire            n23056;
wire            n23057;
wire            n23058;
wire            n23059;
wire      [7:0] n2306;
wire      [7:0] n23060;
wire            n23061;
wire            n23062;
wire            n23063;
wire            n23064;
wire            n23065;
wire      [7:0] n23066;
wire            n23067;
wire            n23068;
wire            n23069;
wire      [7:0] n2307;
wire            n23070;
wire            n23071;
wire      [7:0] n23072;
wire            n23073;
wire            n23074;
wire            n23075;
wire            n23076;
wire            n23077;
wire      [7:0] n23078;
wire            n23079;
wire      [7:0] n2308;
wire            n23080;
wire            n23081;
wire            n23082;
wire            n23083;
wire      [7:0] n23084;
wire            n23085;
wire            n23086;
wire            n23087;
wire            n23088;
wire            n23089;
wire      [7:0] n2309;
wire      [7:0] n23090;
wire            n23091;
wire            n23092;
wire            n23093;
wire            n23094;
wire            n23095;
wire      [7:0] n23096;
wire            n23097;
wire            n23098;
wire            n23099;
wire      [7:0] n2310;
wire            n23100;
wire            n23101;
wire      [7:0] n23102;
wire            n23103;
wire            n23104;
wire            n23105;
wire            n23106;
wire            n23107;
wire      [7:0] n23108;
wire            n23109;
wire      [7:0] n2311;
wire            n23110;
wire            n23111;
wire            n23112;
wire            n23113;
wire      [7:0] n23114;
wire            n23115;
wire            n23116;
wire            n23117;
wire            n23118;
wire            n23119;
wire      [7:0] n2312;
wire      [7:0] n23120;
wire            n23121;
wire            n23122;
wire            n23123;
wire            n23124;
wire            n23125;
wire      [7:0] n23126;
wire            n23127;
wire            n23128;
wire            n23129;
wire      [7:0] n2313;
wire            n23130;
wire            n23131;
wire      [7:0] n23132;
wire            n23133;
wire            n23134;
wire            n23135;
wire            n23136;
wire            n23137;
wire      [7:0] n23138;
wire            n23139;
wire      [7:0] n2314;
wire            n23140;
wire            n23141;
wire            n23142;
wire            n23143;
wire      [7:0] n23144;
wire            n23145;
wire            n23146;
wire            n23147;
wire            n23148;
wire            n23149;
wire      [7:0] n2315;
wire      [7:0] n23150;
wire            n23151;
wire            n23152;
wire            n23153;
wire            n23154;
wire            n23155;
wire      [7:0] n23156;
wire            n23157;
wire            n23158;
wire            n23159;
wire      [7:0] n2316;
wire            n23160;
wire            n23161;
wire      [7:0] n23162;
wire            n23163;
wire            n23164;
wire            n23165;
wire            n23166;
wire            n23167;
wire      [7:0] n23168;
wire            n23169;
wire      [7:0] n2317;
wire            n23170;
wire            n23171;
wire            n23172;
wire            n23173;
wire      [7:0] n23174;
wire            n23175;
wire            n23176;
wire            n23177;
wire            n23178;
wire            n23179;
wire      [7:0] n2318;
wire      [7:0] n23180;
wire            n23181;
wire            n23182;
wire            n23183;
wire            n23184;
wire            n23185;
wire      [7:0] n23186;
wire            n23187;
wire            n23188;
wire            n23189;
wire      [7:0] n2319;
wire            n23190;
wire            n23191;
wire      [7:0] n23192;
wire            n23193;
wire            n23194;
wire            n23195;
wire            n23196;
wire            n23197;
wire      [7:0] n23198;
wire            n23199;
wire            n232;
wire      [7:0] n2320;
wire            n23200;
wire            n23201;
wire            n23202;
wire            n23203;
wire      [7:0] n23204;
wire            n23205;
wire            n23206;
wire            n23207;
wire            n23208;
wire            n23209;
wire      [7:0] n2321;
wire      [7:0] n23210;
wire            n23211;
wire            n23212;
wire            n23213;
wire            n23214;
wire            n23215;
wire      [7:0] n23216;
wire            n23217;
wire            n23218;
wire            n23219;
wire      [7:0] n2322;
wire            n23220;
wire            n23221;
wire      [7:0] n23222;
wire            n23223;
wire            n23224;
wire            n23225;
wire            n23226;
wire            n23227;
wire      [7:0] n23228;
wire            n23229;
wire      [7:0] n2323;
wire            n23230;
wire            n23231;
wire            n23232;
wire            n23233;
wire      [7:0] n23234;
wire            n23235;
wire            n23236;
wire            n23237;
wire            n23238;
wire            n23239;
wire      [7:0] n2324;
wire      [7:0] n23240;
wire            n23241;
wire            n23242;
wire            n23243;
wire            n23244;
wire            n23245;
wire      [7:0] n23246;
wire            n23247;
wire            n23248;
wire            n23249;
wire      [7:0] n2325;
wire            n23250;
wire            n23251;
wire      [7:0] n23252;
wire            n23253;
wire            n23254;
wire            n23255;
wire            n23256;
wire            n23257;
wire      [7:0] n23258;
wire            n23259;
wire      [7:0] n2326;
wire            n23260;
wire            n23261;
wire            n23262;
wire            n23263;
wire      [7:0] n23264;
wire            n23265;
wire            n23266;
wire            n23267;
wire            n23268;
wire            n23269;
wire      [7:0] n2327;
wire      [7:0] n23270;
wire            n23271;
wire            n23272;
wire            n23273;
wire            n23274;
wire            n23275;
wire      [7:0] n23276;
wire            n23277;
wire            n23278;
wire            n23279;
wire      [7:0] n2328;
wire            n23280;
wire            n23281;
wire      [7:0] n23282;
wire            n23283;
wire            n23284;
wire            n23285;
wire            n23286;
wire            n23287;
wire      [7:0] n23288;
wire            n23289;
wire      [7:0] n2329;
wire            n23290;
wire            n23291;
wire            n23292;
wire            n23293;
wire      [7:0] n23294;
wire            n23295;
wire            n23296;
wire            n23297;
wire            n23298;
wire            n23299;
wire      [7:0] n2330;
wire      [7:0] n23300;
wire            n23301;
wire            n23302;
wire            n23303;
wire            n23304;
wire            n23305;
wire      [7:0] n23306;
wire            n23307;
wire            n23308;
wire            n23309;
wire      [7:0] n2331;
wire            n23310;
wire            n23311;
wire      [7:0] n23312;
wire            n23313;
wire            n23314;
wire            n23315;
wire            n23316;
wire            n23317;
wire      [7:0] n23318;
wire            n23319;
wire      [7:0] n2332;
wire            n23320;
wire            n23321;
wire            n23322;
wire            n23323;
wire      [7:0] n23324;
wire            n23325;
wire            n23326;
wire            n23327;
wire            n23328;
wire            n23329;
wire      [7:0] n2333;
wire      [7:0] n23330;
wire            n23331;
wire            n23332;
wire            n23333;
wire            n23334;
wire            n23335;
wire      [7:0] n23336;
wire            n23337;
wire            n23338;
wire            n23339;
wire      [7:0] n2334;
wire            n23340;
wire            n23341;
wire      [7:0] n23342;
wire            n23343;
wire            n23344;
wire            n23345;
wire            n23346;
wire            n23347;
wire      [7:0] n23348;
wire            n23349;
wire      [7:0] n2335;
wire            n23350;
wire            n23351;
wire            n23352;
wire            n23353;
wire      [7:0] n23354;
wire            n23355;
wire            n23356;
wire            n23357;
wire            n23358;
wire            n23359;
wire      [7:0] n2336;
wire      [7:0] n23360;
wire            n23361;
wire            n23362;
wire            n23363;
wire            n23364;
wire            n23365;
wire      [7:0] n23366;
wire            n23367;
wire            n23368;
wire            n23369;
wire      [7:0] n2337;
wire            n23370;
wire            n23371;
wire      [7:0] n23372;
wire            n23373;
wire            n23374;
wire            n23375;
wire            n23376;
wire            n23377;
wire      [7:0] n23378;
wire            n23379;
wire      [7:0] n2338;
wire            n23380;
wire            n23381;
wire            n23382;
wire            n23383;
wire      [7:0] n23384;
wire            n23385;
wire            n23386;
wire            n23387;
wire            n23388;
wire            n23389;
wire      [7:0] n2339;
wire      [7:0] n23390;
wire            n23391;
wire            n23392;
wire            n23393;
wire            n23394;
wire            n23395;
wire      [7:0] n23396;
wire            n23397;
wire            n23398;
wire            n23399;
wire            n234;
wire      [7:0] n2340;
wire            n23400;
wire            n23401;
wire      [7:0] n23402;
wire            n23403;
wire            n23404;
wire            n23405;
wire            n23406;
wire            n23407;
wire      [7:0] n23408;
wire            n23409;
wire      [7:0] n2341;
wire            n23410;
wire            n23411;
wire            n23412;
wire            n23413;
wire      [7:0] n23414;
wire            n23415;
wire            n23416;
wire            n23417;
wire            n23418;
wire            n23419;
wire      [7:0] n2342;
wire      [7:0] n23420;
wire            n23421;
wire            n23422;
wire            n23423;
wire            n23424;
wire            n23425;
wire      [7:0] n23426;
wire            n23427;
wire            n23428;
wire            n23429;
wire      [7:0] n2343;
wire            n23430;
wire            n23431;
wire      [7:0] n23432;
wire            n23433;
wire            n23434;
wire            n23435;
wire            n23436;
wire            n23437;
wire      [7:0] n23438;
wire            n23439;
wire      [7:0] n2344;
wire            n23440;
wire            n23441;
wire            n23442;
wire            n23443;
wire      [7:0] n23444;
wire            n23445;
wire            n23446;
wire            n23447;
wire            n23448;
wire            n23449;
wire      [7:0] n2345;
wire      [7:0] n23450;
wire            n23451;
wire            n23452;
wire            n23453;
wire            n23454;
wire            n23455;
wire      [7:0] n23456;
wire            n23457;
wire            n23458;
wire            n23459;
wire      [7:0] n2346;
wire            n23460;
wire            n23461;
wire      [7:0] n23462;
wire            n23463;
wire            n23464;
wire            n23465;
wire            n23466;
wire            n23467;
wire      [7:0] n23468;
wire            n23469;
wire      [7:0] n2347;
wire            n23470;
wire            n23471;
wire            n23472;
wire            n23473;
wire      [7:0] n23474;
wire            n23475;
wire            n23476;
wire            n23477;
wire            n23478;
wire            n23479;
wire      [7:0] n2348;
wire      [7:0] n23480;
wire            n23481;
wire            n23482;
wire            n23483;
wire            n23484;
wire            n23485;
wire      [7:0] n23486;
wire            n23487;
wire            n23488;
wire            n23489;
wire      [7:0] n2349;
wire            n23490;
wire            n23491;
wire      [7:0] n23492;
wire            n23493;
wire            n23494;
wire            n23495;
wire            n23496;
wire            n23497;
wire      [7:0] n23498;
wire            n23499;
wire      [7:0] n2350;
wire            n23500;
wire            n23501;
wire            n23502;
wire            n23503;
wire      [7:0] n23504;
wire            n23505;
wire            n23506;
wire            n23507;
wire            n23508;
wire            n23509;
wire      [7:0] n2351;
wire      [7:0] n23510;
wire            n23511;
wire            n23512;
wire            n23513;
wire            n23514;
wire            n23515;
wire      [7:0] n23516;
wire            n23517;
wire            n23518;
wire            n23519;
wire      [7:0] n2352;
wire            n23520;
wire            n23521;
wire      [7:0] n23522;
wire            n23523;
wire            n23524;
wire            n23525;
wire            n23526;
wire            n23527;
wire      [7:0] n23528;
wire            n23529;
wire      [7:0] n2353;
wire            n23530;
wire            n23531;
wire            n23532;
wire            n23533;
wire      [7:0] n23534;
wire            n23535;
wire            n23536;
wire            n23537;
wire            n23538;
wire            n23539;
wire      [7:0] n2354;
wire      [7:0] n23540;
wire            n23541;
wire            n23542;
wire            n23543;
wire            n23544;
wire            n23545;
wire      [7:0] n23546;
wire            n23547;
wire            n23548;
wire            n23549;
wire      [7:0] n2355;
wire            n23550;
wire            n23551;
wire      [7:0] n23552;
wire            n23553;
wire            n23554;
wire            n23555;
wire            n23556;
wire            n23557;
wire      [7:0] n23558;
wire            n23559;
wire      [7:0] n2356;
wire            n23560;
wire            n23561;
wire            n23562;
wire            n23563;
wire      [7:0] n23564;
wire            n23565;
wire            n23566;
wire            n23567;
wire            n23568;
wire            n23569;
wire      [7:0] n2357;
wire      [7:0] n23570;
wire            n23571;
wire            n23572;
wire            n23573;
wire            n23574;
wire            n23575;
wire      [7:0] n23576;
wire            n23577;
wire            n23578;
wire            n23579;
wire      [7:0] n2358;
wire            n23580;
wire            n23581;
wire      [7:0] n23582;
wire            n23583;
wire            n23584;
wire            n23585;
wire            n23586;
wire            n23587;
wire      [7:0] n23588;
wire            n23589;
wire      [7:0] n2359;
wire            n23590;
wire            n23591;
wire            n23592;
wire            n23593;
wire      [7:0] n23594;
wire            n23595;
wire            n23596;
wire            n23597;
wire            n23598;
wire            n23599;
wire            n236;
wire      [7:0] n2360;
wire      [7:0] n23600;
wire            n23601;
wire            n23602;
wire            n23603;
wire            n23604;
wire            n23605;
wire      [7:0] n23606;
wire            n23607;
wire            n23608;
wire            n23609;
wire      [7:0] n2361;
wire            n23610;
wire            n23611;
wire      [7:0] n23612;
wire            n23613;
wire            n23614;
wire            n23615;
wire            n23616;
wire            n23617;
wire      [7:0] n23618;
wire            n23619;
wire      [7:0] n2362;
wire            n23620;
wire            n23621;
wire            n23622;
wire            n23623;
wire      [7:0] n23624;
wire            n23625;
wire            n23626;
wire            n23627;
wire            n23628;
wire            n23629;
wire      [7:0] n2363;
wire      [7:0] n23630;
wire            n23631;
wire            n23632;
wire            n23633;
wire            n23634;
wire            n23635;
wire      [7:0] n23636;
wire            n23637;
wire            n23638;
wire            n23639;
wire      [7:0] n2364;
wire            n23640;
wire            n23641;
wire      [7:0] n23642;
wire            n23643;
wire            n23644;
wire            n23645;
wire            n23646;
wire            n23647;
wire      [7:0] n23648;
wire            n23649;
wire      [7:0] n2365;
wire            n23650;
wire            n23651;
wire            n23652;
wire            n23653;
wire      [7:0] n23654;
wire            n23655;
wire            n23656;
wire            n23657;
wire            n23658;
wire            n23659;
wire      [7:0] n2366;
wire      [7:0] n23660;
wire            n23661;
wire            n23662;
wire            n23663;
wire            n23664;
wire            n23665;
wire      [7:0] n23666;
wire            n23667;
wire            n23668;
wire            n23669;
wire      [7:0] n2367;
wire            n23670;
wire            n23671;
wire      [7:0] n23672;
wire            n23673;
wire            n23674;
wire            n23675;
wire            n23676;
wire            n23677;
wire      [7:0] n23678;
wire            n23679;
wire      [7:0] n2368;
wire            n23680;
wire            n23681;
wire            n23682;
wire            n23683;
wire      [7:0] n23684;
wire            n23685;
wire            n23686;
wire            n23687;
wire            n23688;
wire            n23689;
wire      [7:0] n2369;
wire      [7:0] n23690;
wire            n23691;
wire            n23692;
wire            n23693;
wire            n23694;
wire            n23695;
wire      [7:0] n23696;
wire            n23697;
wire            n23698;
wire            n23699;
wire      [7:0] n2370;
wire            n23700;
wire            n23701;
wire      [7:0] n23702;
wire            n23703;
wire            n23704;
wire            n23705;
wire            n23706;
wire            n23707;
wire      [7:0] n23708;
wire            n23709;
wire      [7:0] n2371;
wire            n23710;
wire            n23711;
wire            n23712;
wire            n23713;
wire      [7:0] n23714;
wire            n23715;
wire            n23716;
wire            n23717;
wire            n23718;
wire            n23719;
wire      [7:0] n2372;
wire      [7:0] n23720;
wire            n23721;
wire            n23722;
wire            n23723;
wire            n23724;
wire            n23725;
wire      [7:0] n23726;
wire            n23727;
wire            n23728;
wire            n23729;
wire      [7:0] n2373;
wire            n23730;
wire            n23731;
wire      [7:0] n23732;
wire            n23733;
wire            n23734;
wire            n23735;
wire            n23736;
wire            n23737;
wire      [7:0] n23738;
wire            n23739;
wire      [7:0] n2374;
wire            n23740;
wire            n23741;
wire            n23742;
wire            n23743;
wire      [7:0] n23744;
wire            n23745;
wire            n23746;
wire            n23747;
wire            n23748;
wire            n23749;
wire      [7:0] n2375;
wire      [7:0] n23750;
wire            n23751;
wire            n23752;
wire            n23753;
wire            n23754;
wire            n23755;
wire      [7:0] n23756;
wire            n23757;
wire            n23758;
wire            n23759;
wire      [7:0] n2376;
wire            n23760;
wire            n23761;
wire      [7:0] n23762;
wire            n23763;
wire            n23764;
wire            n23765;
wire            n23766;
wire            n23767;
wire      [7:0] n23768;
wire            n23769;
wire      [7:0] n2377;
wire            n23770;
wire            n23771;
wire            n23772;
wire            n23773;
wire      [7:0] n23774;
wire            n23775;
wire            n23776;
wire            n23777;
wire            n23778;
wire            n23779;
wire      [7:0] n2378;
wire      [7:0] n23780;
wire            n23781;
wire            n23782;
wire            n23783;
wire            n23784;
wire            n23785;
wire      [7:0] n23786;
wire            n23787;
wire            n23788;
wire            n23789;
wire      [7:0] n2379;
wire            n23790;
wire            n23791;
wire      [7:0] n23792;
wire            n23793;
wire            n23794;
wire            n23795;
wire            n23796;
wire            n23797;
wire      [7:0] n23798;
wire            n23799;
wire            n238;
wire      [7:0] n2380;
wire            n23800;
wire            n23801;
wire            n23802;
wire            n23803;
wire      [7:0] n23804;
wire            n23805;
wire            n23806;
wire            n23807;
wire            n23808;
wire            n23809;
wire      [7:0] n2381;
wire      [7:0] n23810;
wire            n23811;
wire            n23812;
wire            n23813;
wire            n23814;
wire            n23815;
wire      [7:0] n23816;
wire            n23817;
wire            n23818;
wire            n23819;
wire      [7:0] n2382;
wire            n23820;
wire            n23821;
wire      [7:0] n23822;
wire            n23823;
wire            n23824;
wire            n23825;
wire            n23826;
wire            n23827;
wire      [7:0] n23828;
wire            n23829;
wire      [7:0] n2383;
wire            n23830;
wire            n23831;
wire            n23832;
wire            n23833;
wire      [7:0] n23834;
wire            n23835;
wire            n23836;
wire            n23837;
wire            n23838;
wire            n23839;
wire      [7:0] n2384;
wire      [7:0] n23840;
wire            n23841;
wire            n23842;
wire            n23843;
wire            n23844;
wire            n23845;
wire      [7:0] n23846;
wire            n23847;
wire            n23848;
wire            n23849;
wire            n2385;
wire            n23850;
wire            n23851;
wire      [7:0] n23852;
wire            n23853;
wire            n23854;
wire            n23855;
wire            n23856;
wire            n23857;
wire      [7:0] n23858;
wire            n23859;
wire            n2386;
wire            n23860;
wire            n23861;
wire            n23862;
wire            n23863;
wire      [7:0] n23864;
wire            n23865;
wire            n23866;
wire            n23867;
wire            n23868;
wire            n23869;
wire      [3:0] n2387;
wire      [7:0] n23870;
wire            n23871;
wire            n23872;
wire            n23873;
wire            n23874;
wire            n23875;
wire      [7:0] n23876;
wire            n23877;
wire            n23878;
wire            n23879;
wire      [4:0] n2388;
wire            n23880;
wire            n23881;
wire      [7:0] n23882;
wire            n23883;
wire            n23884;
wire            n23885;
wire            n23886;
wire            n23887;
wire      [7:0] n23888;
wire            n23889;
wire      [7:0] n2389;
wire            n23890;
wire            n23891;
wire            n23892;
wire            n23893;
wire      [7:0] n23894;
wire            n23895;
wire            n23896;
wire            n23897;
wire            n23898;
wire            n23899;
wire      [3:0] n2390;
wire      [7:0] n23900;
wire            n23901;
wire            n23902;
wire            n23903;
wire            n23904;
wire            n23905;
wire      [7:0] n23906;
wire            n23907;
wire            n23908;
wire            n23909;
wire      [7:0] n2391;
wire            n23910;
wire            n23911;
wire      [7:0] n23912;
wire            n23913;
wire            n23914;
wire            n23915;
wire            n23916;
wire            n23917;
wire      [7:0] n23918;
wire            n23919;
wire      [7:0] n2392;
wire            n23920;
wire            n23921;
wire            n23922;
wire            n23923;
wire      [7:0] n23924;
wire            n23925;
wire            n23926;
wire            n23927;
wire            n23928;
wire            n23929;
wire      [7:0] n2393;
wire      [7:0] n23930;
wire            n23931;
wire            n23932;
wire            n23933;
wire            n23934;
wire            n23935;
wire      [7:0] n23936;
wire            n23937;
wire            n23938;
wire            n23939;
wire            n2394;
wire            n23940;
wire            n23941;
wire      [7:0] n23942;
wire            n23943;
wire            n23944;
wire            n23945;
wire            n23946;
wire            n23947;
wire      [7:0] n23948;
wire            n23949;
wire            n2395;
wire            n23950;
wire            n23951;
wire            n23952;
wire            n23953;
wire      [7:0] n23954;
wire            n23955;
wire            n23956;
wire            n23957;
wire            n23958;
wire            n23959;
wire      [3:0] n2396;
wire      [7:0] n23960;
wire            n23961;
wire            n23962;
wire            n23963;
wire            n23964;
wire            n23965;
wire      [7:0] n23966;
wire            n23967;
wire            n23968;
wire            n23969;
wire      [4:0] n2397;
wire            n23970;
wire            n23971;
wire      [7:0] n23972;
wire            n23973;
wire            n23974;
wire            n23975;
wire            n23976;
wire            n23977;
wire      [7:0] n23978;
wire            n23979;
wire      [7:0] n2398;
wire            n23980;
wire            n23981;
wire            n23982;
wire            n23983;
wire      [7:0] n23984;
wire            n23985;
wire            n23986;
wire            n23987;
wire            n23988;
wire            n23989;
wire      [3:0] n2399;
wire      [7:0] n23990;
wire            n23991;
wire            n23992;
wire            n23993;
wire            n23994;
wire            n23995;
wire      [7:0] n23996;
wire            n23997;
wire            n23998;
wire            n23999;
wire            n240;
wire      [7:0] n2400;
wire            n24000;
wire            n24001;
wire      [7:0] n24002;
wire            n24003;
wire            n24004;
wire            n24005;
wire            n24006;
wire            n24007;
wire      [7:0] n24008;
wire            n24009;
wire      [7:0] n2401;
wire            n24010;
wire            n24011;
wire            n24012;
wire            n24013;
wire      [7:0] n24014;
wire            n24015;
wire            n24016;
wire            n24017;
wire            n24018;
wire            n24019;
wire      [7:0] n2402;
wire      [7:0] n24020;
wire            n24021;
wire            n24022;
wire            n24023;
wire            n24024;
wire            n24025;
wire      [7:0] n24026;
wire            n24027;
wire            n24028;
wire            n24029;
wire            n2403;
wire            n24030;
wire            n24031;
wire      [7:0] n24032;
wire            n24033;
wire            n24034;
wire            n24035;
wire            n24036;
wire            n24037;
wire      [7:0] n24038;
wire            n24039;
wire      [7:0] n2404;
wire            n24040;
wire            n24041;
wire            n24042;
wire            n24043;
wire      [7:0] n24044;
wire            n24045;
wire            n24046;
wire            n24047;
wire            n24048;
wire            n24049;
wire            n2405;
wire      [7:0] n24050;
wire            n24051;
wire            n24052;
wire            n24053;
wire            n24054;
wire            n24055;
wire      [7:0] n24056;
wire            n24057;
wire            n24058;
wire            n24059;
wire            n2406;
wire            n24060;
wire            n24061;
wire      [7:0] n24062;
wire            n24063;
wire            n24064;
wire            n24065;
wire            n24066;
wire            n24067;
wire      [7:0] n24068;
wire            n24069;
wire            n2407;
wire            n24070;
wire            n24071;
wire            n24072;
wire            n24073;
wire      [7:0] n24074;
wire            n24075;
wire            n24076;
wire            n24077;
wire            n24078;
wire            n24079;
wire            n2408;
wire      [7:0] n24080;
wire            n24081;
wire            n24082;
wire            n24083;
wire            n24084;
wire            n24085;
wire      [7:0] n24086;
wire            n24087;
wire            n24088;
wire            n24089;
wire            n2409;
wire            n24090;
wire            n24091;
wire      [7:0] n24092;
wire            n24093;
wire            n24094;
wire            n24095;
wire            n24096;
wire            n24097;
wire      [7:0] n24098;
wire            n24099;
wire            n2410;
wire            n24100;
wire            n24101;
wire            n24102;
wire            n24103;
wire      [7:0] n24104;
wire            n24105;
wire            n24106;
wire            n24107;
wire            n24108;
wire            n24109;
wire            n2411;
wire      [7:0] n24110;
wire            n24111;
wire            n24112;
wire            n24113;
wire            n24114;
wire            n24115;
wire      [7:0] n24116;
wire            n24117;
wire            n24118;
wire            n24119;
wire            n2412;
wire            n24120;
wire            n24121;
wire      [7:0] n24122;
wire            n24123;
wire            n24124;
wire            n24125;
wire            n24126;
wire            n24127;
wire      [7:0] n24128;
wire            n24129;
wire            n2413;
wire            n24130;
wire            n24131;
wire            n24132;
wire            n24133;
wire      [7:0] n24134;
wire            n24135;
wire            n24136;
wire            n24137;
wire            n24138;
wire            n24139;
wire            n2414;
wire      [7:0] n24140;
wire            n24141;
wire            n24142;
wire            n24143;
wire            n24144;
wire            n24145;
wire      [7:0] n24146;
wire            n24147;
wire            n24148;
wire            n24149;
wire            n2415;
wire            n24150;
wire            n24151;
wire      [7:0] n24152;
wire            n24153;
wire            n24154;
wire            n24155;
wire            n24156;
wire            n24157;
wire      [7:0] n24158;
wire            n24159;
wire            n2416;
wire            n24160;
wire            n24161;
wire            n24162;
wire            n24163;
wire      [7:0] n24164;
wire            n24165;
wire            n24166;
wire            n24167;
wire            n24168;
wire            n24169;
wire            n2417;
wire      [7:0] n24170;
wire            n24171;
wire            n24172;
wire            n24173;
wire            n24174;
wire            n24175;
wire      [7:0] n24176;
wire            n24177;
wire            n24178;
wire            n24179;
wire            n2418;
wire            n24180;
wire            n24181;
wire      [7:0] n24182;
wire            n24183;
wire            n24184;
wire            n24185;
wire            n24186;
wire            n24187;
wire      [7:0] n24188;
wire            n24189;
wire            n2419;
wire            n24190;
wire            n24191;
wire            n24192;
wire            n24193;
wire      [7:0] n24194;
wire            n24195;
wire            n24196;
wire            n24197;
wire            n24198;
wire            n24199;
wire            n242;
wire            n2420;
wire      [7:0] n24200;
wire            n24201;
wire            n24202;
wire            n24203;
wire            n24204;
wire            n24205;
wire      [7:0] n24206;
wire            n24207;
wire            n24208;
wire            n24209;
wire            n2421;
wire            n24210;
wire            n24211;
wire      [7:0] n24212;
wire            n24213;
wire            n24214;
wire            n24215;
wire            n24216;
wire            n24217;
wire      [7:0] n24218;
wire            n24219;
wire            n2422;
wire            n24220;
wire            n24221;
wire            n24222;
wire            n24223;
wire      [7:0] n24224;
wire            n24225;
wire            n24226;
wire            n24227;
wire            n24228;
wire            n24229;
wire            n2423;
wire      [7:0] n24230;
wire            n24231;
wire            n24232;
wire            n24233;
wire            n24234;
wire            n24235;
wire      [7:0] n24236;
wire            n24237;
wire            n24238;
wire            n24239;
wire            n2424;
wire            n24240;
wire            n24241;
wire      [7:0] n24242;
wire            n24243;
wire            n24244;
wire            n24245;
wire            n24246;
wire            n24247;
wire      [7:0] n24248;
wire            n24249;
wire            n2425;
wire            n24250;
wire            n24251;
wire            n24252;
wire            n24253;
wire      [7:0] n24254;
wire            n24255;
wire            n24256;
wire            n24257;
wire            n24258;
wire            n24259;
wire            n2426;
wire      [7:0] n24260;
wire            n24261;
wire            n24262;
wire            n24263;
wire            n24264;
wire            n24265;
wire      [7:0] n24266;
wire            n24267;
wire            n24268;
wire            n24269;
wire            n2427;
wire            n24270;
wire            n24271;
wire      [7:0] n24272;
wire            n24273;
wire            n24274;
wire            n24275;
wire            n24276;
wire            n24277;
wire      [7:0] n24278;
wire            n24279;
wire            n2428;
wire            n24280;
wire            n24281;
wire            n24282;
wire            n24283;
wire      [7:0] n24284;
wire            n24285;
wire            n24286;
wire            n24287;
wire            n24288;
wire            n24289;
wire            n2429;
wire      [7:0] n24290;
wire            n24291;
wire            n24292;
wire            n24293;
wire            n24294;
wire            n24295;
wire      [7:0] n24296;
wire            n24297;
wire            n24298;
wire            n24299;
wire            n2430;
wire            n24300;
wire            n24301;
wire      [7:0] n24302;
wire            n24303;
wire            n24304;
wire            n24305;
wire            n24306;
wire            n24307;
wire      [7:0] n24308;
wire            n24309;
wire            n2431;
wire            n24310;
wire            n24311;
wire            n24312;
wire            n24313;
wire      [7:0] n24314;
wire            n24315;
wire            n24316;
wire            n24317;
wire            n24318;
wire            n24319;
wire            n2432;
wire      [7:0] n24320;
wire            n24321;
wire            n24322;
wire            n24323;
wire            n24324;
wire            n24325;
wire      [7:0] n24326;
wire            n24327;
wire            n24328;
wire            n24329;
wire            n2433;
wire            n24330;
wire            n24331;
wire      [7:0] n24332;
wire            n24333;
wire            n24334;
wire            n24335;
wire            n24336;
wire            n24337;
wire      [7:0] n24338;
wire            n24339;
wire            n2434;
wire            n24340;
wire            n24341;
wire            n24342;
wire            n24343;
wire      [7:0] n24344;
wire            n24345;
wire            n24346;
wire            n24347;
wire            n24348;
wire            n24349;
wire            n2435;
wire      [7:0] n24350;
wire            n24351;
wire            n24352;
wire            n24353;
wire            n24354;
wire            n24355;
wire      [7:0] n24356;
wire            n24357;
wire            n24358;
wire            n24359;
wire            n2436;
wire            n24360;
wire            n24361;
wire      [7:0] n24362;
wire            n24363;
wire            n24364;
wire            n24365;
wire            n24366;
wire            n24367;
wire      [7:0] n24368;
wire            n24369;
wire            n2437;
wire            n24370;
wire            n24371;
wire            n24372;
wire            n24373;
wire      [7:0] n24374;
wire            n24375;
wire            n24376;
wire            n24377;
wire            n24378;
wire            n24379;
wire            n2438;
wire      [7:0] n24380;
wire            n24381;
wire            n24382;
wire            n24383;
wire            n24384;
wire            n24385;
wire      [7:0] n24386;
wire            n24387;
wire            n24388;
wire            n24389;
wire            n2439;
wire            n24390;
wire            n24391;
wire      [7:0] n24392;
wire            n24393;
wire            n24394;
wire            n24395;
wire            n24396;
wire            n24397;
wire      [7:0] n24398;
wire            n24399;
wire            n244;
wire            n2440;
wire            n24400;
wire            n24401;
wire            n24402;
wire            n24403;
wire      [7:0] n24404;
wire            n24405;
wire            n24406;
wire            n24407;
wire            n24408;
wire            n24409;
wire            n2441;
wire      [7:0] n24410;
wire            n24411;
wire            n24412;
wire            n24413;
wire            n24414;
wire            n24415;
wire      [7:0] n24416;
wire            n24417;
wire            n24418;
wire            n24419;
wire            n2442;
wire            n24420;
wire            n24421;
wire      [7:0] n24422;
wire            n24423;
wire            n24424;
wire            n24425;
wire            n24426;
wire            n24427;
wire      [7:0] n24428;
wire            n24429;
wire            n2443;
wire            n24430;
wire            n24431;
wire            n24432;
wire            n24433;
wire      [7:0] n24434;
wire            n24435;
wire            n24436;
wire            n24437;
wire            n24438;
wire            n24439;
wire            n2444;
wire      [7:0] n24440;
wire            n24441;
wire            n24442;
wire            n24443;
wire            n24444;
wire            n24445;
wire      [7:0] n24446;
wire            n24447;
wire            n24448;
wire            n24449;
wire            n2445;
wire            n24450;
wire            n24451;
wire      [7:0] n24452;
wire            n24453;
wire            n24454;
wire            n24455;
wire            n24456;
wire            n24457;
wire      [7:0] n24458;
wire            n24459;
wire            n2446;
wire            n24460;
wire            n24461;
wire            n24462;
wire            n24463;
wire      [7:0] n24464;
wire            n24465;
wire            n24466;
wire            n24467;
wire            n24468;
wire            n24469;
wire            n2447;
wire      [7:0] n24470;
wire            n24471;
wire            n24472;
wire            n24473;
wire            n24474;
wire            n24475;
wire      [7:0] n24476;
wire            n24477;
wire            n24478;
wire            n24479;
wire            n2448;
wire            n24480;
wire            n24481;
wire      [7:0] n24482;
wire            n24483;
wire            n24484;
wire            n24485;
wire            n24486;
wire            n24487;
wire      [7:0] n24488;
wire            n24489;
wire            n2449;
wire            n24490;
wire            n24491;
wire            n24492;
wire            n24493;
wire      [7:0] n24494;
wire            n24495;
wire            n24496;
wire            n24497;
wire            n24498;
wire            n24499;
wire            n2450;
wire      [7:0] n24500;
wire            n24501;
wire            n24502;
wire            n24503;
wire            n24504;
wire            n24505;
wire      [7:0] n24506;
wire            n24507;
wire            n24508;
wire            n24509;
wire            n2451;
wire            n24510;
wire            n24511;
wire      [7:0] n24512;
wire            n24513;
wire            n24514;
wire            n24515;
wire            n24516;
wire            n24517;
wire      [7:0] n24518;
wire            n24519;
wire            n2452;
wire            n24520;
wire            n24521;
wire            n24522;
wire            n24523;
wire      [7:0] n24524;
wire            n24525;
wire            n24526;
wire            n24527;
wire            n24528;
wire            n24529;
wire            n2453;
wire      [7:0] n24530;
wire            n24531;
wire            n24532;
wire            n24533;
wire            n24534;
wire            n24535;
wire      [7:0] n24536;
wire            n24537;
wire            n24538;
wire            n24539;
wire            n2454;
wire            n24540;
wire            n24541;
wire      [7:0] n24542;
wire            n24543;
wire            n24544;
wire            n24545;
wire            n24546;
wire            n24547;
wire      [7:0] n24548;
wire            n24549;
wire            n2455;
wire            n24550;
wire            n24551;
wire            n24552;
wire            n24553;
wire      [7:0] n24554;
wire            n24555;
wire            n24556;
wire            n24557;
wire            n24558;
wire            n24559;
wire            n2456;
wire      [7:0] n24560;
wire            n24561;
wire            n24562;
wire            n24563;
wire            n24564;
wire            n24565;
wire      [7:0] n24566;
wire            n24567;
wire            n24568;
wire            n24569;
wire            n2457;
wire            n24570;
wire            n24571;
wire      [7:0] n24572;
wire            n24573;
wire            n24574;
wire            n24575;
wire            n24576;
wire            n24577;
wire      [7:0] n24578;
wire            n24579;
wire            n2458;
wire            n24580;
wire            n24581;
wire            n24582;
wire            n24583;
wire      [7:0] n24584;
wire            n24585;
wire            n24586;
wire            n24587;
wire            n24588;
wire            n24589;
wire            n2459;
wire      [7:0] n24590;
wire            n24591;
wire            n24592;
wire            n24593;
wire            n24594;
wire            n24595;
wire      [7:0] n24596;
wire            n24597;
wire            n24598;
wire            n24599;
wire            n246;
wire            n2460;
wire            n24600;
wire            n24601;
wire      [7:0] n24602;
wire            n24603;
wire            n24604;
wire            n24605;
wire            n24606;
wire            n24607;
wire      [7:0] n24608;
wire            n24609;
wire            n2461;
wire            n24610;
wire            n24611;
wire            n24612;
wire            n24613;
wire      [7:0] n24614;
wire            n24615;
wire            n24616;
wire            n24617;
wire            n24618;
wire            n24619;
wire            n2462;
wire      [7:0] n24620;
wire            n24621;
wire            n24622;
wire            n24623;
wire            n24624;
wire            n24625;
wire      [7:0] n24626;
wire            n24627;
wire            n24628;
wire            n24629;
wire            n2463;
wire            n24630;
wire            n24631;
wire      [7:0] n24632;
wire            n24633;
wire            n24634;
wire            n24635;
wire            n24636;
wire            n24637;
wire      [7:0] n24638;
wire            n24639;
wire            n2464;
wire            n24640;
wire            n24641;
wire            n24642;
wire            n24643;
wire      [7:0] n24644;
wire            n24645;
wire            n24646;
wire            n24647;
wire            n24648;
wire            n24649;
wire            n2465;
wire      [7:0] n24650;
wire            n24651;
wire            n24652;
wire            n24653;
wire            n24654;
wire            n24655;
wire      [7:0] n24656;
wire            n24657;
wire            n24658;
wire            n24659;
wire            n2466;
wire            n24660;
wire            n24661;
wire      [7:0] n24662;
wire            n24663;
wire            n24664;
wire            n24665;
wire            n24666;
wire            n24667;
wire      [7:0] n24668;
wire            n24669;
wire            n2467;
wire            n24670;
wire            n24671;
wire            n24672;
wire            n24673;
wire      [7:0] n24674;
wire            n24675;
wire            n24676;
wire            n24677;
wire            n24678;
wire            n24679;
wire            n2468;
wire      [7:0] n24680;
wire            n24681;
wire            n24682;
wire            n24683;
wire            n24684;
wire            n24685;
wire      [7:0] n24686;
wire            n24687;
wire            n24688;
wire            n24689;
wire            n2469;
wire            n24690;
wire            n24691;
wire      [7:0] n24692;
wire            n24693;
wire            n24694;
wire            n24695;
wire            n24696;
wire            n24697;
wire      [7:0] n24698;
wire            n24699;
wire            n2470;
wire            n24700;
wire            n24701;
wire            n24702;
wire            n24703;
wire      [7:0] n24704;
wire            n24705;
wire            n24706;
wire            n24707;
wire            n24708;
wire            n24709;
wire            n2471;
wire      [7:0] n24710;
wire            n24711;
wire            n24712;
wire            n24713;
wire            n24714;
wire            n24715;
wire      [7:0] n24716;
wire            n24717;
wire            n24718;
wire            n24719;
wire            n2472;
wire            n24720;
wire            n24721;
wire      [7:0] n24722;
wire            n24723;
wire            n24724;
wire            n24725;
wire            n24726;
wire            n24727;
wire      [7:0] n24728;
wire            n24729;
wire            n2473;
wire            n24730;
wire            n24731;
wire            n24732;
wire            n24733;
wire      [7:0] n24734;
wire            n24735;
wire            n24736;
wire            n24737;
wire            n24738;
wire            n24739;
wire            n2474;
wire      [7:0] n24740;
wire            n24741;
wire            n24742;
wire            n24743;
wire            n24744;
wire            n24745;
wire      [7:0] n24746;
wire            n24747;
wire            n24748;
wire            n24749;
wire            n2475;
wire            n24750;
wire            n24751;
wire      [7:0] n24752;
wire            n24753;
wire            n24754;
wire            n24755;
wire            n24756;
wire            n24757;
wire      [7:0] n24758;
wire            n24759;
wire            n2476;
wire            n24760;
wire            n24761;
wire            n24762;
wire            n24763;
wire      [7:0] n24764;
wire            n24765;
wire            n24766;
wire            n24767;
wire            n24768;
wire            n24769;
wire            n2477;
wire      [7:0] n24770;
wire            n24771;
wire            n24772;
wire            n24773;
wire            n24774;
wire            n24775;
wire      [7:0] n24776;
wire            n24777;
wire            n24778;
wire            n24779;
wire            n2478;
wire            n24780;
wire            n24781;
wire      [7:0] n24782;
wire            n24783;
wire            n24784;
wire            n24785;
wire            n24786;
wire            n24787;
wire      [7:0] n24788;
wire            n24789;
wire            n2479;
wire            n24790;
wire            n24791;
wire            n24792;
wire            n24793;
wire      [7:0] n24794;
wire            n24795;
wire            n24796;
wire            n24797;
wire            n24798;
wire            n24799;
wire            n248;
wire            n2480;
wire      [7:0] n24800;
wire            n24801;
wire            n24802;
wire            n24803;
wire            n24804;
wire            n24805;
wire      [7:0] n24806;
wire            n24807;
wire            n24808;
wire            n24809;
wire            n2481;
wire            n24810;
wire            n24811;
wire      [7:0] n24812;
wire            n24813;
wire            n24814;
wire            n24815;
wire            n24816;
wire            n24817;
wire      [7:0] n24818;
wire            n24819;
wire            n2482;
wire            n24820;
wire            n24821;
wire            n24822;
wire            n24823;
wire      [7:0] n24824;
wire            n24825;
wire            n24826;
wire            n24827;
wire            n24828;
wire            n24829;
wire            n2483;
wire      [7:0] n24830;
wire            n24831;
wire            n24832;
wire            n24833;
wire            n24834;
wire            n24835;
wire      [7:0] n24836;
wire            n24837;
wire            n24838;
wire            n24839;
wire            n2484;
wire            n24840;
wire            n24841;
wire      [7:0] n24842;
wire            n24843;
wire            n24844;
wire            n24845;
wire            n24846;
wire            n24847;
wire      [7:0] n24848;
wire            n24849;
wire            n2485;
wire            n24850;
wire            n24851;
wire            n24852;
wire            n24853;
wire      [7:0] n24854;
wire            n24855;
wire            n24856;
wire            n24857;
wire            n24858;
wire            n24859;
wire            n2486;
wire      [7:0] n24860;
wire            n24861;
wire            n24862;
wire            n24863;
wire            n24864;
wire            n24865;
wire      [7:0] n24866;
wire            n24867;
wire            n24868;
wire            n24869;
wire            n2487;
wire            n24870;
wire            n24871;
wire      [7:0] n24872;
wire            n24873;
wire            n24874;
wire            n24875;
wire            n24876;
wire            n24877;
wire      [7:0] n24878;
wire            n24879;
wire            n2488;
wire            n24880;
wire            n24881;
wire            n24882;
wire            n24883;
wire      [7:0] n24884;
wire            n24885;
wire            n24886;
wire            n24887;
wire            n24888;
wire            n24889;
wire            n2489;
wire      [7:0] n24890;
wire            n24891;
wire            n24892;
wire            n24893;
wire            n24894;
wire            n24895;
wire      [7:0] n24896;
wire            n24897;
wire            n24898;
wire            n24899;
wire            n2490;
wire            n24900;
wire            n24901;
wire      [7:0] n24902;
wire            n24903;
wire            n24904;
wire            n24905;
wire            n24906;
wire            n24907;
wire      [7:0] n24908;
wire            n24909;
wire            n2491;
wire            n24910;
wire            n24911;
wire            n24912;
wire            n24913;
wire      [7:0] n24914;
wire            n24915;
wire            n24916;
wire            n24917;
wire            n24918;
wire            n24919;
wire            n2492;
wire      [7:0] n24920;
wire            n24921;
wire            n24922;
wire            n24923;
wire            n24924;
wire            n24925;
wire      [7:0] n24926;
wire            n24927;
wire            n24928;
wire            n24929;
wire            n2493;
wire            n24930;
wire            n24931;
wire      [7:0] n24932;
wire            n24933;
wire            n24934;
wire            n24935;
wire            n24936;
wire            n24937;
wire      [7:0] n24938;
wire            n24939;
wire            n2494;
wire            n24940;
wire            n24941;
wire            n24942;
wire            n24943;
wire      [7:0] n24944;
wire            n24945;
wire            n24946;
wire            n24947;
wire            n24948;
wire            n24949;
wire            n2495;
wire      [7:0] n24950;
wire            n24951;
wire            n24952;
wire            n24953;
wire            n24954;
wire            n24955;
wire      [7:0] n24956;
wire            n24957;
wire            n24958;
wire            n24959;
wire            n2496;
wire            n24960;
wire            n24961;
wire      [7:0] n24962;
wire            n24963;
wire            n24964;
wire            n24965;
wire            n24966;
wire            n24967;
wire      [7:0] n24968;
wire            n24969;
wire            n2497;
wire            n24970;
wire            n24971;
wire            n24972;
wire            n24973;
wire      [7:0] n24974;
wire            n24975;
wire            n24976;
wire            n24977;
wire            n24978;
wire            n24979;
wire            n2498;
wire      [7:0] n24980;
wire            n24981;
wire            n24982;
wire            n24983;
wire            n24984;
wire            n24985;
wire      [7:0] n24986;
wire            n24987;
wire            n24988;
wire            n24989;
wire            n2499;
wire            n24990;
wire            n24991;
wire      [7:0] n24992;
wire            n24993;
wire            n24994;
wire            n24995;
wire            n24996;
wire            n24997;
wire      [7:0] n24998;
wire            n24999;
wire            n25;
wire            n250;
wire            n2500;
wire            n25000;
wire            n25001;
wire            n25002;
wire            n25003;
wire      [7:0] n25004;
wire            n25005;
wire            n25006;
wire            n25007;
wire            n25008;
wire            n25009;
wire            n2501;
wire      [7:0] n25010;
wire            n25011;
wire            n25012;
wire            n25013;
wire            n25014;
wire            n25015;
wire      [7:0] n25016;
wire            n25017;
wire            n25018;
wire            n25019;
wire            n2502;
wire            n25020;
wire            n25021;
wire      [7:0] n25022;
wire            n25023;
wire            n25024;
wire            n25025;
wire            n25026;
wire            n25027;
wire      [7:0] n25028;
wire            n25029;
wire            n2503;
wire            n25030;
wire            n25031;
wire            n25032;
wire            n25033;
wire      [7:0] n25034;
wire            n25035;
wire            n25036;
wire            n25037;
wire            n25038;
wire            n25039;
wire            n2504;
wire      [7:0] n25040;
wire            n25041;
wire            n25042;
wire            n25043;
wire            n25044;
wire            n25045;
wire      [7:0] n25046;
wire            n25047;
wire            n25048;
wire            n25049;
wire            n2505;
wire            n25050;
wire            n25051;
wire      [7:0] n25052;
wire            n25053;
wire            n25054;
wire            n25055;
wire            n25056;
wire            n25057;
wire      [7:0] n25058;
wire            n25059;
wire            n2506;
wire            n25060;
wire            n25061;
wire            n25062;
wire            n25063;
wire      [7:0] n25064;
wire            n25065;
wire            n25066;
wire            n25067;
wire            n25068;
wire            n25069;
wire            n2507;
wire      [7:0] n25070;
wire            n25071;
wire            n25072;
wire            n25073;
wire            n25074;
wire            n25075;
wire      [7:0] n25076;
wire            n25077;
wire            n25078;
wire            n25079;
wire            n2508;
wire            n25080;
wire            n25081;
wire      [7:0] n25082;
wire            n25083;
wire            n25084;
wire            n25085;
wire            n25086;
wire            n25087;
wire      [7:0] n25088;
wire            n25089;
wire            n2509;
wire            n25090;
wire            n25091;
wire            n25092;
wire            n25093;
wire      [7:0] n25094;
wire            n25095;
wire            n25096;
wire            n25097;
wire            n25098;
wire            n25099;
wire            n2510;
wire      [7:0] n25100;
wire            n25101;
wire            n25102;
wire            n25103;
wire            n25104;
wire            n25105;
wire      [7:0] n25106;
wire            n25107;
wire            n25108;
wire            n25109;
wire            n2511;
wire            n25110;
wire            n25111;
wire      [7:0] n25112;
wire            n25113;
wire            n25114;
wire            n25115;
wire            n25116;
wire            n25117;
wire      [7:0] n25118;
wire            n25119;
wire            n2512;
wire            n25120;
wire            n25121;
wire            n25122;
wire            n25123;
wire      [7:0] n25124;
wire            n25125;
wire            n25126;
wire            n25127;
wire            n25128;
wire            n25129;
wire            n2513;
wire      [7:0] n25130;
wire            n25131;
wire            n25132;
wire            n25133;
wire            n25134;
wire            n25135;
wire      [7:0] n25136;
wire            n25137;
wire            n25138;
wire            n25139;
wire            n2514;
wire            n25140;
wire            n25141;
wire      [7:0] n25142;
wire            n25143;
wire            n25144;
wire            n25145;
wire            n25146;
wire            n25147;
wire      [7:0] n25148;
wire            n25149;
wire            n2515;
wire            n25150;
wire            n25151;
wire            n25152;
wire            n25153;
wire      [7:0] n25154;
wire            n25155;
wire            n25156;
wire            n25157;
wire            n25158;
wire            n25159;
wire            n2516;
wire      [7:0] n25160;
wire            n25161;
wire            n25162;
wire            n25163;
wire            n25164;
wire            n25165;
wire      [7:0] n25166;
wire            n25167;
wire            n25168;
wire            n25169;
wire            n2517;
wire            n25170;
wire            n25171;
wire      [7:0] n25172;
wire            n25173;
wire            n25174;
wire            n25175;
wire            n25176;
wire            n25177;
wire      [7:0] n25178;
wire            n25179;
wire            n2518;
wire            n25180;
wire            n25181;
wire            n25182;
wire            n25183;
wire      [7:0] n25184;
wire            n25185;
wire            n25186;
wire            n25187;
wire            n25188;
wire            n25189;
wire            n2519;
wire      [7:0] n25190;
wire            n25191;
wire            n25192;
wire            n25193;
wire            n25194;
wire            n25195;
wire      [7:0] n25196;
wire            n25197;
wire            n25198;
wire            n25199;
wire            n252;
wire            n2520;
wire            n25200;
wire            n25201;
wire      [7:0] n25202;
wire            n25203;
wire            n25204;
wire            n25205;
wire            n25206;
wire            n25207;
wire      [7:0] n25208;
wire            n25209;
wire            n2521;
wire            n25210;
wire            n25211;
wire            n25212;
wire            n25213;
wire      [7:0] n25214;
wire            n25215;
wire            n25216;
wire            n25217;
wire            n25218;
wire            n25219;
wire            n2522;
wire      [7:0] n25220;
wire            n25221;
wire            n25222;
wire            n25223;
wire            n25224;
wire            n25225;
wire      [7:0] n25226;
wire            n25227;
wire            n25228;
wire            n25229;
wire            n2523;
wire            n25230;
wire            n25231;
wire      [7:0] n25232;
wire            n25233;
wire            n25234;
wire            n25235;
wire            n25236;
wire            n25237;
wire      [7:0] n25238;
wire            n25239;
wire            n2524;
wire            n25240;
wire            n25241;
wire            n25242;
wire            n25243;
wire      [7:0] n25244;
wire            n25245;
wire            n25246;
wire            n25247;
wire            n25248;
wire            n25249;
wire            n2525;
wire      [7:0] n25250;
wire            n25251;
wire            n25252;
wire            n25253;
wire            n25254;
wire            n25255;
wire      [7:0] n25256;
wire            n25257;
wire            n25258;
wire            n25259;
wire            n2526;
wire            n25260;
wire            n25261;
wire      [7:0] n25262;
wire            n25263;
wire            n25264;
wire            n25265;
wire            n25266;
wire            n25267;
wire      [7:0] n25268;
wire            n25269;
wire            n2527;
wire            n25270;
wire            n25271;
wire            n25272;
wire            n25273;
wire      [7:0] n25274;
wire            n25275;
wire            n25276;
wire            n25277;
wire            n25278;
wire            n25279;
wire            n2528;
wire      [7:0] n25280;
wire            n25281;
wire            n25282;
wire            n25283;
wire            n25284;
wire            n25285;
wire      [7:0] n25286;
wire            n25287;
wire            n25288;
wire            n25289;
wire            n2529;
wire            n25290;
wire            n25291;
wire      [7:0] n25292;
wire            n25293;
wire            n25294;
wire            n25295;
wire            n25296;
wire            n25297;
wire      [7:0] n25298;
wire            n25299;
wire            n2530;
wire            n25300;
wire            n25301;
wire            n25302;
wire            n25303;
wire      [7:0] n25304;
wire            n25305;
wire            n25306;
wire            n25307;
wire            n25308;
wire            n25309;
wire            n2531;
wire      [7:0] n25310;
wire            n25311;
wire            n25312;
wire            n25313;
wire            n25314;
wire            n25315;
wire      [7:0] n25316;
wire            n25317;
wire            n25318;
wire            n25319;
wire            n2532;
wire            n25320;
wire            n25321;
wire      [7:0] n25322;
wire            n25323;
wire            n25324;
wire            n25325;
wire            n25326;
wire            n25327;
wire      [7:0] n25328;
wire            n25329;
wire            n2533;
wire            n25330;
wire            n25331;
wire            n25332;
wire            n25333;
wire      [7:0] n25334;
wire            n25335;
wire            n25336;
wire            n25337;
wire            n25338;
wire            n25339;
wire            n2534;
wire      [7:0] n25340;
wire            n25341;
wire            n25342;
wire            n25343;
wire            n25344;
wire            n25345;
wire      [7:0] n25346;
wire            n25347;
wire            n25348;
wire            n25349;
wire            n2535;
wire            n25350;
wire            n25351;
wire      [7:0] n25352;
wire            n25353;
wire            n25354;
wire            n25355;
wire            n25356;
wire            n25357;
wire      [7:0] n25358;
wire            n25359;
wire            n2536;
wire            n25360;
wire            n25361;
wire            n25362;
wire            n25363;
wire      [7:0] n25364;
wire            n25365;
wire            n25366;
wire            n25367;
wire            n25368;
wire            n25369;
wire            n2537;
wire      [7:0] n25370;
wire            n25371;
wire            n25372;
wire            n25373;
wire            n25374;
wire            n25375;
wire      [7:0] n25376;
wire            n25377;
wire            n25378;
wire            n25379;
wire            n2538;
wire            n25380;
wire            n25381;
wire      [7:0] n25382;
wire            n25383;
wire            n25384;
wire            n25385;
wire            n25386;
wire            n25387;
wire      [7:0] n25388;
wire            n25389;
wire            n2539;
wire            n25390;
wire            n25391;
wire            n25392;
wire            n25393;
wire      [7:0] n25394;
wire            n25395;
wire            n25396;
wire            n25397;
wire            n25398;
wire            n25399;
wire            n254;
wire            n2540;
wire      [7:0] n25400;
wire            n25401;
wire            n25402;
wire            n25403;
wire            n25404;
wire            n25405;
wire      [7:0] n25406;
wire            n25407;
wire            n25408;
wire            n25409;
wire            n2541;
wire            n25410;
wire            n25411;
wire      [7:0] n25412;
wire            n25413;
wire            n25414;
wire            n25415;
wire            n25416;
wire            n25417;
wire      [7:0] n25418;
wire            n25419;
wire            n2542;
wire            n25420;
wire            n25421;
wire            n25422;
wire            n25423;
wire      [7:0] n25424;
wire            n25425;
wire            n25426;
wire            n25427;
wire            n25428;
wire            n25429;
wire            n2543;
wire      [7:0] n25430;
wire            n25431;
wire            n25432;
wire            n25433;
wire            n25434;
wire            n25435;
wire      [7:0] n25436;
wire            n25437;
wire            n25438;
wire            n25439;
wire            n2544;
wire            n25440;
wire            n25441;
wire      [7:0] n25442;
wire            n25443;
wire            n25444;
wire            n25445;
wire            n25446;
wire            n25447;
wire      [7:0] n25448;
wire            n25449;
wire            n2545;
wire            n25450;
wire            n25451;
wire            n25452;
wire            n25453;
wire      [7:0] n25454;
wire            n25455;
wire            n25456;
wire            n25457;
wire            n25458;
wire            n25459;
wire            n2546;
wire      [7:0] n25460;
wire            n25461;
wire            n25462;
wire            n25463;
wire            n25464;
wire            n25465;
wire      [7:0] n25466;
wire            n25467;
wire            n25468;
wire            n25469;
wire            n2547;
wire            n25470;
wire            n25471;
wire      [7:0] n25472;
wire            n25473;
wire            n25474;
wire            n25475;
wire            n25476;
wire            n25477;
wire      [7:0] n25478;
wire            n25479;
wire            n2548;
wire            n25480;
wire            n25481;
wire            n25482;
wire            n25483;
wire      [7:0] n25484;
wire            n25485;
wire            n25486;
wire            n25487;
wire            n25488;
wire            n25489;
wire            n2549;
wire      [7:0] n25490;
wire            n25491;
wire            n25492;
wire            n25493;
wire            n25494;
wire            n25495;
wire      [7:0] n25496;
wire            n25497;
wire            n25498;
wire            n25499;
wire            n2550;
wire            n25500;
wire            n25501;
wire      [7:0] n25502;
wire            n25503;
wire            n25504;
wire            n25505;
wire            n25506;
wire            n25507;
wire      [7:0] n25508;
wire            n25509;
wire            n2551;
wire            n25510;
wire            n25511;
wire            n25512;
wire            n25513;
wire      [7:0] n25514;
wire            n25515;
wire            n25516;
wire            n25517;
wire            n25518;
wire            n25519;
wire            n2552;
wire      [7:0] n25520;
wire            n25521;
wire            n25522;
wire            n25523;
wire            n25524;
wire            n25525;
wire      [7:0] n25526;
wire            n25527;
wire            n25528;
wire            n25529;
wire            n2553;
wire            n25530;
wire            n25531;
wire      [7:0] n25532;
wire            n25533;
wire            n25534;
wire            n25535;
wire            n25536;
wire            n25537;
wire      [7:0] n25538;
wire            n25539;
wire            n2554;
wire            n25540;
wire            n25541;
wire            n25542;
wire            n25543;
wire      [7:0] n25544;
wire            n25545;
wire            n25546;
wire            n25547;
wire            n25548;
wire            n25549;
wire            n2555;
wire      [7:0] n25550;
wire            n25551;
wire            n25552;
wire            n25553;
wire            n25554;
wire            n25555;
wire      [7:0] n25556;
wire            n25557;
wire            n25558;
wire            n25559;
wire            n2556;
wire            n25560;
wire            n25561;
wire      [7:0] n25562;
wire            n25563;
wire            n25564;
wire            n25565;
wire            n25566;
wire            n25567;
wire      [7:0] n25568;
wire            n25569;
wire            n2557;
wire            n25570;
wire            n25571;
wire            n25572;
wire            n25573;
wire      [7:0] n25574;
wire            n25575;
wire            n25576;
wire            n25577;
wire            n25578;
wire            n25579;
wire            n2558;
wire      [7:0] n25580;
wire            n25581;
wire            n25582;
wire            n25583;
wire            n25584;
wire            n25585;
wire      [7:0] n25586;
wire            n25587;
wire            n25588;
wire            n25589;
wire            n2559;
wire            n25590;
wire            n25591;
wire      [7:0] n25592;
wire            n25593;
wire            n25594;
wire            n25595;
wire            n25596;
wire            n25597;
wire      [7:0] n25598;
wire            n25599;
wire            n256;
wire            n2560;
wire            n25600;
wire            n25601;
wire            n25602;
wire            n25603;
wire      [7:0] n25604;
wire            n25605;
wire            n25606;
wire            n25607;
wire            n25608;
wire            n25609;
wire            n2561;
wire      [7:0] n25610;
wire            n25611;
wire            n25612;
wire            n25613;
wire            n25614;
wire            n25615;
wire      [7:0] n25616;
wire            n25617;
wire            n25618;
wire            n25619;
wire            n2562;
wire            n25620;
wire            n25621;
wire      [7:0] n25622;
wire            n25623;
wire            n25624;
wire            n25625;
wire            n25626;
wire            n25627;
wire      [7:0] n25628;
wire            n25629;
wire            n2563;
wire            n25630;
wire            n25631;
wire            n25632;
wire            n25633;
wire      [7:0] n25634;
wire            n25635;
wire            n25636;
wire            n25637;
wire            n25638;
wire            n25639;
wire            n2564;
wire      [7:0] n25640;
wire            n25641;
wire            n25642;
wire            n25643;
wire            n25644;
wire            n25645;
wire      [7:0] n25646;
wire            n25647;
wire            n25648;
wire            n25649;
wire            n2565;
wire            n25650;
wire            n25651;
wire      [7:0] n25652;
wire            n25653;
wire            n25654;
wire            n25655;
wire            n25656;
wire            n25657;
wire      [7:0] n25658;
wire            n25659;
wire            n2566;
wire            n25660;
wire            n25661;
wire            n25662;
wire            n25663;
wire      [7:0] n25664;
wire            n25665;
wire            n25666;
wire            n25667;
wire            n25668;
wire            n25669;
wire            n2567;
wire      [7:0] n25670;
wire            n25671;
wire            n25672;
wire            n25673;
wire            n25674;
wire            n25675;
wire      [7:0] n25676;
wire            n25677;
wire            n25678;
wire            n25679;
wire            n2568;
wire            n25680;
wire            n25681;
wire      [7:0] n25682;
wire            n25683;
wire            n25684;
wire            n25685;
wire            n25686;
wire            n25687;
wire      [7:0] n25688;
wire            n25689;
wire            n2569;
wire            n25690;
wire            n25691;
wire            n25692;
wire            n25693;
wire      [7:0] n25694;
wire            n25695;
wire            n25696;
wire            n25697;
wire            n25698;
wire            n25699;
wire            n2570;
wire      [7:0] n25700;
wire            n25701;
wire            n25702;
wire            n25703;
wire            n25704;
wire            n25705;
wire      [7:0] n25706;
wire            n25707;
wire            n25708;
wire            n25709;
wire            n2571;
wire            n25710;
wire            n25711;
wire      [7:0] n25712;
wire            n25713;
wire            n25714;
wire            n25715;
wire            n25716;
wire            n25717;
wire      [7:0] n25718;
wire            n25719;
wire            n2572;
wire            n25720;
wire            n25721;
wire            n25722;
wire            n25723;
wire      [7:0] n25724;
wire            n25725;
wire            n25726;
wire            n25727;
wire            n25728;
wire            n25729;
wire            n2573;
wire      [7:0] n25730;
wire            n25731;
wire            n25732;
wire            n25733;
wire            n25734;
wire            n25735;
wire      [7:0] n25736;
wire            n25737;
wire            n25738;
wire            n25739;
wire            n2574;
wire            n25740;
wire            n25741;
wire      [7:0] n25742;
wire            n25743;
wire            n25744;
wire            n25745;
wire            n25746;
wire            n25747;
wire      [7:0] n25748;
wire            n25749;
wire            n2575;
wire            n25750;
wire            n25751;
wire            n25752;
wire            n25753;
wire      [7:0] n25754;
wire            n25755;
wire            n25756;
wire            n25757;
wire            n25758;
wire            n25759;
wire            n2576;
wire      [7:0] n25760;
wire            n25761;
wire            n25762;
wire            n25763;
wire            n25764;
wire            n25765;
wire      [7:0] n25766;
wire            n25767;
wire            n25768;
wire            n25769;
wire            n2577;
wire            n25770;
wire            n25771;
wire      [7:0] n25772;
wire            n25773;
wire            n25774;
wire            n25775;
wire            n25776;
wire            n25777;
wire      [7:0] n25778;
wire            n25779;
wire            n2578;
wire            n25780;
wire            n25781;
wire            n25782;
wire            n25783;
wire      [7:0] n25784;
wire            n25785;
wire            n25786;
wire            n25787;
wire            n25788;
wire            n25789;
wire            n2579;
wire      [7:0] n25790;
wire            n25791;
wire            n25792;
wire            n25793;
wire            n25794;
wire            n25795;
wire      [7:0] n25796;
wire            n25797;
wire            n25798;
wire            n25799;
wire            n258;
wire            n2580;
wire            n25800;
wire            n25801;
wire      [7:0] n25802;
wire            n25803;
wire            n25804;
wire            n25805;
wire            n25806;
wire            n25807;
wire      [7:0] n25808;
wire            n25809;
wire            n2581;
wire            n25810;
wire            n25811;
wire            n25812;
wire            n25813;
wire      [7:0] n25814;
wire            n25815;
wire            n25816;
wire            n25817;
wire            n25818;
wire            n25819;
wire            n2582;
wire      [7:0] n25820;
wire            n25821;
wire            n25822;
wire            n25823;
wire            n25824;
wire            n25825;
wire      [7:0] n25826;
wire            n25827;
wire            n25828;
wire            n25829;
wire            n2583;
wire            n25830;
wire            n25831;
wire      [7:0] n25832;
wire            n25833;
wire            n25834;
wire            n25835;
wire            n25836;
wire            n25837;
wire      [7:0] n25838;
wire            n25839;
wire            n2584;
wire            n25840;
wire            n25841;
wire            n25842;
wire            n25843;
wire      [7:0] n25844;
wire            n25845;
wire            n25846;
wire            n25847;
wire            n25848;
wire            n25849;
wire            n2585;
wire      [7:0] n25850;
wire            n25851;
wire            n25852;
wire            n25853;
wire            n25854;
wire            n25855;
wire      [7:0] n25856;
wire            n25857;
wire            n25858;
wire            n25859;
wire            n2586;
wire            n25860;
wire            n25861;
wire      [7:0] n25862;
wire            n25863;
wire            n25864;
wire            n25865;
wire            n25866;
wire            n25867;
wire      [7:0] n25868;
wire            n25869;
wire            n2587;
wire            n25870;
wire            n25871;
wire            n25872;
wire            n25873;
wire      [7:0] n25874;
wire            n25875;
wire            n25876;
wire            n25877;
wire            n25878;
wire            n25879;
wire            n2588;
wire      [7:0] n25880;
wire            n25881;
wire            n25882;
wire            n25883;
wire            n25884;
wire            n25885;
wire      [7:0] n25886;
wire            n25887;
wire            n25888;
wire            n25889;
wire            n2589;
wire            n25890;
wire            n25891;
wire      [7:0] n25892;
wire            n25893;
wire            n25894;
wire            n25895;
wire            n25896;
wire            n25897;
wire      [7:0] n25898;
wire            n25899;
wire            n2590;
wire            n25900;
wire            n25901;
wire            n25902;
wire            n25903;
wire      [7:0] n25904;
wire            n25905;
wire            n25906;
wire            n25907;
wire            n25908;
wire            n25909;
wire            n2591;
wire      [7:0] n25910;
wire            n25911;
wire            n25912;
wire            n25913;
wire            n25914;
wire            n25915;
wire      [7:0] n25916;
wire            n25917;
wire            n25918;
wire            n25919;
wire            n2592;
wire            n25920;
wire            n25921;
wire      [7:0] n25922;
wire            n25923;
wire            n25924;
wire            n25925;
wire            n25926;
wire            n25927;
wire      [7:0] n25928;
wire            n25929;
wire            n2593;
wire            n25930;
wire            n25931;
wire            n25932;
wire            n25933;
wire      [7:0] n25934;
wire            n25935;
wire            n25936;
wire            n25937;
wire            n25938;
wire            n25939;
wire            n2594;
wire      [7:0] n25940;
wire            n25941;
wire            n25942;
wire            n25943;
wire            n25944;
wire            n25945;
wire      [7:0] n25946;
wire            n25947;
wire            n25948;
wire            n25949;
wire            n2595;
wire            n25950;
wire            n25951;
wire      [7:0] n25952;
wire            n25953;
wire            n25954;
wire            n25955;
wire            n25956;
wire            n25957;
wire      [7:0] n25958;
wire            n25959;
wire            n2596;
wire            n25960;
wire            n25961;
wire            n25962;
wire            n25963;
wire      [7:0] n25964;
wire            n25965;
wire            n25966;
wire            n25967;
wire            n25968;
wire            n25969;
wire            n2597;
wire      [7:0] n25970;
wire            n25971;
wire            n25972;
wire            n25973;
wire            n25974;
wire            n25975;
wire      [7:0] n25976;
wire            n25977;
wire            n25978;
wire            n25979;
wire            n2598;
wire            n25980;
wire            n25981;
wire      [7:0] n25982;
wire            n25983;
wire            n25984;
wire            n25985;
wire            n25986;
wire            n25987;
wire      [7:0] n25988;
wire            n25989;
wire            n2599;
wire            n25990;
wire            n25991;
wire            n25992;
wire            n25993;
wire      [7:0] n25994;
wire            n25995;
wire            n25996;
wire            n25997;
wire            n25998;
wire            n25999;
wire            n260;
wire            n2600;
wire      [7:0] n26000;
wire            n26001;
wire            n26002;
wire            n26003;
wire            n26004;
wire            n26005;
wire      [7:0] n26006;
wire            n26007;
wire            n26008;
wire            n26009;
wire            n2601;
wire            n26010;
wire            n26011;
wire      [7:0] n26012;
wire            n26013;
wire            n26014;
wire            n26015;
wire            n26016;
wire            n26017;
wire      [7:0] n26018;
wire            n26019;
wire            n2602;
wire            n26020;
wire            n26021;
wire            n26022;
wire            n26023;
wire      [7:0] n26024;
wire            n26025;
wire            n26026;
wire            n26027;
wire            n26028;
wire            n26029;
wire            n2603;
wire      [7:0] n26030;
wire            n26031;
wire            n26032;
wire            n26033;
wire            n26034;
wire            n26035;
wire      [7:0] n26036;
wire            n26037;
wire            n26038;
wire            n26039;
wire            n2604;
wire            n26040;
wire            n26041;
wire      [7:0] n26042;
wire            n26043;
wire            n26044;
wire            n26045;
wire            n26046;
wire            n26047;
wire      [7:0] n26048;
wire            n26049;
wire            n2605;
wire            n26050;
wire            n26051;
wire            n26052;
wire            n26053;
wire      [7:0] n26054;
wire            n26055;
wire            n26056;
wire            n26057;
wire            n26058;
wire            n26059;
wire            n2606;
wire      [7:0] n26060;
wire            n26061;
wire            n26062;
wire            n26063;
wire            n26064;
wire            n26065;
wire      [7:0] n26066;
wire            n26067;
wire            n26068;
wire            n26069;
wire            n2607;
wire            n26070;
wire            n26071;
wire      [7:0] n26072;
wire            n26073;
wire            n26074;
wire            n26075;
wire            n26076;
wire            n26077;
wire      [7:0] n26078;
wire            n26079;
wire            n2608;
wire            n26080;
wire            n26081;
wire            n26082;
wire            n26083;
wire      [7:0] n26084;
wire            n26085;
wire            n26086;
wire            n26087;
wire            n26088;
wire            n26089;
wire            n2609;
wire      [7:0] n26090;
wire            n26091;
wire            n26092;
wire            n26093;
wire            n26094;
wire            n26095;
wire      [7:0] n26096;
wire            n26097;
wire            n26098;
wire            n26099;
wire            n2610;
wire            n26100;
wire            n26101;
wire      [7:0] n26102;
wire            n26103;
wire            n26104;
wire            n26105;
wire            n26106;
wire            n26107;
wire      [7:0] n26108;
wire            n26109;
wire            n2611;
wire            n26110;
wire            n26111;
wire            n26112;
wire            n26113;
wire      [7:0] n26114;
wire            n26115;
wire            n26116;
wire            n26117;
wire            n26118;
wire            n26119;
wire            n2612;
wire      [7:0] n26120;
wire            n26121;
wire            n26122;
wire            n26123;
wire            n26124;
wire            n26125;
wire      [7:0] n26126;
wire            n26127;
wire            n26128;
wire            n26129;
wire            n2613;
wire            n26130;
wire            n26131;
wire      [7:0] n26132;
wire            n26133;
wire            n26134;
wire            n26135;
wire            n26136;
wire            n26137;
wire      [7:0] n26138;
wire            n26139;
wire            n2614;
wire            n26140;
wire            n26141;
wire            n26142;
wire            n26143;
wire      [7:0] n26144;
wire            n26145;
wire            n26146;
wire            n26147;
wire            n26148;
wire            n26149;
wire            n2615;
wire      [7:0] n26150;
wire            n26151;
wire            n26152;
wire            n26153;
wire            n26154;
wire            n26155;
wire      [7:0] n26156;
wire            n26157;
wire            n26158;
wire            n26159;
wire            n2616;
wire            n26160;
wire            n26161;
wire      [7:0] n26162;
wire            n26163;
wire            n26164;
wire            n26165;
wire            n26166;
wire            n26167;
wire      [7:0] n26168;
wire            n26169;
wire            n2617;
wire            n26170;
wire            n26171;
wire            n26172;
wire            n26173;
wire      [7:0] n26174;
wire            n26175;
wire            n26176;
wire            n26177;
wire            n26178;
wire            n26179;
wire            n2618;
wire      [7:0] n26180;
wire            n26181;
wire            n26182;
wire            n26183;
wire            n26184;
wire            n26185;
wire      [7:0] n26186;
wire            n26187;
wire            n26188;
wire            n26189;
wire            n2619;
wire            n26190;
wire            n26191;
wire      [7:0] n26192;
wire            n26193;
wire            n26194;
wire            n26195;
wire            n26196;
wire            n26197;
wire      [7:0] n26198;
wire            n26199;
wire            n262;
wire            n2620;
wire            n26200;
wire            n26201;
wire            n26202;
wire            n26203;
wire      [7:0] n26204;
wire            n26205;
wire            n26206;
wire            n26207;
wire            n26208;
wire            n26209;
wire            n2621;
wire      [7:0] n26210;
wire            n26211;
wire            n26212;
wire            n26213;
wire            n26214;
wire            n26215;
wire      [7:0] n26216;
wire            n26217;
wire            n26218;
wire            n26219;
wire            n2622;
wire            n26220;
wire            n26221;
wire      [7:0] n26222;
wire            n26223;
wire            n26224;
wire            n26225;
wire            n26226;
wire            n26227;
wire      [7:0] n26228;
wire            n26229;
wire            n2623;
wire            n26230;
wire            n26231;
wire            n26232;
wire            n26233;
wire      [7:0] n26234;
wire            n26235;
wire            n26236;
wire            n26237;
wire            n26238;
wire            n26239;
wire            n2624;
wire      [7:0] n26240;
wire            n26241;
wire            n26242;
wire            n26243;
wire            n26244;
wire            n26245;
wire      [7:0] n26246;
wire            n26247;
wire            n26248;
wire            n26249;
wire            n2625;
wire            n26250;
wire            n26251;
wire      [7:0] n26252;
wire            n26253;
wire            n26254;
wire            n26255;
wire            n26256;
wire            n26257;
wire      [7:0] n26258;
wire            n26259;
wire            n2626;
wire            n26260;
wire            n26261;
wire            n26262;
wire            n26263;
wire      [7:0] n26264;
wire            n26265;
wire            n26266;
wire            n26267;
wire            n26268;
wire            n26269;
wire            n2627;
wire      [7:0] n26270;
wire            n26271;
wire            n26272;
wire            n26273;
wire            n26274;
wire            n26275;
wire      [7:0] n26276;
wire            n26277;
wire            n26278;
wire            n26279;
wire            n2628;
wire            n26280;
wire            n26281;
wire      [7:0] n26282;
wire            n26283;
wire            n26284;
wire            n26285;
wire            n26286;
wire            n26287;
wire      [7:0] n26288;
wire            n26289;
wire            n2629;
wire            n26290;
wire            n26291;
wire            n26292;
wire            n26293;
wire      [7:0] n26294;
wire            n26295;
wire            n26296;
wire            n26297;
wire            n26298;
wire            n26299;
wire            n2630;
wire      [7:0] n26300;
wire            n26301;
wire            n26302;
wire            n26303;
wire            n26304;
wire            n26305;
wire      [7:0] n26306;
wire            n26307;
wire            n26308;
wire            n26309;
wire            n2631;
wire            n26310;
wire            n26311;
wire      [7:0] n26312;
wire            n26313;
wire            n26314;
wire            n26315;
wire            n26316;
wire            n26317;
wire      [7:0] n26318;
wire            n26319;
wire            n2632;
wire            n26320;
wire            n26321;
wire            n26322;
wire            n26323;
wire      [7:0] n26324;
wire            n26325;
wire            n26326;
wire            n26327;
wire            n26328;
wire            n26329;
wire            n2633;
wire      [7:0] n26330;
wire            n26331;
wire            n26332;
wire            n26333;
wire            n26334;
wire            n26335;
wire      [7:0] n26336;
wire            n26337;
wire            n26338;
wire            n26339;
wire            n2634;
wire            n26340;
wire            n26341;
wire      [7:0] n26342;
wire            n26343;
wire            n26344;
wire            n26345;
wire            n26346;
wire            n26347;
wire      [7:0] n26348;
wire            n26349;
wire            n2635;
wire            n26350;
wire            n26351;
wire            n26352;
wire            n26353;
wire      [7:0] n26354;
wire            n26355;
wire            n26356;
wire            n26357;
wire            n26358;
wire            n26359;
wire            n2636;
wire      [7:0] n26360;
wire            n26361;
wire            n26362;
wire            n26363;
wire            n26364;
wire            n26365;
wire      [7:0] n26366;
wire            n26367;
wire            n26368;
wire            n26369;
wire            n2637;
wire            n26370;
wire            n26371;
wire      [7:0] n26372;
wire            n26373;
wire            n26374;
wire            n26375;
wire            n26376;
wire            n26377;
wire      [7:0] n26378;
wire            n26379;
wire            n2638;
wire            n26380;
wire            n26381;
wire            n26382;
wire            n26383;
wire      [7:0] n26384;
wire            n26385;
wire            n26386;
wire            n26387;
wire            n26388;
wire            n26389;
wire            n2639;
wire      [7:0] n26390;
wire            n26391;
wire            n26392;
wire            n26393;
wire            n26394;
wire            n26395;
wire      [7:0] n26396;
wire            n26397;
wire            n26398;
wire            n26399;
wire            n264;
wire            n2640;
wire            n26400;
wire            n26401;
wire      [7:0] n26402;
wire            n26403;
wire            n26404;
wire            n26405;
wire            n26406;
wire            n26407;
wire      [7:0] n26408;
wire            n26409;
wire            n2641;
wire            n26410;
wire            n26411;
wire            n26412;
wire            n26413;
wire      [7:0] n26414;
wire            n26415;
wire            n26416;
wire            n26417;
wire            n26418;
wire            n26419;
wire            n2642;
wire      [7:0] n26420;
wire            n26421;
wire            n26422;
wire            n26423;
wire            n26424;
wire            n26425;
wire      [7:0] n26426;
wire            n26427;
wire            n26428;
wire            n26429;
wire            n2643;
wire            n26430;
wire            n26431;
wire      [7:0] n26432;
wire            n26433;
wire            n26434;
wire            n26435;
wire            n26436;
wire            n26437;
wire      [7:0] n26438;
wire            n26439;
wire            n2644;
wire            n26440;
wire            n26441;
wire            n26442;
wire            n26443;
wire      [7:0] n26444;
wire            n26445;
wire            n26446;
wire            n26447;
wire            n26448;
wire            n26449;
wire            n2645;
wire      [7:0] n26450;
wire            n26451;
wire            n26452;
wire            n26453;
wire            n26454;
wire            n26455;
wire      [7:0] n26456;
wire            n26457;
wire            n26458;
wire            n26459;
wire            n2646;
wire            n26460;
wire            n26461;
wire      [7:0] n26462;
wire            n26463;
wire            n26464;
wire            n26465;
wire            n26466;
wire            n26467;
wire      [7:0] n26468;
wire            n26469;
wire            n2647;
wire            n26470;
wire            n26471;
wire            n26472;
wire            n26473;
wire      [7:0] n26474;
wire            n26475;
wire            n26476;
wire            n26477;
wire            n26478;
wire            n26479;
wire            n2648;
wire      [7:0] n26480;
wire            n26481;
wire            n26482;
wire            n26483;
wire            n26484;
wire            n26485;
wire      [7:0] n26486;
wire            n26487;
wire            n26488;
wire            n26489;
wire            n2649;
wire            n26490;
wire            n26491;
wire      [7:0] n26492;
wire            n26493;
wire            n26494;
wire            n26495;
wire            n26496;
wire            n26497;
wire      [7:0] n26498;
wire            n26499;
wire            n2650;
wire            n26500;
wire            n26501;
wire            n26502;
wire            n26503;
wire      [7:0] n26504;
wire            n26505;
wire            n26506;
wire            n26507;
wire            n26508;
wire            n26509;
wire            n2651;
wire      [7:0] n26510;
wire            n26511;
wire            n26512;
wire            n26513;
wire            n26514;
wire            n26515;
wire      [7:0] n26516;
wire            n26517;
wire            n26518;
wire            n26519;
wire            n2652;
wire            n26520;
wire            n26521;
wire      [7:0] n26522;
wire            n26523;
wire            n26524;
wire            n26525;
wire            n26526;
wire            n26527;
wire      [7:0] n26528;
wire            n26529;
wire            n2653;
wire            n26530;
wire            n26531;
wire            n26532;
wire            n26533;
wire      [7:0] n26534;
wire            n26535;
wire            n26536;
wire            n26537;
wire            n26538;
wire            n26539;
wire            n2654;
wire      [7:0] n26540;
wire            n26541;
wire            n26542;
wire            n26543;
wire            n26544;
wire            n26545;
wire      [7:0] n26546;
wire            n26547;
wire            n26548;
wire            n26549;
wire            n2655;
wire            n26550;
wire            n26551;
wire      [7:0] n26552;
wire            n26553;
wire            n26554;
wire            n26555;
wire            n26556;
wire            n26557;
wire      [7:0] n26558;
wire            n26559;
wire            n2656;
wire            n26560;
wire            n26561;
wire            n26562;
wire            n26563;
wire      [7:0] n26564;
wire            n26565;
wire            n26566;
wire            n26567;
wire            n26568;
wire            n26569;
wire            n2657;
wire      [7:0] n26570;
wire            n26571;
wire            n26572;
wire            n26573;
wire            n26574;
wire            n26575;
wire      [7:0] n26576;
wire            n26577;
wire            n26578;
wire            n26579;
wire            n2658;
wire            n26580;
wire            n26581;
wire      [7:0] n26582;
wire            n26583;
wire            n26584;
wire            n26585;
wire            n26586;
wire            n26587;
wire      [7:0] n26588;
wire            n26589;
wire            n2659;
wire            n26590;
wire            n26591;
wire            n26592;
wire            n26593;
wire      [7:0] n26594;
wire            n26595;
wire            n26596;
wire            n26597;
wire            n26598;
wire            n26599;
wire            n266;
wire      [7:0] n2660;
wire      [7:0] n26600;
wire            n26601;
wire            n26602;
wire            n26603;
wire            n26604;
wire            n26605;
wire      [7:0] n26606;
wire            n26607;
wire            n26608;
wire            n26609;
wire      [7:0] n2661;
wire            n26610;
wire            n26611;
wire      [7:0] n26612;
wire            n26613;
wire            n26614;
wire            n26615;
wire            n26616;
wire            n26617;
wire      [7:0] n26618;
wire            n26619;
wire      [7:0] n2662;
wire            n26620;
wire            n26621;
wire            n26622;
wire            n26623;
wire      [7:0] n26624;
wire            n26625;
wire            n26626;
wire            n26627;
wire            n26628;
wire            n26629;
wire      [7:0] n2663;
wire      [7:0] n26630;
wire            n26631;
wire            n26632;
wire            n26633;
wire            n26634;
wire            n26635;
wire      [7:0] n26636;
wire            n26637;
wire            n26638;
wire            n26639;
wire      [7:0] n2664;
wire            n26640;
wire            n26641;
wire      [7:0] n26642;
wire            n26643;
wire            n26644;
wire            n26645;
wire            n26646;
wire            n26647;
wire      [7:0] n26648;
wire            n26649;
wire      [7:0] n2665;
wire            n26650;
wire            n26651;
wire            n26652;
wire            n26653;
wire      [7:0] n26654;
wire            n26655;
wire            n26656;
wire            n26657;
wire            n26658;
wire            n26659;
wire      [7:0] n2666;
wire      [7:0] n26660;
wire            n26661;
wire            n26662;
wire            n26663;
wire            n26664;
wire            n26665;
wire      [7:0] n26666;
wire            n26667;
wire            n26668;
wire            n26669;
wire      [7:0] n2667;
wire            n26670;
wire            n26671;
wire      [7:0] n26672;
wire            n26673;
wire            n26674;
wire            n26675;
wire            n26676;
wire            n26677;
wire      [7:0] n26678;
wire            n26679;
wire      [7:0] n2668;
wire            n26680;
wire            n26681;
wire            n26682;
wire            n26683;
wire      [7:0] n26684;
wire            n26685;
wire            n26686;
wire            n26687;
wire            n26688;
wire            n26689;
wire      [7:0] n2669;
wire      [7:0] n26690;
wire            n26691;
wire            n26692;
wire            n26693;
wire            n26694;
wire            n26695;
wire      [7:0] n26696;
wire            n26697;
wire            n26698;
wire            n26699;
wire      [7:0] n2670;
wire            n26700;
wire            n26701;
wire      [7:0] n26702;
wire            n26703;
wire            n26704;
wire            n26705;
wire            n26706;
wire            n26707;
wire      [7:0] n26708;
wire            n26709;
wire      [7:0] n2671;
wire            n26710;
wire            n26711;
wire            n26712;
wire            n26713;
wire      [7:0] n26714;
wire            n26715;
wire            n26716;
wire            n26717;
wire            n26718;
wire            n26719;
wire      [7:0] n2672;
wire      [7:0] n26720;
wire            n26721;
wire            n26722;
wire            n26723;
wire            n26724;
wire            n26725;
wire      [7:0] n26726;
wire            n26727;
wire            n26728;
wire            n26729;
wire      [7:0] n2673;
wire            n26730;
wire            n26731;
wire      [7:0] n26732;
wire            n26733;
wire            n26734;
wire            n26735;
wire            n26736;
wire            n26737;
wire      [7:0] n26738;
wire            n26739;
wire      [7:0] n2674;
wire            n26740;
wire            n26741;
wire            n26742;
wire            n26743;
wire      [7:0] n26744;
wire            n26745;
wire            n26746;
wire            n26747;
wire            n26748;
wire            n26749;
wire      [7:0] n2675;
wire      [7:0] n26750;
wire            n26751;
wire            n26752;
wire            n26753;
wire            n26754;
wire            n26755;
wire      [7:0] n26756;
wire            n26757;
wire            n26758;
wire            n26759;
wire      [7:0] n2676;
wire            n26760;
wire            n26761;
wire      [7:0] n26762;
wire            n26763;
wire            n26764;
wire            n26765;
wire            n26766;
wire            n26767;
wire      [7:0] n26768;
wire            n26769;
wire      [7:0] n2677;
wire            n26770;
wire            n26771;
wire            n26772;
wire            n26773;
wire      [7:0] n26774;
wire            n26775;
wire            n26776;
wire            n26777;
wire            n26778;
wire            n26779;
wire      [7:0] n2678;
wire      [7:0] n26780;
wire            n26781;
wire            n26782;
wire            n26783;
wire            n26784;
wire            n26785;
wire      [7:0] n26786;
wire            n26787;
wire            n26788;
wire            n26789;
wire      [7:0] n2679;
wire            n26790;
wire            n26791;
wire      [7:0] n26792;
wire            n26793;
wire            n26794;
wire            n26795;
wire            n26796;
wire            n26797;
wire      [7:0] n26798;
wire            n26799;
wire            n268;
wire      [7:0] n2680;
wire            n26800;
wire            n26801;
wire            n26802;
wire            n26803;
wire      [7:0] n26804;
wire            n26805;
wire            n26806;
wire            n26807;
wire            n26808;
wire            n26809;
wire      [7:0] n2681;
wire      [7:0] n26810;
wire            n26811;
wire            n26812;
wire            n26813;
wire            n26814;
wire            n26815;
wire      [7:0] n26816;
wire            n26817;
wire            n26818;
wire            n26819;
wire      [7:0] n2682;
wire            n26820;
wire            n26821;
wire      [7:0] n26822;
wire            n26823;
wire            n26824;
wire            n26825;
wire            n26826;
wire            n26827;
wire      [7:0] n26828;
wire            n26829;
wire      [7:0] n2683;
wire            n26830;
wire            n26831;
wire            n26832;
wire            n26833;
wire      [7:0] n26834;
wire            n26835;
wire            n26836;
wire            n26837;
wire            n26838;
wire            n26839;
wire      [7:0] n2684;
wire      [7:0] n26840;
wire            n26841;
wire            n26842;
wire            n26843;
wire            n26844;
wire            n26845;
wire      [7:0] n26846;
wire            n26847;
wire            n26848;
wire            n26849;
wire      [7:0] n2685;
wire            n26850;
wire            n26851;
wire      [7:0] n26852;
wire            n26853;
wire            n26854;
wire            n26855;
wire            n26856;
wire            n26857;
wire      [7:0] n26858;
wire            n26859;
wire      [7:0] n2686;
wire            n26860;
wire            n26861;
wire            n26862;
wire            n26863;
wire      [7:0] n26864;
wire            n26865;
wire            n26866;
wire            n26867;
wire            n26868;
wire            n26869;
wire      [7:0] n2687;
wire      [7:0] n26870;
wire            n26871;
wire            n26872;
wire            n26873;
wire            n26874;
wire            n26875;
wire      [7:0] n26876;
wire            n26877;
wire            n26878;
wire            n26879;
wire      [7:0] n2688;
wire            n26880;
wire            n26881;
wire      [7:0] n26882;
wire            n26883;
wire            n26884;
wire            n26885;
wire            n26886;
wire            n26887;
wire      [7:0] n26888;
wire            n26889;
wire      [7:0] n2689;
wire            n26890;
wire            n26891;
wire            n26892;
wire            n26893;
wire      [7:0] n26894;
wire            n26895;
wire            n26896;
wire            n26897;
wire            n26898;
wire            n26899;
wire      [7:0] n2690;
wire      [7:0] n26900;
wire            n26901;
wire            n26902;
wire            n26903;
wire            n26904;
wire            n26905;
wire      [7:0] n26906;
wire            n26907;
wire            n26908;
wire            n26909;
wire      [7:0] n2691;
wire            n26910;
wire            n26911;
wire      [7:0] n26912;
wire            n26913;
wire            n26914;
wire            n26915;
wire            n26916;
wire            n26917;
wire      [7:0] n26918;
wire            n26919;
wire      [7:0] n2692;
wire            n26920;
wire            n26921;
wire            n26922;
wire            n26923;
wire      [7:0] n26924;
wire            n26925;
wire            n26926;
wire            n26927;
wire            n26928;
wire            n26929;
wire      [7:0] n2693;
wire      [7:0] n26930;
wire            n26931;
wire            n26932;
wire            n26933;
wire            n26934;
wire            n26935;
wire      [7:0] n26936;
wire            n26937;
wire            n26938;
wire            n26939;
wire      [7:0] n2694;
wire            n26940;
wire            n26941;
wire      [7:0] n26942;
wire            n26943;
wire            n26944;
wire            n26945;
wire            n26946;
wire            n26947;
wire      [7:0] n26948;
wire            n26949;
wire      [7:0] n2695;
wire            n26950;
wire            n26951;
wire            n26952;
wire            n26953;
wire      [7:0] n26954;
wire            n26955;
wire            n26956;
wire            n26957;
wire            n26958;
wire            n26959;
wire      [7:0] n2696;
wire      [7:0] n26960;
wire            n26961;
wire            n26962;
wire            n26963;
wire            n26964;
wire            n26965;
wire      [7:0] n26966;
wire            n26967;
wire            n26968;
wire            n26969;
wire      [7:0] n2697;
wire            n26970;
wire            n26971;
wire      [7:0] n26972;
wire            n26973;
wire            n26974;
wire            n26975;
wire            n26976;
wire            n26977;
wire      [7:0] n26978;
wire            n26979;
wire      [7:0] n2698;
wire            n26980;
wire            n26981;
wire            n26982;
wire            n26983;
wire      [7:0] n26984;
wire            n26985;
wire            n26986;
wire            n26987;
wire            n26988;
wire            n26989;
wire      [7:0] n2699;
wire      [7:0] n26990;
wire            n26991;
wire            n26992;
wire            n26993;
wire            n26994;
wire            n26995;
wire      [7:0] n26996;
wire            n26997;
wire            n26998;
wire            n26999;
wire            n27;
wire            n270;
wire      [7:0] n2700;
wire            n27000;
wire            n27001;
wire      [7:0] n27002;
wire            n27003;
wire            n27004;
wire            n27005;
wire            n27006;
wire            n27007;
wire      [7:0] n27008;
wire            n27009;
wire      [7:0] n2701;
wire            n27010;
wire            n27011;
wire            n27012;
wire            n27013;
wire      [7:0] n27014;
wire            n27015;
wire            n27016;
wire            n27017;
wire            n27018;
wire            n27019;
wire      [7:0] n2702;
wire      [7:0] n27020;
wire            n27021;
wire            n27022;
wire            n27023;
wire            n27024;
wire            n27025;
wire      [7:0] n27026;
wire            n27027;
wire            n27028;
wire            n27029;
wire      [7:0] n2703;
wire            n27030;
wire            n27031;
wire      [7:0] n27032;
wire            n27033;
wire            n27034;
wire            n27035;
wire            n27036;
wire            n27037;
wire      [7:0] n27038;
wire            n27039;
wire      [7:0] n2704;
wire            n27040;
wire            n27041;
wire            n27042;
wire            n27043;
wire      [7:0] n27044;
wire            n27045;
wire            n27046;
wire            n27047;
wire            n27048;
wire            n27049;
wire      [7:0] n2705;
wire      [7:0] n27050;
wire            n27051;
wire            n27052;
wire            n27053;
wire            n27054;
wire            n27055;
wire      [7:0] n27056;
wire            n27057;
wire            n27058;
wire            n27059;
wire      [7:0] n2706;
wire            n27060;
wire            n27061;
wire      [7:0] n27062;
wire            n27063;
wire            n27064;
wire            n27065;
wire            n27066;
wire            n27067;
wire      [7:0] n27068;
wire            n27069;
wire      [7:0] n2707;
wire            n27070;
wire            n27071;
wire            n27072;
wire            n27073;
wire      [7:0] n27074;
wire            n27075;
wire            n27076;
wire            n27077;
wire            n27078;
wire            n27079;
wire      [7:0] n2708;
wire      [7:0] n27080;
wire            n27081;
wire            n27082;
wire            n27083;
wire            n27084;
wire            n27085;
wire      [7:0] n27086;
wire            n27087;
wire            n27088;
wire            n27089;
wire      [7:0] n2709;
wire            n27090;
wire            n27091;
wire      [7:0] n27092;
wire            n27093;
wire            n27094;
wire            n27095;
wire            n27096;
wire            n27097;
wire      [7:0] n27098;
wire            n27099;
wire      [7:0] n2710;
wire            n27100;
wire            n27101;
wire            n27102;
wire            n27103;
wire      [7:0] n27104;
wire            n27105;
wire            n27106;
wire            n27107;
wire            n27108;
wire            n27109;
wire      [7:0] n2711;
wire      [7:0] n27110;
wire            n27111;
wire            n27112;
wire            n27113;
wire            n27114;
wire            n27115;
wire      [7:0] n27116;
wire            n27117;
wire            n27118;
wire            n27119;
wire      [7:0] n2712;
wire            n27120;
wire            n27121;
wire      [7:0] n27122;
wire            n27123;
wire            n27124;
wire            n27125;
wire            n27126;
wire            n27127;
wire      [7:0] n27128;
wire            n27129;
wire      [7:0] n2713;
wire            n27130;
wire            n27131;
wire            n27132;
wire            n27133;
wire      [7:0] n27134;
wire            n27135;
wire            n27136;
wire            n27137;
wire            n27138;
wire            n27139;
wire      [7:0] n2714;
wire      [7:0] n27140;
wire            n27141;
wire            n27142;
wire            n27143;
wire            n27144;
wire            n27145;
wire      [7:0] n27146;
wire            n27147;
wire            n27148;
wire            n27149;
wire      [7:0] n2715;
wire            n27150;
wire            n27151;
wire      [7:0] n27152;
wire            n27153;
wire            n27154;
wire            n27155;
wire            n27156;
wire            n27157;
wire      [7:0] n27158;
wire            n27159;
wire      [7:0] n2716;
wire            n27160;
wire            n27161;
wire            n27162;
wire            n27163;
wire      [7:0] n27164;
wire            n27165;
wire            n27166;
wire            n27167;
wire            n27168;
wire            n27169;
wire      [7:0] n2717;
wire      [7:0] n27170;
wire            n27171;
wire            n27172;
wire            n27173;
wire            n27174;
wire            n27175;
wire      [7:0] n27176;
wire            n27177;
wire            n27178;
wire            n27179;
wire      [7:0] n2718;
wire            n27180;
wire            n27181;
wire      [7:0] n27182;
wire            n27183;
wire            n27184;
wire            n27185;
wire            n27186;
wire            n27187;
wire      [7:0] n27188;
wire            n27189;
wire      [7:0] n2719;
wire            n27190;
wire            n27191;
wire            n27192;
wire            n27193;
wire      [7:0] n27194;
wire            n27195;
wire            n27196;
wire            n27197;
wire            n27198;
wire            n27199;
wire            n272;
wire      [7:0] n2720;
wire      [7:0] n27200;
wire            n27201;
wire            n27202;
wire            n27203;
wire            n27204;
wire            n27205;
wire      [7:0] n27206;
wire            n27207;
wire            n27208;
wire            n27209;
wire      [7:0] n2721;
wire            n27210;
wire            n27211;
wire      [7:0] n27212;
wire            n27213;
wire            n27214;
wire            n27215;
wire            n27216;
wire            n27217;
wire      [7:0] n27218;
wire            n27219;
wire      [7:0] n2722;
wire            n27220;
wire            n27221;
wire            n27222;
wire            n27223;
wire      [7:0] n27224;
wire            n27225;
wire            n27226;
wire            n27227;
wire            n27228;
wire            n27229;
wire      [7:0] n2723;
wire      [7:0] n27230;
wire            n27231;
wire            n27232;
wire            n27233;
wire            n27234;
wire            n27235;
wire      [7:0] n27236;
wire            n27237;
wire            n27238;
wire            n27239;
wire      [7:0] n2724;
wire            n27240;
wire            n27241;
wire      [7:0] n27242;
wire            n27243;
wire            n27244;
wire            n27245;
wire            n27246;
wire            n27247;
wire      [7:0] n27248;
wire            n27249;
wire      [7:0] n2725;
wire            n27250;
wire            n27251;
wire            n27252;
wire            n27253;
wire      [7:0] n27254;
wire            n27255;
wire            n27256;
wire            n27257;
wire            n27258;
wire            n27259;
wire      [7:0] n2726;
wire      [7:0] n27260;
wire            n27261;
wire            n27262;
wire            n27263;
wire            n27264;
wire            n27265;
wire      [7:0] n27266;
wire            n27267;
wire            n27268;
wire            n27269;
wire      [7:0] n2727;
wire            n27270;
wire            n27271;
wire      [7:0] n27272;
wire            n27273;
wire            n27274;
wire            n27275;
wire            n27276;
wire            n27277;
wire      [7:0] n27278;
wire            n27279;
wire      [7:0] n2728;
wire            n27280;
wire            n27281;
wire            n27282;
wire            n27283;
wire      [7:0] n27284;
wire            n27285;
wire            n27286;
wire            n27287;
wire            n27288;
wire            n27289;
wire      [7:0] n2729;
wire      [7:0] n27290;
wire            n27291;
wire            n27292;
wire            n27293;
wire            n27294;
wire            n27295;
wire      [7:0] n27296;
wire            n27297;
wire            n27298;
wire            n27299;
wire      [7:0] n2730;
wire            n27300;
wire            n27301;
wire      [7:0] n27302;
wire            n27303;
wire            n27304;
wire            n27305;
wire            n27306;
wire            n27307;
wire      [7:0] n27308;
wire            n27309;
wire      [7:0] n2731;
wire            n27310;
wire            n27311;
wire            n27312;
wire            n27313;
wire      [7:0] n27314;
wire            n27315;
wire            n27316;
wire            n27317;
wire            n27318;
wire            n27319;
wire      [7:0] n2732;
wire      [7:0] n27320;
wire            n27321;
wire            n27322;
wire            n27323;
wire            n27324;
wire            n27325;
wire      [7:0] n27326;
wire            n27327;
wire            n27328;
wire            n27329;
wire      [7:0] n2733;
wire            n27330;
wire            n27331;
wire      [7:0] n27332;
wire            n27333;
wire            n27334;
wire            n27335;
wire            n27336;
wire            n27337;
wire      [7:0] n27338;
wire            n27339;
wire      [7:0] n2734;
wire            n27340;
wire            n27341;
wire            n27342;
wire            n27343;
wire      [7:0] n27344;
wire            n27345;
wire            n27346;
wire            n27347;
wire            n27348;
wire            n27349;
wire      [7:0] n2735;
wire      [7:0] n27350;
wire            n27351;
wire            n27352;
wire            n27353;
wire            n27354;
wire            n27355;
wire      [7:0] n27356;
wire            n27357;
wire            n27358;
wire            n27359;
wire      [7:0] n2736;
wire            n27360;
wire            n27361;
wire      [7:0] n27362;
wire            n27363;
wire            n27364;
wire            n27365;
wire            n27366;
wire            n27367;
wire      [7:0] n27368;
wire            n27369;
wire      [7:0] n2737;
wire            n27370;
wire            n27371;
wire            n27372;
wire            n27373;
wire      [7:0] n27374;
wire            n27375;
wire            n27376;
wire            n27377;
wire            n27378;
wire            n27379;
wire      [7:0] n2738;
wire      [7:0] n27380;
wire            n27381;
wire            n27382;
wire            n27383;
wire            n27384;
wire            n27385;
wire      [7:0] n27386;
wire            n27387;
wire            n27388;
wire            n27389;
wire      [7:0] n2739;
wire            n27390;
wire            n27391;
wire      [7:0] n27392;
wire            n27393;
wire            n27394;
wire            n27395;
wire            n27396;
wire            n27397;
wire      [7:0] n27398;
wire            n27399;
wire            n274;
wire      [7:0] n2740;
wire            n27400;
wire            n27401;
wire            n27402;
wire            n27403;
wire      [7:0] n27404;
wire            n27405;
wire            n27406;
wire            n27407;
wire            n27408;
wire            n27409;
wire      [7:0] n2741;
wire      [7:0] n27410;
wire            n27411;
wire            n27412;
wire            n27413;
wire            n27414;
wire            n27415;
wire      [7:0] n27416;
wire            n27417;
wire            n27418;
wire            n27419;
wire      [7:0] n2742;
wire            n27420;
wire            n27421;
wire      [7:0] n27422;
wire            n27423;
wire            n27424;
wire            n27425;
wire            n27426;
wire            n27427;
wire      [7:0] n27428;
wire            n27429;
wire      [7:0] n2743;
wire            n27430;
wire            n27431;
wire            n27432;
wire            n27433;
wire      [7:0] n27434;
wire            n27435;
wire            n27436;
wire            n27437;
wire            n27438;
wire            n27439;
wire      [7:0] n2744;
wire      [7:0] n27440;
wire            n27441;
wire            n27442;
wire            n27443;
wire            n27444;
wire            n27445;
wire      [7:0] n27446;
wire            n27447;
wire            n27448;
wire            n27449;
wire      [7:0] n2745;
wire            n27450;
wire            n27451;
wire      [7:0] n27452;
wire            n27453;
wire            n27454;
wire            n27455;
wire            n27456;
wire            n27457;
wire      [7:0] n27458;
wire            n27459;
wire      [7:0] n2746;
wire            n27460;
wire            n27461;
wire            n27462;
wire            n27463;
wire      [7:0] n27464;
wire            n27465;
wire            n27466;
wire            n27467;
wire            n27468;
wire            n27469;
wire      [7:0] n2747;
wire      [7:0] n27470;
wire            n27471;
wire            n27472;
wire            n27473;
wire            n27474;
wire            n27475;
wire      [7:0] n27476;
wire            n27477;
wire            n27478;
wire            n27479;
wire      [7:0] n2748;
wire            n27480;
wire            n27481;
wire      [7:0] n27482;
wire            n27483;
wire            n27484;
wire            n27485;
wire            n27486;
wire            n27487;
wire      [7:0] n27488;
wire            n27489;
wire      [7:0] n2749;
wire            n27490;
wire            n27491;
wire            n27492;
wire            n27493;
wire      [7:0] n27494;
wire            n27495;
wire            n27496;
wire            n27497;
wire            n27498;
wire            n27499;
wire      [7:0] n2750;
wire      [7:0] n27500;
wire            n27501;
wire            n27502;
wire            n27503;
wire            n27504;
wire            n27505;
wire      [7:0] n27506;
wire            n27507;
wire            n27508;
wire            n27509;
wire      [7:0] n2751;
wire            n27510;
wire            n27511;
wire      [7:0] n27512;
wire            n27513;
wire            n27514;
wire            n27515;
wire            n27516;
wire            n27517;
wire      [7:0] n27518;
wire            n27519;
wire      [7:0] n2752;
wire            n27520;
wire            n27521;
wire            n27522;
wire            n27523;
wire      [7:0] n27524;
wire            n27525;
wire            n27526;
wire            n27527;
wire            n27528;
wire            n27529;
wire      [7:0] n2753;
wire      [7:0] n27530;
wire            n27531;
wire            n27532;
wire            n27533;
wire            n27534;
wire            n27535;
wire      [7:0] n27536;
wire            n27537;
wire            n27538;
wire            n27539;
wire      [7:0] n2754;
wire            n27540;
wire            n27541;
wire      [7:0] n27542;
wire            n27543;
wire            n27544;
wire            n27545;
wire            n27546;
wire            n27547;
wire      [7:0] n27548;
wire            n27549;
wire      [7:0] n2755;
wire            n27550;
wire            n27551;
wire            n27552;
wire            n27553;
wire      [7:0] n27554;
wire            n27555;
wire            n27556;
wire            n27557;
wire            n27558;
wire            n27559;
wire      [7:0] n2756;
wire      [7:0] n27560;
wire            n27561;
wire            n27562;
wire            n27563;
wire            n27564;
wire            n27565;
wire      [7:0] n27566;
wire            n27567;
wire            n27568;
wire            n27569;
wire      [7:0] n2757;
wire            n27570;
wire            n27571;
wire      [7:0] n27572;
wire            n27573;
wire            n27574;
wire            n27575;
wire            n27576;
wire            n27577;
wire      [7:0] n27578;
wire            n27579;
wire      [7:0] n2758;
wire            n27580;
wire            n27581;
wire            n27582;
wire            n27583;
wire      [7:0] n27584;
wire            n27585;
wire            n27586;
wire            n27587;
wire            n27588;
wire            n27589;
wire      [7:0] n2759;
wire      [7:0] n27590;
wire            n27591;
wire            n27592;
wire            n27593;
wire            n27594;
wire            n27595;
wire      [7:0] n27596;
wire            n27597;
wire            n27598;
wire            n27599;
wire            n276;
wire      [7:0] n2760;
wire            n27600;
wire            n27601;
wire      [7:0] n27602;
wire            n27603;
wire            n27604;
wire            n27605;
wire            n27606;
wire            n27607;
wire      [7:0] n27608;
wire            n27609;
wire      [7:0] n2761;
wire            n27610;
wire            n27611;
wire            n27612;
wire            n27613;
wire      [7:0] n27614;
wire            n27615;
wire            n27616;
wire            n27617;
wire            n27618;
wire            n27619;
wire      [7:0] n2762;
wire      [7:0] n27620;
wire            n27621;
wire            n27622;
wire            n27623;
wire            n27624;
wire            n27625;
wire      [7:0] n27626;
wire            n27627;
wire            n27628;
wire            n27629;
wire      [7:0] n2763;
wire            n27630;
wire            n27631;
wire      [7:0] n27632;
wire            n27633;
wire            n27634;
wire            n27635;
wire            n27636;
wire            n27637;
wire      [7:0] n27638;
wire            n27639;
wire      [7:0] n2764;
wire            n27640;
wire            n27641;
wire            n27642;
wire            n27643;
wire      [7:0] n27644;
wire            n27645;
wire            n27646;
wire            n27647;
wire            n27648;
wire            n27649;
wire      [7:0] n2765;
wire      [7:0] n27650;
wire            n27651;
wire            n27652;
wire            n27653;
wire            n27654;
wire            n27655;
wire      [7:0] n27656;
wire            n27657;
wire            n27658;
wire            n27659;
wire      [7:0] n2766;
wire            n27660;
wire            n27661;
wire      [7:0] n27662;
wire            n27663;
wire            n27664;
wire            n27665;
wire            n27666;
wire            n27667;
wire      [7:0] n27668;
wire            n27669;
wire      [7:0] n2767;
wire            n27670;
wire            n27671;
wire            n27672;
wire            n27673;
wire      [7:0] n27674;
wire            n27675;
wire            n27676;
wire            n27677;
wire            n27678;
wire            n27679;
wire      [7:0] n2768;
wire      [7:0] n27680;
wire            n27681;
wire            n27682;
wire            n27683;
wire            n27684;
wire            n27685;
wire      [7:0] n27686;
wire            n27687;
wire            n27688;
wire            n27689;
wire      [7:0] n2769;
wire            n27690;
wire            n27691;
wire      [7:0] n27692;
wire            n27693;
wire            n27694;
wire            n27695;
wire            n27696;
wire            n27697;
wire      [7:0] n27698;
wire            n27699;
wire      [7:0] n2770;
wire            n27700;
wire            n27701;
wire            n27702;
wire            n27703;
wire      [7:0] n27704;
wire            n27705;
wire            n27706;
wire            n27707;
wire            n27708;
wire            n27709;
wire      [7:0] n2771;
wire      [7:0] n27710;
wire            n27711;
wire            n27712;
wire            n27713;
wire            n27714;
wire            n27715;
wire      [7:0] n27716;
wire            n27717;
wire            n27718;
wire            n27719;
wire      [7:0] n2772;
wire            n27720;
wire            n27721;
wire      [7:0] n27722;
wire            n27723;
wire            n27724;
wire            n27725;
wire            n27726;
wire            n27727;
wire      [7:0] n27728;
wire            n27729;
wire      [7:0] n2773;
wire            n27730;
wire            n27731;
wire            n27732;
wire            n27733;
wire      [7:0] n27734;
wire            n27735;
wire            n27736;
wire            n27737;
wire            n27738;
wire            n27739;
wire      [7:0] n2774;
wire      [7:0] n27740;
wire            n27741;
wire            n27742;
wire            n27743;
wire            n27744;
wire            n27745;
wire      [7:0] n27746;
wire            n27747;
wire            n27748;
wire            n27749;
wire      [7:0] n2775;
wire            n27750;
wire            n27751;
wire      [7:0] n27752;
wire            n27753;
wire            n27754;
wire            n27755;
wire            n27756;
wire            n27757;
wire      [7:0] n27758;
wire            n27759;
wire      [7:0] n2776;
wire            n27760;
wire            n27761;
wire            n27762;
wire            n27763;
wire      [7:0] n27764;
wire            n27765;
wire            n27766;
wire            n27767;
wire            n27768;
wire            n27769;
wire      [7:0] n2777;
wire      [7:0] n27770;
wire            n27771;
wire            n27772;
wire            n27773;
wire            n27774;
wire            n27775;
wire      [7:0] n27776;
wire            n27777;
wire            n27778;
wire            n27779;
wire      [7:0] n2778;
wire            n27780;
wire            n27781;
wire      [7:0] n27782;
wire            n27783;
wire            n27784;
wire            n27785;
wire            n27786;
wire            n27787;
wire      [7:0] n27788;
wire            n27789;
wire      [7:0] n2779;
wire            n27790;
wire            n27791;
wire            n27792;
wire            n27793;
wire      [7:0] n27794;
wire            n27795;
wire            n27796;
wire            n27797;
wire            n27798;
wire            n27799;
wire            n278;
wire      [7:0] n2780;
wire      [7:0] n27800;
wire            n27801;
wire            n27802;
wire            n27803;
wire            n27804;
wire            n27805;
wire      [7:0] n27806;
wire            n27807;
wire            n27808;
wire            n27809;
wire      [7:0] n2781;
wire            n27810;
wire            n27811;
wire      [7:0] n27812;
wire            n27813;
wire            n27814;
wire            n27815;
wire            n27816;
wire            n27817;
wire      [7:0] n27818;
wire            n27819;
wire      [7:0] n2782;
wire            n27820;
wire            n27821;
wire            n27822;
wire            n27823;
wire      [7:0] n27824;
wire            n27825;
wire            n27826;
wire            n27827;
wire            n27828;
wire            n27829;
wire      [7:0] n2783;
wire      [7:0] n27830;
wire            n27831;
wire            n27832;
wire            n27833;
wire            n27834;
wire            n27835;
wire      [7:0] n27836;
wire            n27837;
wire            n27838;
wire            n27839;
wire      [7:0] n2784;
wire            n27840;
wire            n27841;
wire      [7:0] n27842;
wire            n27843;
wire            n27844;
wire            n27845;
wire            n27846;
wire            n27847;
wire      [7:0] n27848;
wire            n27849;
wire      [7:0] n2785;
wire            n27850;
wire            n27851;
wire            n27852;
wire            n27853;
wire      [7:0] n27854;
wire            n27855;
wire            n27856;
wire            n27857;
wire            n27858;
wire            n27859;
wire      [7:0] n2786;
wire      [7:0] n27860;
wire            n27861;
wire            n27862;
wire            n27863;
wire            n27864;
wire            n27865;
wire      [7:0] n27866;
wire            n27867;
wire            n27868;
wire            n27869;
wire      [7:0] n2787;
wire            n27870;
wire            n27871;
wire      [7:0] n27872;
wire            n27873;
wire            n27874;
wire            n27875;
wire            n27876;
wire            n27877;
wire      [7:0] n27878;
wire            n27879;
wire      [7:0] n2788;
wire            n27880;
wire            n27881;
wire            n27882;
wire            n27883;
wire      [7:0] n27884;
wire            n27885;
wire            n27886;
wire            n27887;
wire            n27888;
wire            n27889;
wire      [7:0] n2789;
wire      [7:0] n27890;
wire            n27891;
wire            n27892;
wire            n27893;
wire            n27894;
wire            n27895;
wire      [7:0] n27896;
wire            n27897;
wire            n27898;
wire            n27899;
wire      [7:0] n2790;
wire            n27900;
wire            n27901;
wire      [7:0] n27902;
wire            n27903;
wire            n27904;
wire            n27905;
wire            n27906;
wire            n27907;
wire      [7:0] n27908;
wire            n27909;
wire      [7:0] n2791;
wire            n27910;
wire            n27911;
wire            n27912;
wire            n27913;
wire      [7:0] n27914;
wire            n27915;
wire            n27916;
wire            n27917;
wire            n27918;
wire            n27919;
wire      [7:0] n2792;
wire      [7:0] n27920;
wire            n27921;
wire            n27922;
wire            n27923;
wire            n27924;
wire            n27925;
wire      [7:0] n27926;
wire            n27927;
wire            n27928;
wire            n27929;
wire      [7:0] n2793;
wire            n27930;
wire            n27931;
wire      [7:0] n27932;
wire            n27933;
wire            n27934;
wire            n27935;
wire            n27936;
wire            n27937;
wire      [7:0] n27938;
wire            n27939;
wire      [7:0] n2794;
wire            n27940;
wire            n27941;
wire            n27942;
wire            n27943;
wire      [7:0] n27944;
wire            n27945;
wire            n27946;
wire            n27947;
wire            n27948;
wire            n27949;
wire      [7:0] n2795;
wire      [7:0] n27950;
wire            n27951;
wire            n27952;
wire            n27953;
wire            n27954;
wire            n27955;
wire      [7:0] n27956;
wire            n27957;
wire            n27958;
wire            n27959;
wire      [7:0] n2796;
wire            n27960;
wire            n27961;
wire      [7:0] n27962;
wire            n27963;
wire            n27964;
wire            n27965;
wire            n27966;
wire            n27967;
wire      [7:0] n27968;
wire            n27969;
wire      [7:0] n2797;
wire            n27970;
wire            n27971;
wire            n27972;
wire            n27973;
wire      [7:0] n27974;
wire            n27975;
wire            n27976;
wire            n27977;
wire            n27978;
wire            n27979;
wire      [7:0] n2798;
wire      [7:0] n27980;
wire            n27981;
wire            n27982;
wire            n27983;
wire            n27984;
wire            n27985;
wire      [7:0] n27986;
wire            n27987;
wire            n27988;
wire            n27989;
wire      [7:0] n2799;
wire            n27990;
wire            n27991;
wire      [7:0] n27992;
wire            n27993;
wire            n27994;
wire            n27995;
wire            n27996;
wire            n27997;
wire      [7:0] n27998;
wire            n27999;
wire            n280;
wire      [7:0] n2800;
wire            n28000;
wire            n28001;
wire            n28002;
wire            n28003;
wire      [7:0] n28004;
wire            n28005;
wire            n28006;
wire            n28007;
wire            n28008;
wire            n28009;
wire      [7:0] n2801;
wire      [7:0] n28010;
wire            n28011;
wire            n28012;
wire            n28013;
wire            n28014;
wire            n28015;
wire      [7:0] n28016;
wire            n28017;
wire            n28018;
wire            n28019;
wire      [7:0] n2802;
wire            n28020;
wire            n28021;
wire      [7:0] n28022;
wire            n28023;
wire            n28024;
wire            n28025;
wire            n28026;
wire            n28027;
wire      [7:0] n28028;
wire            n28029;
wire      [7:0] n2803;
wire            n28030;
wire            n28031;
wire            n28032;
wire            n28033;
wire      [7:0] n28034;
wire            n28035;
wire            n28036;
wire            n28037;
wire            n28038;
wire            n28039;
wire      [7:0] n2804;
wire      [7:0] n28040;
wire            n28041;
wire            n28042;
wire            n28043;
wire            n28044;
wire            n28045;
wire      [7:0] n28046;
wire            n28047;
wire            n28048;
wire            n28049;
wire      [7:0] n2805;
wire            n28050;
wire            n28051;
wire      [7:0] n28052;
wire            n28053;
wire            n28054;
wire            n28055;
wire            n28056;
wire            n28057;
wire      [7:0] n28058;
wire            n28059;
wire      [7:0] n2806;
wire            n28060;
wire            n28061;
wire            n28062;
wire            n28063;
wire      [7:0] n28064;
wire            n28065;
wire            n28066;
wire            n28067;
wire            n28068;
wire            n28069;
wire      [7:0] n2807;
wire      [7:0] n28070;
wire            n28071;
wire            n28072;
wire            n28073;
wire            n28074;
wire            n28075;
wire      [7:0] n28076;
wire            n28077;
wire            n28078;
wire            n28079;
wire      [7:0] n2808;
wire            n28080;
wire            n28081;
wire      [7:0] n28082;
wire            n28083;
wire            n28084;
wire            n28085;
wire            n28086;
wire            n28087;
wire      [7:0] n28088;
wire            n28089;
wire      [7:0] n2809;
wire            n28090;
wire            n28091;
wire            n28092;
wire            n28093;
wire      [7:0] n28094;
wire            n28095;
wire            n28096;
wire            n28097;
wire            n28098;
wire            n28099;
wire      [7:0] n2810;
wire      [7:0] n28100;
wire            n28101;
wire            n28102;
wire            n28103;
wire            n28104;
wire            n28105;
wire      [7:0] n28106;
wire            n28107;
wire            n28108;
wire            n28109;
wire      [7:0] n2811;
wire            n28110;
wire            n28111;
wire      [7:0] n28112;
wire            n28113;
wire            n28114;
wire            n28115;
wire            n28116;
wire            n28117;
wire      [7:0] n28118;
wire            n28119;
wire      [7:0] n2812;
wire            n28120;
wire            n28121;
wire            n28122;
wire            n28123;
wire      [7:0] n28124;
wire            n28125;
wire            n28126;
wire            n28127;
wire            n28128;
wire            n28129;
wire      [7:0] n2813;
wire      [7:0] n28130;
wire            n28131;
wire            n28132;
wire            n28133;
wire            n28134;
wire            n28135;
wire      [7:0] n28136;
wire            n28137;
wire            n28138;
wire            n28139;
wire      [7:0] n2814;
wire            n28140;
wire            n28141;
wire      [7:0] n28142;
wire            n28143;
wire            n28144;
wire            n28145;
wire            n28146;
wire            n28147;
wire      [7:0] n28148;
wire            n28149;
wire      [7:0] n2815;
wire            n28150;
wire            n28151;
wire            n28152;
wire            n28153;
wire      [7:0] n28154;
wire            n28155;
wire            n28156;
wire            n28157;
wire            n28158;
wire            n28159;
wire      [7:0] n2816;
wire      [7:0] n28160;
wire            n28161;
wire            n28162;
wire            n28163;
wire            n28164;
wire            n28165;
wire      [7:0] n28166;
wire            n28167;
wire            n28168;
wire            n28169;
wire      [7:0] n2817;
wire            n28170;
wire            n28171;
wire      [7:0] n28172;
wire            n28173;
wire            n28174;
wire            n28175;
wire            n28176;
wire            n28177;
wire      [7:0] n28178;
wire            n28179;
wire      [7:0] n2818;
wire            n28180;
wire            n28181;
wire            n28182;
wire            n28183;
wire      [7:0] n28184;
wire            n28185;
wire            n28186;
wire            n28187;
wire            n28188;
wire            n28189;
wire      [7:0] n2819;
wire      [7:0] n28190;
wire            n28191;
wire            n28192;
wire            n28193;
wire            n28194;
wire            n28195;
wire      [7:0] n28196;
wire            n28197;
wire            n28198;
wire            n28199;
wire            n282;
wire      [7:0] n2820;
wire            n28200;
wire            n28201;
wire      [7:0] n28202;
wire            n28203;
wire            n28204;
wire            n28205;
wire            n28206;
wire            n28207;
wire      [7:0] n28208;
wire            n28209;
wire      [7:0] n2821;
wire            n28210;
wire            n28211;
wire            n28212;
wire            n28213;
wire      [7:0] n28214;
wire            n28215;
wire            n28216;
wire            n28217;
wire            n28218;
wire            n28219;
wire      [7:0] n2822;
wire      [7:0] n28220;
wire            n28221;
wire            n28222;
wire            n28223;
wire            n28224;
wire            n28225;
wire      [7:0] n28226;
wire            n28227;
wire            n28228;
wire            n28229;
wire      [7:0] n2823;
wire            n28230;
wire            n28231;
wire      [7:0] n28232;
wire            n28233;
wire            n28234;
wire            n28235;
wire            n28236;
wire            n28237;
wire      [7:0] n28238;
wire            n28239;
wire      [7:0] n2824;
wire            n28240;
wire            n28241;
wire            n28242;
wire            n28243;
wire      [7:0] n28244;
wire            n28245;
wire            n28246;
wire            n28247;
wire            n28248;
wire            n28249;
wire      [7:0] n2825;
wire      [7:0] n28250;
wire            n28251;
wire            n28252;
wire            n28253;
wire            n28254;
wire            n28255;
wire      [7:0] n28256;
wire            n28257;
wire            n28258;
wire            n28259;
wire      [7:0] n2826;
wire            n28260;
wire            n28261;
wire      [7:0] n28262;
wire            n28263;
wire            n28264;
wire            n28265;
wire            n28266;
wire            n28267;
wire      [7:0] n28268;
wire            n28269;
wire      [7:0] n2827;
wire            n28270;
wire            n28271;
wire            n28272;
wire            n28273;
wire      [7:0] n28274;
wire            n28275;
wire            n28276;
wire            n28277;
wire            n28278;
wire            n28279;
wire      [7:0] n2828;
wire      [7:0] n28280;
wire            n28281;
wire            n28282;
wire            n28283;
wire            n28284;
wire            n28285;
wire      [7:0] n28286;
wire            n28287;
wire            n28288;
wire            n28289;
wire      [7:0] n2829;
wire            n28290;
wire            n28291;
wire      [7:0] n28292;
wire            n28293;
wire            n28294;
wire            n28295;
wire            n28296;
wire            n28297;
wire      [7:0] n28298;
wire            n28299;
wire      [7:0] n2830;
wire            n28300;
wire            n28301;
wire            n28302;
wire            n28303;
wire      [7:0] n28304;
wire            n28305;
wire            n28306;
wire            n28307;
wire            n28308;
wire            n28309;
wire      [7:0] n2831;
wire      [7:0] n28310;
wire            n28311;
wire            n28312;
wire            n28313;
wire            n28314;
wire            n28315;
wire      [7:0] n28316;
wire            n28317;
wire            n28318;
wire            n28319;
wire      [7:0] n2832;
wire            n28320;
wire            n28321;
wire      [7:0] n28322;
wire            n28323;
wire            n28324;
wire            n28325;
wire            n28326;
wire            n28327;
wire      [7:0] n28328;
wire            n28329;
wire      [7:0] n2833;
wire            n28330;
wire            n28331;
wire            n28332;
wire            n28333;
wire      [7:0] n28334;
wire            n28335;
wire            n28336;
wire            n28337;
wire            n28338;
wire            n28339;
wire      [7:0] n2834;
wire      [7:0] n28340;
wire            n28341;
wire            n28342;
wire            n28343;
wire            n28344;
wire            n28345;
wire      [7:0] n28346;
wire            n28347;
wire            n28348;
wire            n28349;
wire      [7:0] n2835;
wire            n28350;
wire            n28351;
wire      [7:0] n28352;
wire            n28353;
wire            n28354;
wire            n28355;
wire            n28356;
wire            n28357;
wire      [7:0] n28358;
wire            n28359;
wire      [7:0] n2836;
wire            n28360;
wire            n28361;
wire            n28362;
wire            n28363;
wire      [7:0] n28364;
wire            n28365;
wire            n28366;
wire            n28367;
wire            n28368;
wire            n28369;
wire      [7:0] n2837;
wire      [7:0] n28370;
wire            n28371;
wire            n28372;
wire            n28373;
wire            n28374;
wire            n28375;
wire      [7:0] n28376;
wire            n28377;
wire            n28378;
wire            n28379;
wire      [7:0] n2838;
wire            n28380;
wire            n28381;
wire      [7:0] n28382;
wire            n28383;
wire            n28384;
wire            n28385;
wire            n28386;
wire            n28387;
wire      [7:0] n28388;
wire            n28389;
wire      [7:0] n2839;
wire            n28390;
wire            n28391;
wire            n28392;
wire            n28393;
wire      [7:0] n28394;
wire            n28395;
wire            n28396;
wire            n28397;
wire            n28398;
wire            n28399;
wire            n284;
wire      [7:0] n2840;
wire      [7:0] n28400;
wire            n28401;
wire            n28402;
wire            n28403;
wire            n28404;
wire            n28405;
wire      [7:0] n28406;
wire            n28407;
wire            n28408;
wire            n28409;
wire      [7:0] n2841;
wire            n28410;
wire            n28411;
wire      [7:0] n28412;
wire            n28413;
wire            n28414;
wire            n28415;
wire            n28416;
wire            n28417;
wire      [7:0] n28418;
wire            n28419;
wire      [7:0] n2842;
wire            n28420;
wire            n28421;
wire            n28422;
wire            n28423;
wire      [7:0] n28424;
wire            n28425;
wire            n28426;
wire            n28427;
wire            n28428;
wire            n28429;
wire      [7:0] n2843;
wire      [7:0] n28430;
wire            n28431;
wire            n28432;
wire            n28433;
wire            n28434;
wire            n28435;
wire      [7:0] n28436;
wire            n28437;
wire            n28438;
wire            n28439;
wire      [7:0] n2844;
wire            n28440;
wire            n28441;
wire      [7:0] n28442;
wire            n28443;
wire            n28444;
wire            n28445;
wire            n28446;
wire            n28447;
wire      [7:0] n28448;
wire            n28449;
wire      [7:0] n2845;
wire            n28450;
wire            n28451;
wire            n28452;
wire            n28453;
wire      [7:0] n28454;
wire            n28455;
wire            n28456;
wire            n28457;
wire            n28458;
wire            n28459;
wire      [7:0] n2846;
wire      [7:0] n28460;
wire            n28461;
wire            n28462;
wire            n28463;
wire            n28464;
wire            n28465;
wire      [7:0] n28466;
wire            n28467;
wire            n28468;
wire            n28469;
wire      [7:0] n2847;
wire            n28470;
wire            n28471;
wire      [7:0] n28472;
wire            n28473;
wire            n28474;
wire            n28475;
wire            n28476;
wire            n28477;
wire      [7:0] n28478;
wire            n28479;
wire      [7:0] n2848;
wire            n28480;
wire            n28481;
wire            n28482;
wire            n28483;
wire      [7:0] n28484;
wire            n28485;
wire            n28486;
wire            n28487;
wire            n28488;
wire            n28489;
wire      [7:0] n2849;
wire      [7:0] n28490;
wire            n28491;
wire            n28492;
wire            n28493;
wire            n28494;
wire            n28495;
wire      [7:0] n28496;
wire            n28497;
wire            n28498;
wire            n28499;
wire      [7:0] n2850;
wire            n28500;
wire            n28501;
wire      [7:0] n28502;
wire            n28503;
wire            n28504;
wire            n28505;
wire            n28506;
wire            n28507;
wire      [7:0] n28508;
wire            n28509;
wire      [7:0] n2851;
wire            n28510;
wire            n28511;
wire            n28512;
wire            n28513;
wire      [7:0] n28514;
wire            n28515;
wire            n28516;
wire            n28517;
wire            n28518;
wire            n28519;
wire      [7:0] n2852;
wire      [7:0] n28520;
wire            n28521;
wire            n28522;
wire            n28523;
wire            n28524;
wire            n28525;
wire      [7:0] n28526;
wire            n28527;
wire            n28528;
wire            n28529;
wire      [7:0] n2853;
wire            n28530;
wire            n28531;
wire      [7:0] n28532;
wire            n28533;
wire            n28534;
wire            n28535;
wire            n28536;
wire            n28537;
wire      [7:0] n28538;
wire            n28539;
wire      [7:0] n2854;
wire            n28540;
wire            n28541;
wire            n28542;
wire            n28543;
wire      [7:0] n28544;
wire            n28545;
wire            n28546;
wire            n28547;
wire            n28548;
wire            n28549;
wire      [7:0] n2855;
wire      [7:0] n28550;
wire            n28551;
wire            n28552;
wire            n28553;
wire            n28554;
wire            n28555;
wire      [7:0] n28556;
wire            n28557;
wire            n28558;
wire            n28559;
wire      [7:0] n2856;
wire            n28560;
wire            n28561;
wire      [7:0] n28562;
wire            n28563;
wire            n28564;
wire            n28565;
wire            n28566;
wire            n28567;
wire      [7:0] n28568;
wire            n28569;
wire      [7:0] n2857;
wire            n28570;
wire            n28571;
wire            n28572;
wire            n28573;
wire      [7:0] n28574;
wire            n28575;
wire            n28576;
wire            n28577;
wire            n28578;
wire            n28579;
wire      [7:0] n2858;
wire      [7:0] n28580;
wire            n28581;
wire            n28582;
wire            n28583;
wire            n28584;
wire            n28585;
wire      [7:0] n28586;
wire            n28587;
wire            n28588;
wire            n28589;
wire      [7:0] n2859;
wire            n28590;
wire            n28591;
wire      [7:0] n28592;
wire            n28593;
wire            n28594;
wire            n28595;
wire            n28596;
wire            n28597;
wire      [7:0] n28598;
wire            n28599;
wire            n286;
wire      [7:0] n2860;
wire            n28600;
wire            n28601;
wire            n28602;
wire            n28603;
wire      [7:0] n28604;
wire            n28605;
wire            n28606;
wire            n28607;
wire            n28608;
wire            n28609;
wire      [7:0] n2861;
wire      [7:0] n28610;
wire            n28611;
wire            n28612;
wire            n28613;
wire            n28614;
wire            n28615;
wire      [7:0] n28616;
wire            n28617;
wire            n28618;
wire            n28619;
wire      [7:0] n2862;
wire            n28620;
wire            n28621;
wire      [7:0] n28622;
wire            n28623;
wire            n28624;
wire            n28625;
wire            n28626;
wire            n28627;
wire      [7:0] n28628;
wire            n28629;
wire      [7:0] n2863;
wire            n28630;
wire            n28631;
wire            n28632;
wire            n28633;
wire      [7:0] n28634;
wire            n28635;
wire            n28636;
wire            n28637;
wire            n28638;
wire            n28639;
wire      [7:0] n2864;
wire      [7:0] n28640;
wire            n28641;
wire            n28642;
wire            n28643;
wire            n28644;
wire            n28645;
wire      [7:0] n28646;
wire            n28647;
wire            n28648;
wire            n28649;
wire      [7:0] n2865;
wire            n28650;
wire            n28651;
wire      [7:0] n28652;
wire            n28653;
wire            n28654;
wire            n28655;
wire            n28656;
wire            n28657;
wire      [7:0] n28658;
wire            n28659;
wire      [7:0] n2866;
wire            n28660;
wire            n28661;
wire            n28662;
wire            n28663;
wire      [7:0] n28664;
wire            n28665;
wire            n28666;
wire            n28667;
wire            n28668;
wire            n28669;
wire      [7:0] n2867;
wire      [7:0] n28670;
wire            n28671;
wire            n28672;
wire            n28673;
wire            n28674;
wire            n28675;
wire      [7:0] n28676;
wire            n28677;
wire            n28678;
wire            n28679;
wire      [7:0] n2868;
wire            n28680;
wire            n28681;
wire      [7:0] n28682;
wire            n28683;
wire            n28684;
wire            n28685;
wire            n28686;
wire            n28687;
wire      [7:0] n28688;
wire            n28689;
wire      [7:0] n2869;
wire            n28690;
wire            n28691;
wire            n28692;
wire            n28693;
wire      [7:0] n28694;
wire            n28695;
wire            n28696;
wire            n28697;
wire            n28698;
wire            n28699;
wire      [7:0] n2870;
wire      [7:0] n28700;
wire            n28701;
wire            n28702;
wire            n28703;
wire            n28704;
wire            n28705;
wire      [7:0] n28706;
wire            n28707;
wire            n28708;
wire            n28709;
wire      [7:0] n2871;
wire            n28710;
wire            n28711;
wire      [7:0] n28712;
wire            n28713;
wire            n28714;
wire            n28715;
wire            n28716;
wire            n28717;
wire      [7:0] n28718;
wire            n28719;
wire      [7:0] n2872;
wire            n28720;
wire            n28721;
wire            n28722;
wire            n28723;
wire      [7:0] n28724;
wire            n28725;
wire            n28726;
wire            n28727;
wire            n28728;
wire            n28729;
wire      [7:0] n2873;
wire      [7:0] n28730;
wire            n28731;
wire            n28732;
wire            n28733;
wire            n28734;
wire            n28735;
wire      [7:0] n28736;
wire            n28737;
wire            n28738;
wire            n28739;
wire      [7:0] n2874;
wire            n28740;
wire            n28741;
wire      [7:0] n28742;
wire            n28743;
wire            n28744;
wire            n28745;
wire            n28746;
wire            n28747;
wire      [7:0] n28748;
wire            n28749;
wire      [7:0] n2875;
wire            n28750;
wire            n28751;
wire            n28752;
wire            n28753;
wire      [7:0] n28754;
wire            n28755;
wire            n28756;
wire            n28757;
wire            n28758;
wire            n28759;
wire      [7:0] n2876;
wire      [7:0] n28760;
wire            n28761;
wire            n28762;
wire            n28763;
wire            n28764;
wire            n28765;
wire      [7:0] n28766;
wire            n28767;
wire            n28768;
wire            n28769;
wire      [7:0] n2877;
wire            n28770;
wire            n28771;
wire      [7:0] n28772;
wire            n28773;
wire            n28774;
wire            n28775;
wire            n28776;
wire            n28777;
wire      [7:0] n28778;
wire            n28779;
wire      [7:0] n2878;
wire            n28780;
wire            n28781;
wire            n28782;
wire            n28783;
wire      [7:0] n28784;
wire            n28785;
wire            n28786;
wire            n28787;
wire            n28788;
wire            n28789;
wire      [7:0] n2879;
wire      [7:0] n28790;
wire            n28791;
wire            n28792;
wire            n28793;
wire            n28794;
wire            n28795;
wire      [7:0] n28796;
wire            n28797;
wire            n28798;
wire            n28799;
wire            n288;
wire      [7:0] n2880;
wire            n28800;
wire            n28801;
wire      [7:0] n28802;
wire            n28803;
wire            n28804;
wire            n28805;
wire            n28806;
wire            n28807;
wire      [7:0] n28808;
wire            n28809;
wire      [7:0] n2881;
wire            n28810;
wire            n28811;
wire            n28812;
wire            n28813;
wire      [7:0] n28814;
wire            n28815;
wire            n28816;
wire            n28817;
wire            n28818;
wire            n28819;
wire      [7:0] n2882;
wire      [7:0] n28820;
wire            n28821;
wire            n28822;
wire            n28823;
wire            n28824;
wire            n28825;
wire      [7:0] n28826;
wire            n28827;
wire            n28828;
wire            n28829;
wire      [7:0] n2883;
wire            n28830;
wire            n28831;
wire      [7:0] n28832;
wire            n28833;
wire            n28834;
wire            n28835;
wire            n28836;
wire            n28837;
wire      [7:0] n28838;
wire            n28839;
wire      [7:0] n2884;
wire            n28840;
wire            n28841;
wire            n28842;
wire            n28843;
wire      [7:0] n28844;
wire            n28845;
wire            n28846;
wire            n28847;
wire            n28848;
wire            n28849;
wire      [7:0] n2885;
wire      [7:0] n28850;
wire            n28851;
wire            n28852;
wire            n28853;
wire            n28854;
wire            n28855;
wire      [7:0] n28856;
wire            n28857;
wire            n28858;
wire            n28859;
wire      [7:0] n2886;
wire            n28860;
wire            n28861;
wire      [7:0] n28862;
wire            n28863;
wire            n28864;
wire            n28865;
wire            n28866;
wire            n28867;
wire      [7:0] n28868;
wire            n28869;
wire      [7:0] n2887;
wire            n28870;
wire            n28871;
wire            n28872;
wire            n28873;
wire      [7:0] n28874;
wire            n28875;
wire            n28876;
wire            n28877;
wire            n28878;
wire            n28879;
wire      [7:0] n2888;
wire      [7:0] n28880;
wire            n28881;
wire            n28882;
wire            n28883;
wire            n28884;
wire            n28885;
wire      [7:0] n28886;
wire            n28887;
wire            n28888;
wire            n28889;
wire      [7:0] n2889;
wire            n28890;
wire            n28891;
wire      [7:0] n28892;
wire            n28893;
wire            n28894;
wire            n28895;
wire            n28896;
wire            n28897;
wire      [7:0] n28898;
wire            n28899;
wire      [7:0] n2890;
wire            n28900;
wire            n28901;
wire            n28902;
wire            n28903;
wire      [7:0] n28904;
wire            n28905;
wire            n28906;
wire            n28907;
wire            n28908;
wire            n28909;
wire      [7:0] n2891;
wire      [7:0] n28910;
wire            n28911;
wire            n28912;
wire            n28913;
wire            n28914;
wire            n28915;
wire      [7:0] n28916;
wire            n28917;
wire            n28918;
wire            n28919;
wire      [7:0] n2892;
wire            n28920;
wire            n28921;
wire      [7:0] n28922;
wire            n28923;
wire            n28924;
wire            n28925;
wire            n28926;
wire            n28927;
wire      [7:0] n28928;
wire            n28929;
wire      [7:0] n2893;
wire            n28930;
wire            n28931;
wire            n28932;
wire            n28933;
wire      [7:0] n28934;
wire            n28935;
wire            n28936;
wire            n28937;
wire            n28938;
wire            n28939;
wire      [7:0] n2894;
wire      [7:0] n28940;
wire            n28941;
wire            n28942;
wire            n28943;
wire            n28944;
wire            n28945;
wire      [7:0] n28946;
wire            n28947;
wire            n28948;
wire            n28949;
wire      [7:0] n2895;
wire            n28950;
wire            n28951;
wire      [7:0] n28952;
wire            n28953;
wire            n28954;
wire            n28955;
wire            n28956;
wire            n28957;
wire      [7:0] n28958;
wire            n28959;
wire      [7:0] n2896;
wire            n28960;
wire            n28961;
wire            n28962;
wire            n28963;
wire      [7:0] n28964;
wire            n28965;
wire            n28966;
wire            n28967;
wire            n28968;
wire            n28969;
wire      [7:0] n2897;
wire      [7:0] n28970;
wire            n28971;
wire            n28972;
wire            n28973;
wire            n28974;
wire            n28975;
wire      [7:0] n28976;
wire            n28977;
wire            n28978;
wire            n28979;
wire      [7:0] n2898;
wire            n28980;
wire            n28981;
wire      [7:0] n28982;
wire            n28983;
wire            n28984;
wire            n28985;
wire            n28986;
wire            n28987;
wire      [7:0] n28988;
wire            n28989;
wire      [7:0] n2899;
wire            n28990;
wire            n28991;
wire            n28992;
wire            n28993;
wire      [7:0] n28994;
wire            n28995;
wire            n28996;
wire            n28997;
wire            n28998;
wire            n28999;
wire            n29;
wire            n290;
wire      [7:0] n2900;
wire      [7:0] n29000;
wire            n29001;
wire            n29002;
wire            n29003;
wire            n29004;
wire            n29005;
wire      [7:0] n29006;
wire            n29007;
wire            n29008;
wire            n29009;
wire      [7:0] n2901;
wire            n29010;
wire            n29011;
wire      [7:0] n29012;
wire            n29013;
wire            n29014;
wire            n29015;
wire            n29016;
wire            n29017;
wire      [7:0] n29018;
wire            n29019;
wire      [7:0] n2902;
wire            n29020;
wire            n29021;
wire            n29022;
wire            n29023;
wire      [7:0] n29024;
wire            n29025;
wire            n29026;
wire            n29027;
wire            n29028;
wire            n29029;
wire      [7:0] n2903;
wire      [7:0] n29030;
wire            n29031;
wire            n29032;
wire            n29033;
wire            n29034;
wire            n29035;
wire      [7:0] n29036;
wire            n29037;
wire            n29038;
wire            n29039;
wire      [7:0] n2904;
wire            n29040;
wire            n29041;
wire      [7:0] n29042;
wire            n29043;
wire            n29044;
wire            n29045;
wire            n29046;
wire            n29047;
wire      [7:0] n29048;
wire            n29049;
wire      [7:0] n2905;
wire            n29050;
wire            n29051;
wire            n29052;
wire            n29053;
wire      [7:0] n29054;
wire            n29055;
wire            n29056;
wire            n29057;
wire            n29058;
wire            n29059;
wire      [7:0] n2906;
wire      [7:0] n29060;
wire            n29061;
wire            n29062;
wire            n29063;
wire            n29064;
wire            n29065;
wire      [7:0] n29066;
wire            n29067;
wire            n29068;
wire            n29069;
wire      [7:0] n2907;
wire            n29070;
wire            n29071;
wire      [7:0] n29072;
wire            n29073;
wire            n29074;
wire            n29075;
wire            n29076;
wire            n29077;
wire      [7:0] n29078;
wire            n29079;
wire      [7:0] n2908;
wire            n29080;
wire            n29081;
wire            n29082;
wire            n29083;
wire      [7:0] n29084;
wire            n29085;
wire            n29086;
wire            n29087;
wire            n29088;
wire            n29089;
wire      [7:0] n2909;
wire      [7:0] n29090;
wire            n29091;
wire            n29092;
wire            n29093;
wire            n29094;
wire            n29095;
wire      [7:0] n29096;
wire            n29097;
wire            n29098;
wire            n29099;
wire      [7:0] n2910;
wire            n29100;
wire            n29101;
wire      [7:0] n29102;
wire            n29103;
wire            n29104;
wire            n29105;
wire            n29106;
wire            n29107;
wire      [7:0] n29108;
wire            n29109;
wire      [7:0] n2911;
wire            n29110;
wire            n29111;
wire            n29112;
wire            n29113;
wire      [7:0] n29114;
wire            n29115;
wire            n29116;
wire            n29117;
wire            n29118;
wire            n29119;
wire      [7:0] n2912;
wire      [7:0] n29120;
wire            n29121;
wire            n29122;
wire            n29123;
wire            n29124;
wire            n29125;
wire      [7:0] n29126;
wire            n29127;
wire            n29128;
wire            n29129;
wire      [7:0] n2913;
wire            n29130;
wire            n29131;
wire      [7:0] n29132;
wire            n29133;
wire            n29134;
wire            n29135;
wire            n29136;
wire            n29137;
wire      [7:0] n29138;
wire            n29139;
wire      [7:0] n2914;
wire            n29140;
wire            n29141;
wire            n29142;
wire            n29143;
wire      [7:0] n29144;
wire            n29145;
wire            n29146;
wire            n29147;
wire            n29148;
wire            n29149;
wire      [7:0] n2915;
wire      [7:0] n29150;
wire            n29151;
wire            n29152;
wire            n29153;
wire            n29154;
wire            n29155;
wire      [7:0] n29156;
wire            n29157;
wire            n29158;
wire            n29159;
wire            n2916;
wire            n29160;
wire            n29161;
wire      [7:0] n29162;
wire            n29163;
wire            n29164;
wire            n29165;
wire            n29166;
wire            n29167;
wire      [7:0] n29168;
wire            n29169;
wire            n2917;
wire            n29170;
wire            n29171;
wire            n29172;
wire            n29173;
wire      [7:0] n29174;
wire            n29175;
wire            n29176;
wire            n29177;
wire            n29178;
wire            n29179;
wire      [3:0] n2918;
wire      [7:0] n29180;
wire            n29181;
wire            n29182;
wire            n29183;
wire            n29184;
wire            n29185;
wire      [7:0] n29186;
wire            n29187;
wire            n29188;
wire            n29189;
wire      [4:0] n2919;
wire            n29190;
wire            n29191;
wire      [7:0] n29192;
wire            n29193;
wire            n29194;
wire            n29195;
wire            n29196;
wire            n29197;
wire      [7:0] n29198;
wire            n29199;
wire            n292;
wire      [7:0] n2920;
wire            n29200;
wire            n29201;
wire            n29202;
wire            n29203;
wire      [7:0] n29204;
wire            n29205;
wire            n29206;
wire            n29207;
wire            n29208;
wire            n29209;
wire      [3:0] n2921;
wire      [7:0] n29210;
wire            n29211;
wire            n29212;
wire            n29213;
wire            n29214;
wire            n29215;
wire      [7:0] n29216;
wire            n29217;
wire            n29218;
wire            n29219;
wire      [7:0] n2922;
wire            n29220;
wire            n29221;
wire      [7:0] n29222;
wire            n29223;
wire            n29224;
wire            n29225;
wire            n29226;
wire            n29227;
wire      [7:0] n29228;
wire            n29229;
wire      [7:0] n2923;
wire            n29230;
wire            n29231;
wire            n29232;
wire            n29233;
wire      [7:0] n29234;
wire            n29235;
wire            n29236;
wire            n29237;
wire            n29238;
wire            n29239;
wire      [7:0] n2924;
wire      [7:0] n29240;
wire            n29241;
wire            n29242;
wire            n29243;
wire            n29244;
wire            n29245;
wire      [7:0] n29246;
wire            n29247;
wire            n29248;
wire            n29249;
wire            n2925;
wire            n29250;
wire            n29251;
wire      [7:0] n29252;
wire            n29253;
wire            n29254;
wire            n29255;
wire            n29256;
wire            n29257;
wire      [7:0] n29258;
wire            n29259;
wire      [7:0] n2926;
wire            n29260;
wire            n29261;
wire            n29262;
wire            n29263;
wire      [7:0] n29264;
wire            n29265;
wire            n29266;
wire            n29267;
wire            n29268;
wire            n29269;
wire            n2927;
wire      [7:0] n29270;
wire            n29271;
wire            n29272;
wire            n29273;
wire            n29274;
wire            n29275;
wire      [7:0] n29276;
wire            n29277;
wire            n29278;
wire            n2928;
wire            n29280;
wire            n29281;
wire            n29282;
wire      [7:0] n29283;
wire            n29284;
wire            n29285;
wire            n29286;
wire            n29287;
wire            n29288;
wire      [7:0] n29289;
wire            n2929;
wire            n29290;
wire            n29291;
wire            n29292;
wire            n29293;
wire            n29294;
wire      [7:0] n29295;
wire            n29296;
wire            n29297;
wire            n29298;
wire            n29299;
wire            n2930;
wire            n29300;
wire      [7:0] n29301;
wire            n29302;
wire            n29303;
wire            n29304;
wire            n29305;
wire            n29306;
wire      [7:0] n29307;
wire            n29308;
wire            n29309;
wire            n2931;
wire            n29310;
wire            n29311;
wire            n29312;
wire      [7:0] n29313;
wire            n29314;
wire            n29315;
wire            n29316;
wire            n29317;
wire            n29318;
wire      [7:0] n29319;
wire            n2932;
wire            n29320;
wire            n29321;
wire            n29322;
wire            n29323;
wire            n29324;
wire      [7:0] n29325;
wire            n29326;
wire            n29327;
wire            n29328;
wire            n29329;
wire            n2933;
wire            n29330;
wire      [7:0] n29331;
wire            n29332;
wire            n29333;
wire            n29334;
wire            n29335;
wire            n29336;
wire      [7:0] n29337;
wire            n29338;
wire            n29339;
wire            n2934;
wire            n29340;
wire            n29341;
wire            n29342;
wire      [7:0] n29343;
wire            n29344;
wire            n29345;
wire            n29346;
wire            n29347;
wire            n29348;
wire      [7:0] n29349;
wire            n2935;
wire            n29350;
wire            n29351;
wire            n29352;
wire            n29353;
wire            n29354;
wire      [7:0] n29355;
wire            n29356;
wire            n29357;
wire            n29358;
wire            n29359;
wire            n2936;
wire            n29360;
wire      [7:0] n29361;
wire            n29362;
wire            n29363;
wire            n29364;
wire            n29365;
wire            n29366;
wire      [7:0] n29367;
wire            n2937;
wire            n2938;
wire            n2939;
wire            n294;
wire            n2940;
wire            n2941;
wire            n2942;
wire            n2943;
wire            n2944;
wire            n2945;
wire            n2946;
wire            n2947;
wire            n2948;
wire            n2949;
wire            n2950;
wire            n2951;
wire            n2952;
wire            n2953;
wire            n2954;
wire            n2955;
wire            n2956;
wire            n2957;
wire            n2958;
wire            n2959;
wire            n296;
wire            n2960;
wire            n2961;
wire            n2962;
wire            n2963;
wire            n2964;
wire            n2965;
wire            n2966;
wire            n2967;
wire            n2968;
wire            n2969;
wire            n2970;
wire            n2971;
wire            n2972;
wire            n2973;
wire            n2974;
wire            n2975;
wire            n2976;
wire            n2977;
wire            n2978;
wire            n2979;
wire            n298;
wire            n2980;
wire            n2981;
wire            n2982;
wire            n2983;
wire            n2984;
wire            n2985;
wire            n2986;
wire            n2987;
wire            n2988;
wire            n2989;
wire            n2990;
wire            n2991;
wire            n2992;
wire            n2993;
wire            n2994;
wire            n2995;
wire            n2996;
wire            n2997;
wire            n2998;
wire            n2999;
wire            n3;
wire            n300;
wire            n3000;
wire            n3001;
wire            n3002;
wire            n3003;
wire            n3004;
wire            n3005;
wire            n3006;
wire            n3007;
wire            n3008;
wire            n3009;
wire            n3010;
wire            n3011;
wire            n3012;
wire            n3013;
wire            n3014;
wire            n3015;
wire            n3016;
wire            n3017;
wire            n3018;
wire            n3019;
wire            n302;
wire            n3020;
wire            n3021;
wire            n3022;
wire            n3023;
wire            n3024;
wire            n3025;
wire            n3026;
wire            n3027;
wire            n3028;
wire            n3029;
wire            n3030;
wire            n3031;
wire            n3032;
wire            n3033;
wire            n3034;
wire            n3035;
wire            n3036;
wire            n3037;
wire            n3038;
wire            n3039;
wire            n304;
wire            n3040;
wire            n3041;
wire            n3042;
wire            n3043;
wire            n3044;
wire            n3045;
wire            n3046;
wire            n3047;
wire            n3048;
wire            n3049;
wire            n3050;
wire            n3051;
wire            n3052;
wire            n3053;
wire            n3054;
wire            n3055;
wire            n3056;
wire            n3057;
wire            n3058;
wire            n3059;
wire            n306;
wire            n3060;
wire            n3061;
wire            n3062;
wire            n3063;
wire            n3064;
wire            n3065;
wire            n3066;
wire            n3067;
wire            n3068;
wire            n3069;
wire            n3070;
wire            n3071;
wire            n3072;
wire            n3073;
wire            n3074;
wire            n3075;
wire            n3076;
wire            n3077;
wire            n3078;
wire            n3079;
wire            n308;
wire            n3080;
wire            n3081;
wire            n3082;
wire            n3083;
wire            n3084;
wire            n3085;
wire            n3086;
wire            n3087;
wire            n3088;
wire            n3089;
wire            n3090;
wire            n3091;
wire            n3092;
wire            n3093;
wire            n3094;
wire            n3095;
wire            n3096;
wire            n3097;
wire            n3098;
wire            n3099;
wire            n31;
wire            n310;
wire            n3100;
wire            n3101;
wire            n3102;
wire            n3103;
wire            n3104;
wire            n3105;
wire            n3106;
wire            n3107;
wire            n3108;
wire            n3109;
wire            n3110;
wire            n3111;
wire            n3112;
wire            n3113;
wire            n3114;
wire            n3115;
wire            n3116;
wire            n3117;
wire            n3118;
wire            n3119;
wire            n312;
wire            n3120;
wire            n3121;
wire            n3122;
wire            n3123;
wire            n3124;
wire            n3125;
wire            n3126;
wire            n3127;
wire            n3128;
wire            n3129;
wire            n3130;
wire            n3131;
wire            n3132;
wire            n3133;
wire            n3134;
wire            n3135;
wire            n3136;
wire            n3137;
wire            n3138;
wire            n3139;
wire            n314;
wire            n3140;
wire            n3141;
wire            n3142;
wire            n3143;
wire            n3144;
wire            n3145;
wire            n3146;
wire            n3147;
wire            n3148;
wire            n3149;
wire            n3150;
wire            n3151;
wire            n3152;
wire            n3153;
wire            n3154;
wire            n3155;
wire            n3156;
wire            n3157;
wire            n3158;
wire            n3159;
wire            n316;
wire            n3160;
wire            n3161;
wire            n3162;
wire            n3163;
wire            n3164;
wire            n3165;
wire            n3166;
wire            n3167;
wire            n3168;
wire            n3169;
wire            n3170;
wire            n3171;
wire            n3172;
wire            n3173;
wire            n3174;
wire            n3175;
wire            n3176;
wire            n3177;
wire            n3178;
wire            n3179;
wire            n318;
wire            n3180;
wire            n3181;
wire      [7:0] n3182;
wire      [7:0] n3183;
wire      [7:0] n3184;
wire      [7:0] n3185;
wire      [7:0] n3186;
wire      [7:0] n3187;
wire      [7:0] n3188;
wire      [7:0] n3189;
wire      [7:0] n3190;
wire      [7:0] n3191;
wire      [7:0] n3192;
wire      [7:0] n3193;
wire      [7:0] n3194;
wire      [7:0] n3195;
wire      [7:0] n3196;
wire      [7:0] n3197;
wire      [7:0] n3198;
wire      [7:0] n3199;
wire            n32;
wire            n320;
wire      [7:0] n3200;
wire      [7:0] n3201;
wire      [7:0] n3202;
wire      [7:0] n3203;
wire      [7:0] n3204;
wire      [7:0] n3205;
wire      [7:0] n3206;
wire      [7:0] n3207;
wire      [7:0] n3208;
wire      [7:0] n3209;
wire      [7:0] n3210;
wire      [7:0] n3211;
wire      [7:0] n3212;
wire      [7:0] n3213;
wire      [7:0] n3214;
wire      [7:0] n3215;
wire      [7:0] n3216;
wire      [7:0] n3217;
wire      [7:0] n3218;
wire      [7:0] n3219;
wire            n322;
wire      [7:0] n3220;
wire      [7:0] n3221;
wire      [7:0] n3222;
wire      [7:0] n3223;
wire      [7:0] n3224;
wire      [7:0] n3225;
wire      [7:0] n3226;
wire      [7:0] n3227;
wire      [7:0] n3228;
wire      [7:0] n3229;
wire      [7:0] n3230;
wire      [7:0] n3231;
wire      [7:0] n3232;
wire      [7:0] n3233;
wire      [7:0] n3234;
wire      [7:0] n3235;
wire      [7:0] n3236;
wire      [7:0] n3237;
wire      [7:0] n3238;
wire      [7:0] n3239;
wire            n324;
wire      [7:0] n3240;
wire      [7:0] n3241;
wire      [7:0] n3242;
wire      [7:0] n3243;
wire      [7:0] n3244;
wire      [7:0] n3245;
wire      [7:0] n3246;
wire      [7:0] n3247;
wire      [7:0] n3248;
wire      [7:0] n3249;
wire      [7:0] n3250;
wire      [7:0] n3251;
wire      [7:0] n3252;
wire      [7:0] n3253;
wire      [7:0] n3254;
wire      [7:0] n3255;
wire      [7:0] n3256;
wire      [7:0] n3257;
wire      [7:0] n3258;
wire      [7:0] n3259;
wire            n326;
wire      [7:0] n3260;
wire      [7:0] n3261;
wire      [7:0] n3262;
wire      [7:0] n3263;
wire      [7:0] n3264;
wire      [7:0] n3265;
wire      [7:0] n3266;
wire      [7:0] n3267;
wire      [7:0] n3268;
wire      [7:0] n3269;
wire      [7:0] n3270;
wire      [7:0] n3271;
wire      [7:0] n3272;
wire      [7:0] n3273;
wire      [7:0] n3274;
wire      [7:0] n3275;
wire      [7:0] n3276;
wire      [7:0] n3277;
wire      [7:0] n3278;
wire      [7:0] n3279;
wire            n328;
wire      [7:0] n3280;
wire      [7:0] n3281;
wire      [7:0] n3282;
wire      [7:0] n3283;
wire      [7:0] n3284;
wire      [7:0] n3285;
wire      [7:0] n3286;
wire      [7:0] n3287;
wire      [7:0] n3288;
wire      [7:0] n3289;
wire      [7:0] n3290;
wire      [7:0] n3291;
wire      [7:0] n3292;
wire      [7:0] n3293;
wire      [7:0] n3294;
wire      [7:0] n3295;
wire      [7:0] n3296;
wire      [7:0] n3297;
wire      [7:0] n3298;
wire      [7:0] n3299;
wire            n33;
wire            n330;
wire      [7:0] n3300;
wire      [7:0] n3301;
wire      [7:0] n3302;
wire      [7:0] n3303;
wire      [7:0] n3304;
wire      [7:0] n3305;
wire      [7:0] n3306;
wire      [7:0] n3307;
wire      [7:0] n3308;
wire      [7:0] n3309;
wire      [7:0] n3310;
wire      [7:0] n3311;
wire      [7:0] n3312;
wire      [7:0] n3313;
wire      [7:0] n3314;
wire      [7:0] n3315;
wire      [7:0] n3316;
wire      [7:0] n3317;
wire      [7:0] n3318;
wire      [7:0] n3319;
wire            n332;
wire      [7:0] n3320;
wire      [7:0] n3321;
wire      [7:0] n3322;
wire      [7:0] n3323;
wire      [7:0] n3324;
wire      [7:0] n3325;
wire      [7:0] n3326;
wire      [7:0] n3327;
wire      [7:0] n3328;
wire      [7:0] n3329;
wire      [7:0] n3330;
wire      [7:0] n3331;
wire      [7:0] n3332;
wire      [7:0] n3333;
wire      [7:0] n3334;
wire      [7:0] n3335;
wire      [7:0] n3336;
wire      [7:0] n3337;
wire      [7:0] n3338;
wire      [7:0] n3339;
wire            n334;
wire      [7:0] n3340;
wire      [7:0] n3341;
wire      [7:0] n3342;
wire      [7:0] n3343;
wire      [7:0] n3344;
wire      [7:0] n3345;
wire      [7:0] n3346;
wire      [7:0] n3347;
wire      [7:0] n3348;
wire      [7:0] n3349;
wire      [7:0] n3350;
wire      [7:0] n3351;
wire      [7:0] n3352;
wire      [7:0] n3353;
wire      [7:0] n3354;
wire      [7:0] n3355;
wire      [7:0] n3356;
wire      [7:0] n3357;
wire      [7:0] n3358;
wire      [7:0] n3359;
wire            n336;
wire      [7:0] n3360;
wire      [7:0] n3361;
wire      [7:0] n3362;
wire      [7:0] n3363;
wire      [7:0] n3364;
wire      [7:0] n3365;
wire      [7:0] n3366;
wire      [7:0] n3367;
wire      [7:0] n3368;
wire      [7:0] n3369;
wire      [7:0] n3370;
wire      [7:0] n3371;
wire      [7:0] n3372;
wire      [7:0] n3373;
wire      [7:0] n3374;
wire      [7:0] n3375;
wire      [7:0] n3376;
wire      [7:0] n3377;
wire      [7:0] n3378;
wire      [7:0] n3379;
wire            n338;
wire      [7:0] n3380;
wire      [7:0] n3381;
wire      [7:0] n3382;
wire      [7:0] n3383;
wire      [7:0] n3384;
wire      [7:0] n3385;
wire      [7:0] n3386;
wire      [7:0] n3387;
wire      [7:0] n3388;
wire      [7:0] n3389;
wire      [7:0] n3390;
wire      [7:0] n3391;
wire      [7:0] n3392;
wire      [7:0] n3393;
wire      [7:0] n3394;
wire      [7:0] n3395;
wire      [7:0] n3396;
wire      [7:0] n3397;
wire      [7:0] n3398;
wire      [7:0] n3399;
wire            n340;
wire      [7:0] n3400;
wire      [7:0] n3401;
wire      [7:0] n3402;
wire      [7:0] n3403;
wire      [7:0] n3404;
wire      [7:0] n3405;
wire      [7:0] n3406;
wire      [7:0] n3407;
wire      [7:0] n3408;
wire      [7:0] n3409;
wire      [7:0] n3410;
wire      [7:0] n3411;
wire      [7:0] n3412;
wire      [7:0] n3413;
wire      [7:0] n3414;
wire      [7:0] n3415;
wire      [7:0] n3416;
wire      [7:0] n3417;
wire      [7:0] n3418;
wire      [7:0] n3419;
wire            n342;
wire      [7:0] n3420;
wire      [7:0] n3421;
wire      [7:0] n3422;
wire      [7:0] n3423;
wire      [7:0] n3424;
wire      [7:0] n3425;
wire      [7:0] n3426;
wire      [7:0] n3427;
wire      [7:0] n3428;
wire      [7:0] n3429;
wire      [7:0] n3430;
wire      [7:0] n3431;
wire      [7:0] n3432;
wire      [7:0] n3433;
wire      [7:0] n3434;
wire      [7:0] n3435;
wire      [7:0] n3436;
wire      [7:0] n3437;
wire      [4:0] n3438;
wire      [7:0] n3439;
wire            n344;
wire            n3440;
wire            n3441;
wire            n3442;
wire      [7:0] n3443;
wire            n3444;
wire            n3445;
wire            n3446;
wire            n3447;
wire            n3448;
wire            n3449;
wire            n3450;
wire            n3451;
wire            n3452;
wire            n3453;
wire            n3454;
wire      [7:0] n3455;
wire      [7:0] n3456;
wire      [7:0] n3457;
wire      [7:0] n3458;
wire      [7:0] n3459;
wire            n346;
wire      [7:0] n3460;
wire      [7:0] n3461;
wire      [7:0] n3462;
wire      [7:0] n3463;
wire      [7:0] n3464;
wire      [7:0] n3465;
wire      [7:0] n3466;
wire      [7:0] n3467;
wire      [7:0] n3468;
wire            n3469;
wire            n3470;
wire            n3471;
wire      [7:0] n3472;
wire            n3473;
wire            n3474;
wire            n3475;
wire            n3476;
wire            n3477;
wire            n3478;
wire            n3479;
wire            n348;
wire            n3480;
wire            n3481;
wire      [7:0] n3482;
wire      [7:0] n3483;
wire      [7:0] n3484;
wire      [7:0] n3485;
wire      [7:0] n3486;
wire      [7:0] n3487;
wire      [7:0] n3488;
wire      [7:0] n3489;
wire      [7:0] n3490;
wire      [7:0] n3491;
wire      [7:0] n3492;
wire      [7:0] n3493;
wire      [7:0] n3494;
wire            n3496;
wire            n3497;
wire            n3498;
wire            n35;
wire            n350;
wire      [7:0] n3500;
wire            n3502;
wire            n3503;
wire            n3504;
wire            n3506;
wire            n3507;
wire            n3508;
wire            n3509;
wire            n3510;
wire            n3511;
wire            n3512;
wire            n3513;
wire            n3514;
wire            n3515;
wire            n3516;
wire            n3518;
wire      [7:0] n3519;
wire            n352;
wire            n3521;
wire      [7:0] n3522;
wire      [7:0] n3523;
wire      [7:0] n3524;
wire      [7:0] n3525;
wire      [7:0] n3526;
wire      [7:0] n3527;
wire            n3528;
wire            n3529;
wire            n3530;
wire            n3531;
wire            n3532;
wire            n3533;
wire            n3534;
wire            n3535;
wire            n3536;
wire            n3537;
wire            n3538;
wire            n3539;
wire            n354;
wire            n3540;
wire            n3541;
wire            n3542;
wire            n3543;
wire            n3544;
wire            n3545;
wire            n3546;
wire            n3547;
wire            n3548;
wire            n3549;
wire            n3550;
wire      [4:0] n3551;
wire      [4:0] n3552;
wire            n3553;
wire            n3554;
wire            n3555;
wire      [2:0] n3556;
wire            n3558;
wire            n3559;
wire            n356;
wire            n3560;
wire            n3561;
wire            n3562;
wire            n3563;
wire            n3564;
wire            n3565;
wire      [7:0] n3566;
wire            n3567;
wire      [7:0] n3568;
wire      [7:0] n3569;
wire      [7:0] n3570;
wire      [7:0] n3571;
wire      [7:0] n3572;
wire      [7:0] n3573;
wire            n3574;
wire            n3575;
wire            n3576;
wire            n3577;
wire            n3578;
wire            n3579;
wire            n358;
wire            n3580;
wire            n3581;
wire            n3582;
wire            n3583;
wire            n3584;
wire            n3585;
wire            n3586;
wire            n3587;
wire            n3588;
wire            n3589;
wire            n3590;
wire            n3591;
wire      [7:0] n3592;
wire            n3593;
wire      [7:0] n3594;
wire      [7:0] n3595;
wire      [7:0] n3596;
wire      [7:0] n3597;
wire      [7:0] n3598;
wire      [7:0] n3599;
wire            n36;
wire            n360;
wire            n3600;
wire            n3601;
wire            n3602;
wire            n3603;
wire            n3604;
wire            n3605;
wire            n3606;
wire            n3607;
wire            n3608;
wire            n3609;
wire            n3610;
wire            n3611;
wire            n3612;
wire            n3613;
wire            n3614;
wire            n3615;
wire            n3616;
wire            n3617;
wire            n3618;
wire            n3619;
wire            n362;
wire            n3620;
wire            n3621;
wire            n3622;
wire      [4:0] n3623;
wire      [4:0] n3624;
wire            n3625;
wire            n3626;
wire            n3627;
wire      [2:0] n3628;
wire            n3629;
wire            n3630;
wire            n3631;
wire            n3632;
wire            n3633;
wire            n3634;
wire            n3635;
wire            n3636;
wire      [7:0] n3637;
wire            n3638;
wire      [7:0] n3639;
wire            n364;
wire      [7:0] n3640;
wire      [7:0] n3641;
wire      [7:0] n3642;
wire      [7:0] n3643;
wire      [7:0] n3644;
wire            n3645;
wire      [4:0] n3646;
wire            n3648;
wire            n3649;
wire      [2:0] n3650;
wire            n3651;
wire            n3652;
wire            n3654;
wire            n3655;
wire            n3657;
wire            n3658;
wire            n366;
wire            n3660;
wire            n3661;
wire            n3662;
wire            n3663;
wire            n3665;
wire            n3666;
wire            n3668;
wire            n3669;
wire            n3670;
wire            n3671;
wire            n3672;
wire            n3673;
wire            n3674;
wire            n3675;
wire            n3676;
wire            n3677;
wire            n3678;
wire            n3679;
wire            n368;
wire            n3680;
wire            n3681;
wire            n3682;
wire            n3683;
wire            n3684;
wire            n3685;
wire            n3686;
wire            n3687;
wire            n3688;
wire            n3689;
wire            n3690;
wire            n3691;
wire            n3692;
wire            n3693;
wire            n3694;
wire            n3695;
wire            n3696;
wire            n3697;
wire            n3698;
wire            n3699;
wire            n37;
wire            n370;
wire            n3700;
wire            n3702;
wire            n3703;
wire      [7:0] n3705;
wire            n3706;
wire            n3707;
wire            n3708;
wire            n3709;
wire            n3710;
wire            n3711;
wire            n3712;
wire            n3713;
wire            n3714;
wire            n3715;
wire            n3716;
wire            n3717;
wire            n3718;
wire            n3719;
wire            n372;
wire            n3720;
wire            n3721;
wire            n3722;
wire            n3723;
wire            n3724;
wire            n3725;
wire            n3726;
wire            n3728;
wire            n3729;
wire            n3730;
wire            n3731;
wire            n3732;
wire            n3733;
wire            n3734;
wire            n3735;
wire            n3736;
wire            n3737;
wire            n3738;
wire            n3739;
wire            n374;
wire            n3740;
wire            n3741;
wire            n3742;
wire            n3743;
wire            n3744;
wire            n3745;
wire            n3746;
wire            n3747;
wire            n3748;
wire            n3749;
wire            n3750;
wire            n3752;
wire            n3753;
wire            n3754;
wire            n3755;
wire            n3756;
wire            n3757;
wire            n3758;
wire            n3759;
wire            n376;
wire            n3760;
wire            n3761;
wire            n3762;
wire            n3763;
wire            n3764;
wire            n3765;
wire            n3766;
wire            n3767;
wire            n3768;
wire            n3769;
wire            n3770;
wire            n3771;
wire            n3772;
wire            n3773;
wire            n3774;
wire            n3776;
wire            n3777;
wire            n3778;
wire            n3779;
wire            n378;
wire            n3780;
wire            n3781;
wire            n3782;
wire            n3783;
wire            n3784;
wire            n3785;
wire            n3786;
wire            n3787;
wire            n3788;
wire            n3789;
wire            n3790;
wire            n3791;
wire            n3792;
wire            n3793;
wire            n3794;
wire            n3795;
wire            n3796;
wire            n3797;
wire            n3798;
wire            n38;
wire            n380;
wire            n3800;
wire            n3801;
wire            n3802;
wire            n3803;
wire            n3804;
wire            n3805;
wire            n3806;
wire            n3807;
wire            n3808;
wire            n3809;
wire            n3810;
wire            n3811;
wire            n3812;
wire            n3813;
wire            n3814;
wire            n3815;
wire            n3816;
wire            n3817;
wire            n3818;
wire            n3819;
wire            n382;
wire            n3820;
wire            n3821;
wire            n3822;
wire            n3824;
wire            n3825;
wire            n3826;
wire            n3827;
wire            n3828;
wire            n3829;
wire            n3830;
wire            n3831;
wire            n3832;
wire            n3833;
wire            n3834;
wire            n3835;
wire            n3836;
wire            n3837;
wire            n3838;
wire            n3839;
wire            n384;
wire            n3840;
wire            n3841;
wire            n3842;
wire            n3843;
wire            n3844;
wire            n3845;
wire            n3846;
wire            n3848;
wire            n3849;
wire            n3850;
wire            n3851;
wire            n3852;
wire            n3853;
wire            n3854;
wire            n3855;
wire            n3856;
wire            n3857;
wire            n3858;
wire            n3859;
wire            n386;
wire            n3860;
wire            n3861;
wire            n3862;
wire            n3863;
wire            n3864;
wire            n3865;
wire            n3866;
wire            n3867;
wire            n3868;
wire            n3869;
wire            n3870;
wire            n3872;
wire            n3873;
wire            n3874;
wire            n3875;
wire            n3876;
wire            n3877;
wire            n3878;
wire            n3879;
wire            n388;
wire            n3880;
wire            n3881;
wire            n3882;
wire            n3883;
wire            n3884;
wire            n3885;
wire            n3886;
wire            n3887;
wire            n3888;
wire            n3889;
wire            n3890;
wire            n3891;
wire            n3892;
wire            n3893;
wire            n3894;
wire            n3895;
wire            n3896;
wire            n3897;
wire            n3898;
wire            n3899;
wire            n39;
wire            n390;
wire            n3900;
wire            n3901;
wire            n3902;
wire            n3903;
wire            n3904;
wire      [4:0] n3905;
wire      [4:0] n3906;
wire            n3907;
wire            n3908;
wire            n3909;
wire      [2:0] n3910;
wire            n3911;
wire            n3912;
wire      [4:0] n3913;
wire            n3914;
wire      [4:0] n3915;
wire            n3916;
wire            n3917;
wire      [4:0] n3918;
wire            n3919;
wire            n392;
wire            n3920;
wire      [4:0] n3921;
wire            n3922;
wire            n3923;
wire      [4:0] n3924;
wire            n3925;
wire            n3926;
wire      [4:0] n3927;
wire            n3928;
wire            n3929;
wire      [4:0] n3930;
wire            n3931;
wire            n3932;
wire            n3933;
wire      [2:0] n3934;
wire            n3935;
wire      [7:0] n3937;
wire            n3938;
wire            n3939;
wire            n394;
wire            n3940;
wire            n3941;
wire            n3942;
wire            n3943;
wire            n3944;
wire            n3945;
wire            n3946;
wire            n3947;
wire            n3948;
wire            n3949;
wire            n3950;
wire            n3951;
wire            n3952;
wire            n3953;
wire            n3954;
wire            n3955;
wire            n3956;
wire            n3957;
wire            n3958;
wire            n3959;
wire            n396;
wire      [4:0] n3960;
wire            n3961;
wire            n3962;
wire            n3963;
wire            n3964;
wire            n3965;
wire            n3966;
wire            n3967;
wire            n3968;
wire            n3969;
wire            n3970;
wire            n3971;
wire            n3972;
wire            n3973;
wire            n3974;
wire            n3975;
wire            n3976;
wire            n3977;
wire            n3978;
wire            n3979;
wire            n398;
wire            n3980;
wire            n3981;
wire            n3982;
wire            n3983;
wire            n3984;
wire            n3985;
wire            n3986;
wire            n3987;
wire            n3989;
wire            n3990;
wire            n3991;
wire            n3992;
wire            n3993;
wire            n3994;
wire            n3995;
wire            n3996;
wire            n3997;
wire            n3998;
wire            n3999;
wire            n40;
wire            n400;
wire            n4000;
wire            n4001;
wire            n4002;
wire            n4003;
wire            n4004;
wire            n4005;
wire            n4006;
wire            n4007;
wire            n4008;
wire            n4009;
wire            n4010;
wire            n4011;
wire            n4012;
wire            n4013;
wire            n4014;
wire            n4015;
wire            n4016;
wire            n4017;
wire            n4018;
wire            n4019;
wire            n402;
wire            n4020;
wire            n4021;
wire            n4022;
wire            n4023;
wire            n4024;
wire            n4025;
wire            n4026;
wire            n4027;
wire            n4028;
wire            n4029;
wire            n4030;
wire            n4031;
wire            n4032;
wire            n4033;
wire            n4034;
wire            n4035;
wire            n4036;
wire            n4037;
wire            n4038;
wire            n4039;
wire            n404;
wire            n4040;
wire            n4041;
wire            n4042;
wire            n4043;
wire            n4044;
wire            n4045;
wire            n4046;
wire            n4047;
wire            n4048;
wire            n4049;
wire            n4050;
wire            n4051;
wire            n4052;
wire            n4053;
wire            n4054;
wire            n4055;
wire            n4056;
wire            n4057;
wire            n4058;
wire            n4059;
wire            n406;
wire            n4060;
wire            n4061;
wire            n4062;
wire            n4063;
wire            n4064;
wire            n4065;
wire            n4066;
wire            n4067;
wire            n4068;
wire            n4069;
wire            n4070;
wire            n4071;
wire            n4072;
wire            n4073;
wire            n4074;
wire            n4075;
wire            n4076;
wire            n4077;
wire            n4078;
wire            n4079;
wire            n408;
wire            n4080;
wire            n4081;
wire            n4082;
wire            n4083;
wire            n4084;
wire            n4085;
wire            n4086;
wire            n4087;
wire            n4088;
wire            n4089;
wire            n4090;
wire            n4091;
wire            n4092;
wire            n4093;
wire            n4094;
wire            n4095;
wire            n4096;
wire            n4097;
wire            n4098;
wire            n4099;
wire            n41;
wire            n410;
wire            n4100;
wire            n4101;
wire            n4102;
wire            n4103;
wire            n4104;
wire            n4105;
wire            n4106;
wire            n4107;
wire            n4108;
wire            n4109;
wire            n4110;
wire            n4111;
wire            n4112;
wire            n4113;
wire            n4114;
wire            n4115;
wire            n4116;
wire            n4117;
wire            n4118;
wire            n4119;
wire            n412;
wire            n4120;
wire            n4121;
wire            n4122;
wire            n4123;
wire            n4124;
wire            n4125;
wire            n4126;
wire            n4127;
wire            n4128;
wire            n4129;
wire            n4130;
wire            n4131;
wire            n4132;
wire            n4133;
wire            n4134;
wire            n4135;
wire            n4136;
wire            n4137;
wire            n4138;
wire            n4139;
wire            n414;
wire            n4140;
wire            n4141;
wire            n4142;
wire            n4143;
wire            n4144;
wire            n4145;
wire            n4146;
wire            n4147;
wire            n4148;
wire            n4149;
wire            n4150;
wire            n4151;
wire            n4152;
wire            n4153;
wire            n4154;
wire            n4155;
wire            n4156;
wire            n4157;
wire            n4158;
wire            n4159;
wire            n416;
wire            n4160;
wire            n4161;
wire            n4162;
wire            n4163;
wire            n4164;
wire            n4165;
wire            n4166;
wire            n4167;
wire            n4168;
wire            n4169;
wire            n4170;
wire            n4171;
wire            n4172;
wire            n4173;
wire            n4174;
wire            n4175;
wire            n4176;
wire            n4177;
wire            n4178;
wire            n4179;
wire            n418;
wire            n4180;
wire            n4181;
wire            n4182;
wire            n4183;
wire            n4184;
wire            n4185;
wire            n4186;
wire            n4187;
wire            n4188;
wire            n4189;
wire            n4190;
wire            n4191;
wire            n4192;
wire            n4193;
wire            n4194;
wire            n4195;
wire            n4196;
wire            n4197;
wire            n4198;
wire            n4199;
wire            n42;
wire            n420;
wire            n4200;
wire            n4201;
wire            n4202;
wire            n4203;
wire            n4204;
wire            n4205;
wire            n4206;
wire            n4207;
wire            n4208;
wire            n4209;
wire      [4:0] n4210;
wire            n4211;
wire            n4212;
wire      [2:0] n4213;
wire            n4214;
wire            n4215;
wire            n4216;
wire            n4217;
wire            n4218;
wire            n4219;
wire            n422;
wire            n4220;
wire            n4221;
wire            n4222;
wire            n4223;
wire            n4224;
wire            n4225;
wire            n4226;
wire            n4227;
wire            n4228;
wire            n4229;
wire            n4230;
wire            n4231;
wire            n4232;
wire            n4233;
wire            n4234;
wire            n4235;
wire            n4236;
wire            n4237;
wire            n4238;
wire            n4239;
wire            n424;
wire            n4240;
wire            n4241;
wire            n4242;
wire            n4243;
wire            n4244;
wire            n4245;
wire            n4246;
wire            n4247;
wire            n4248;
wire            n4249;
wire            n4250;
wire            n4251;
wire            n4252;
wire            n4253;
wire            n4254;
wire            n4255;
wire            n4256;
wire            n4257;
wire            n4258;
wire            n4259;
wire            n426;
wire            n4260;
wire            n4261;
wire            n4262;
wire            n4263;
wire            n4264;
wire            n4265;
wire            n4266;
wire            n4267;
wire            n4268;
wire            n4269;
wire            n4270;
wire            n4271;
wire            n4272;
wire            n4273;
wire            n4274;
wire            n4275;
wire            n4276;
wire            n4277;
wire            n4278;
wire            n4279;
wire            n428;
wire            n4280;
wire            n4281;
wire            n4282;
wire            n4283;
wire            n4284;
wire            n4285;
wire            n4286;
wire            n4287;
wire            n4288;
wire            n4289;
wire            n4290;
wire            n4291;
wire            n4292;
wire            n4293;
wire            n4294;
wire            n4295;
wire            n4296;
wire            n4297;
wire            n4298;
wire            n4299;
wire            n43;
wire            n430;
wire            n4300;
wire            n4301;
wire            n4302;
wire            n4303;
wire            n4304;
wire            n4305;
wire            n4306;
wire            n4307;
wire            n4308;
wire            n4309;
wire            n4310;
wire            n4311;
wire            n4312;
wire            n4313;
wire            n4314;
wire            n4315;
wire            n4316;
wire            n4317;
wire            n4318;
wire            n4319;
wire            n432;
wire            n4320;
wire            n4321;
wire            n4322;
wire            n4323;
wire            n4324;
wire            n4325;
wire            n4326;
wire            n4327;
wire            n4328;
wire            n4329;
wire            n4330;
wire            n4331;
wire            n4332;
wire            n4333;
wire            n4334;
wire            n4335;
wire            n4336;
wire            n4337;
wire            n4338;
wire            n4339;
wire            n434;
wire            n4340;
wire            n4341;
wire            n4342;
wire            n4343;
wire            n4344;
wire            n4345;
wire            n4346;
wire            n4347;
wire            n4348;
wire            n4349;
wire            n4350;
wire            n4351;
wire            n4352;
wire            n4353;
wire            n4354;
wire            n4355;
wire            n4356;
wire            n4357;
wire            n4358;
wire            n4359;
wire            n436;
wire            n4360;
wire            n4361;
wire            n4362;
wire            n4363;
wire            n4364;
wire            n4365;
wire            n4366;
wire            n4367;
wire            n4368;
wire            n4369;
wire            n4370;
wire            n4371;
wire            n4372;
wire            n4373;
wire            n4374;
wire            n4375;
wire            n4376;
wire            n4377;
wire            n4378;
wire            n4379;
wire            n438;
wire            n4380;
wire            n4381;
wire            n4382;
wire            n4383;
wire            n4384;
wire            n4385;
wire            n4386;
wire            n4387;
wire            n4388;
wire            n4389;
wire            n4390;
wire            n4391;
wire            n4392;
wire            n4393;
wire            n4394;
wire            n4395;
wire            n4396;
wire            n4397;
wire            n4398;
wire            n4399;
wire      [3:0] n44;
wire            n440;
wire            n4400;
wire            n4401;
wire            n4402;
wire            n4403;
wire            n4404;
wire            n4405;
wire            n4406;
wire            n4407;
wire            n4408;
wire            n4409;
wire            n4410;
wire            n4411;
wire            n4412;
wire            n4413;
wire            n4414;
wire            n4415;
wire            n4416;
wire            n4417;
wire            n4418;
wire            n4419;
wire            n442;
wire            n4420;
wire            n4421;
wire            n4422;
wire            n4423;
wire            n4424;
wire            n4425;
wire            n4426;
wire            n4427;
wire            n4428;
wire            n4429;
wire            n4430;
wire            n4431;
wire            n4432;
wire            n4433;
wire            n4434;
wire            n4435;
wire            n4436;
wire            n4437;
wire            n4438;
wire            n4439;
wire            n444;
wire            n4440;
wire            n4441;
wire            n4442;
wire            n4443;
wire            n4444;
wire            n4445;
wire            n4446;
wire            n4447;
wire            n4448;
wire            n4449;
wire            n4450;
wire            n4451;
wire            n4452;
wire      [4:0] n4453;
wire      [4:0] n4454;
wire            n4455;
wire            n4456;
wire            n4457;
wire      [2:0] n4458;
wire            n4459;
wire            n446;
wire            n4460;
wire            n4461;
wire      [2:0] n4462;
wire            n4463;
wire            n4464;
wire            n4465;
wire            n4466;
wire            n4467;
wire            n4468;
wire            n4469;
wire            n4470;
wire            n4471;
wire            n4472;
wire            n4473;
wire            n4474;
wire            n4475;
wire            n4476;
wire            n4477;
wire            n4478;
wire            n4479;
wire            n448;
wire            n4480;
wire            n4481;
wire            n4482;
wire            n4483;
wire            n4484;
wire            n4485;
wire      [4:0] n4486;
wire            n4487;
wire            n4488;
wire            n4489;
wire            n4490;
wire            n4491;
wire            n4492;
wire            n4493;
wire            n4494;
wire            n4495;
wire            n4496;
wire            n4497;
wire            n4498;
wire            n4499;
wire      [4:0] n45;
wire            n450;
wire            n4500;
wire            n4501;
wire            n4502;
wire            n4503;
wire            n4504;
wire            n4505;
wire            n4506;
wire            n4507;
wire            n4508;
wire            n4509;
wire            n4510;
wire            n4511;
wire            n4512;
wire            n4513;
wire            n4514;
wire            n4515;
wire            n4516;
wire            n4517;
wire            n4518;
wire            n4519;
wire            n452;
wire            n4520;
wire            n4521;
wire            n4522;
wire            n4523;
wire            n4524;
wire            n4525;
wire            n4526;
wire            n4527;
wire            n4528;
wire            n4529;
wire            n4530;
wire            n4531;
wire            n4532;
wire            n4533;
wire            n4534;
wire            n4535;
wire            n4536;
wire            n4537;
wire            n4538;
wire            n4539;
wire            n454;
wire            n4540;
wire            n4541;
wire            n4542;
wire            n4543;
wire            n4544;
wire            n4545;
wire            n4546;
wire            n4547;
wire            n4548;
wire            n4549;
wire            n4550;
wire            n4551;
wire            n4552;
wire            n4553;
wire            n4554;
wire            n4555;
wire            n4556;
wire            n4557;
wire            n4558;
wire            n4559;
wire            n456;
wire            n4560;
wire            n4561;
wire            n4562;
wire            n4563;
wire            n4564;
wire            n4565;
wire            n4566;
wire            n4567;
wire            n4568;
wire            n4569;
wire            n4570;
wire            n4571;
wire            n4572;
wire            n4573;
wire            n4574;
wire            n4575;
wire            n4576;
wire            n4577;
wire            n4578;
wire            n4579;
wire            n458;
wire            n4580;
wire            n4581;
wire            n4582;
wire            n4583;
wire            n4584;
wire            n4585;
wire            n4586;
wire            n4587;
wire            n4588;
wire            n4589;
wire            n4590;
wire            n4591;
wire            n4592;
wire            n4593;
wire            n4594;
wire            n4595;
wire            n4596;
wire            n4597;
wire            n4598;
wire            n4599;
wire            n460;
wire            n4600;
wire            n4601;
wire            n4602;
wire            n4603;
wire            n4604;
wire            n4605;
wire            n4606;
wire            n4607;
wire            n4608;
wire            n4609;
wire            n4610;
wire            n4611;
wire            n4612;
wire            n4613;
wire            n4614;
wire            n4615;
wire            n4616;
wire            n4617;
wire            n4618;
wire            n4619;
wire            n462;
wire            n4620;
wire            n4621;
wire            n4622;
wire            n4623;
wire            n4624;
wire            n4625;
wire            n4626;
wire            n4627;
wire            n4628;
wire            n4629;
wire            n4630;
wire            n4631;
wire            n4632;
wire            n4633;
wire            n4634;
wire            n4635;
wire            n4636;
wire            n4637;
wire            n4638;
wire            n4639;
wire            n464;
wire            n4640;
wire            n4641;
wire            n4642;
wire            n4643;
wire            n4644;
wire            n4645;
wire            n4646;
wire            n4647;
wire            n4648;
wire            n4649;
wire            n4650;
wire            n4651;
wire            n4652;
wire            n4653;
wire            n4654;
wire            n4655;
wire            n4656;
wire            n4657;
wire            n4658;
wire            n4659;
wire            n466;
wire            n4660;
wire            n4661;
wire            n4662;
wire            n4663;
wire            n4664;
wire            n4665;
wire            n4666;
wire            n4667;
wire            n4668;
wire            n4669;
wire            n4670;
wire            n4671;
wire            n4672;
wire            n4673;
wire            n4674;
wire            n4675;
wire            n4676;
wire            n4677;
wire            n4678;
wire            n4679;
wire            n468;
wire            n4680;
wire            n4681;
wire            n4682;
wire            n4683;
wire            n4684;
wire            n4685;
wire            n4686;
wire            n4687;
wire            n4688;
wire            n4689;
wire            n4690;
wire            n4691;
wire            n4692;
wire            n4693;
wire            n4694;
wire            n4695;
wire            n4696;
wire            n4697;
wire            n4698;
wire            n4699;
wire      [7:0] n47;
wire            n470;
wire            n4700;
wire            n4701;
wire            n4702;
wire            n4703;
wire            n4704;
wire            n4705;
wire            n4706;
wire            n4707;
wire            n4708;
wire            n4709;
wire            n4710;
wire            n4711;
wire            n4712;
wire            n4713;
wire            n4714;
wire            n4715;
wire            n4716;
wire            n4717;
wire            n4718;
wire            n4719;
wire            n472;
wire            n4720;
wire            n4721;
wire            n4722;
wire            n4723;
wire            n4724;
wire            n4725;
wire            n4726;
wire            n4727;
wire            n4728;
wire            n4729;
wire            n4730;
wire            n4731;
wire            n4732;
wire            n4733;
wire            n4734;
wire            n4735;
wire            n4736;
wire            n4737;
wire            n4738;
wire            n4739;
wire            n474;
wire            n4740;
wire            n4741;
wire            n4742;
wire            n4743;
wire            n4744;
wire            n4745;
wire            n4746;
wire            n4747;
wire            n4748;
wire            n4749;
wire            n4750;
wire            n4751;
wire            n4752;
wire            n4753;
wire            n4754;
wire            n4755;
wire            n4756;
wire            n4757;
wire      [7:0] n4758;
wire            n4759;
wire            n476;
wire            n4760;
wire      [7:0] n4761;
wire            n4762;
wire      [7:0] n4763;
wire            n4764;
wire      [7:0] n4765;
wire      [7:0] n4766;
wire      [7:0] n4767;
wire      [7:0] n4768;
wire      [7:0] n4769;
wire      [7:0] n4770;
wire            n4772;
wire            n4773;
wire            n4774;
wire            n4775;
wire      [7:0] n4776;
wire            n4777;
wire            n4778;
wire      [7:0] n4779;
wire            n478;
wire      [7:0] n4780;
wire      [7:0] n4781;
wire      [7:0] n4782;
wire            n4783;
wire            n4784;
wire      [7:0] n4785;
wire      [7:0] n4786;
wire      [7:0] n4787;
wire            n4788;
wire            n4789;
wire            n4790;
wire            n4791;
wire            n4792;
wire            n4793;
wire            n4794;
wire            n4795;
wire            n4796;
wire            n4797;
wire            n4798;
wire            n4799;
wire      [3:0] n48;
wire            n480;
wire            n4800;
wire            n4801;
wire            n4802;
wire            n4803;
wire            n4804;
wire      [7:0] n4805;
wire            n4806;
wire            n4807;
wire      [7:0] n4808;
wire      [7:0] n4809;
wire      [7:0] n4810;
wire            n4811;
wire            n4812;
wire            n4813;
wire            n4814;
wire            n4815;
wire      [7:0] n4816;
wire            n4817;
wire            n4818;
wire      [7:0] n4819;
wire            n482;
wire            n4820;
wire      [7:0] n4821;
wire            n4822;
wire      [7:0] n4823;
wire      [7:0] n4824;
wire      [7:0] n4825;
wire      [7:0] n4826;
wire      [7:0] n4827;
wire      [7:0] n4828;
wire     [15:0] n4829;
wire     [15:0] n4831;
wire      [7:0] n4832;
wire     [15:0] n4833;
wire     [15:0] n4834;
wire      [7:0] n4835;
wire      [7:0] n4836;
wire            n4837;
wire            n4838;
wire      [7:0] n4839;
wire            n484;
wire      [7:0] n4840;
wire      [7:0] n4841;
wire            n4842;
wire            n4843;
wire      [7:0] n4844;
wire      [7:0] n4845;
wire      [7:0] n4846;
wire            n4847;
wire            n4848;
wire            n4849;
wire            n4850;
wire            n4851;
wire            n4852;
wire            n4853;
wire      [7:0] n4854;
wire            n4855;
wire            n4856;
wire      [7:0] n4857;
wire            n4858;
wire      [7:0] n4859;
wire            n486;
wire            n4860;
wire      [7:0] n4861;
wire      [7:0] n4862;
wire      [7:0] n4863;
wire      [7:0] n4864;
wire      [7:0] n4865;
wire      [7:0] n4866;
wire      [7:0] n4867;
wire            n4868;
wire            n4869;
wire      [7:0] n4870;
wire      [7:0] n4871;
wire      [7:0] n4872;
wire            n4873;
wire            n4874;
wire            n4875;
wire            n4876;
wire            n4877;
wire            n4878;
wire            n4879;
wire            n488;
wire            n4880;
wire            n4881;
wire            n4882;
wire            n4883;
wire            n4884;
wire            n4885;
wire            n4886;
wire            n4887;
wire            n4888;
wire            n4889;
wire            n4890;
wire            n4891;
wire            n4892;
wire            n4893;
wire      [7:0] n4894;
wire            n4895;
wire            n4896;
wire      [7:0] n4897;
wire            n4898;
wire      [7:0] n4899;
wire      [7:0] n49;
wire            n490;
wire            n4900;
wire      [7:0] n4901;
wire      [7:0] n4902;
wire      [7:0] n4903;
wire      [7:0] n4904;
wire      [7:0] n4905;
wire      [7:0] n4906;
wire      [3:0] n4907;
wire            n4908;
wire            n4909;
wire      [3:0] n4910;
wire      [4:0] n4911;
wire      [4:0] n4913;
wire      [3:0] n4914;
wire      [4:0] n4915;
wire      [4:0] n4916;
wire            n4917;
wire            n4918;
wire            n4919;
wire            n492;
wire      [3:0] n4920;
wire            n4921;
wire            n4922;
wire      [3:0] n4923;
wire      [4:0] n4924;
wire      [4:0] n4925;
wire            n4926;
wire      [4:0] n4927;
wire      [4:0] n4928;
wire      [3:0] n4929;
wire      [4:0] n4930;
wire            n4931;
wire      [4:0] n4932;
wire      [4:0] n4933;
wire      [4:0] n4934;
wire      [3:0] n4935;
wire      [3:0] n4936;
wire      [7:0] n4937;
wire            n4938;
wire            n4939;
wire            n494;
wire      [7:0] n4940;
wire      [7:0] n4941;
wire      [7:0] n4942;
wire            n4943;
wire      [7:0] n4945;
wire            n4946;
wire      [7:0] n4948;
wire            n4949;
wire            n4950;
wire      [7:0] n4951;
wire      [7:0] n4952;
wire      [7:0] n4953;
wire            n4954;
wire      [7:0] n4956;
wire            n4957;
wire      [7:0] n4959;
wire            n496;
wire            n4960;
wire            n4961;
wire      [7:0] n4962;
wire      [7:0] n4963;
wire      [7:0] n4964;
wire            n4965;
wire            n4966;
wire            n4967;
wire            n4968;
wire            n4969;
wire            n4970;
wire            n4971;
wire      [7:0] n4972;
wire            n4973;
wire            n4974;
wire      [7:0] n4975;
wire            n4976;
wire      [7:0] n4977;
wire            n4978;
wire      [7:0] n4979;
wire            n498;
wire      [7:0] n4980;
wire      [7:0] n4981;
wire      [7:0] n4982;
wire      [7:0] n4983;
wire      [7:0] n4984;
wire            n4985;
wire      [1:0] n4986;
wire            n4987;
wire            n4988;
wire            n4989;
wire            n4990;
wire      [7:0] n4991;
wire            n4992;
wire            n4993;
wire      [7:0] n4994;
wire      [7:0] n4995;
wire      [7:0] n4996;
wire            n4997;
wire      [1:0] n4998;
wire      [1:0] n4999;
wire            n5;
wire      [7:0] n50;
wire            n500;
wire      [2:0] n5000;
wire      [3:0] n5001;
wire      [2:0] n5002;
wire      [3:0] n5003;
wire      [3:0] n5004;
wire      [3:0] n5005;
wire      [4:0] n5006;
wire      [3:0] n5007;
wire      [4:0] n5008;
wire      [4:0] n5009;
wire            n5010;
wire            n5011;
wire            n5012;
wire            n5013;
wire            n5014;
wire            n5015;
wire            n5016;
wire            n5017;
wire            n5018;
wire            n5019;
wire            n502;
wire            n5020;
wire      [4:0] n5021;
wire      [4:0] n5022;
wire            n5023;
wire            n5024;
wire      [3:0] n5025;
wire      [3:0] n5026;
wire            n5027;
wire            n5028;
wire      [1:0] n5029;
wire      [1:0] n5030;
wire            n5031;
wire      [2:0] n5032;
wire      [3:0] n5033;
wire      [3:0] n5034;
wire      [7:0] n5035;
wire            n5036;
wire            n5037;
wire      [7:0] n5038;
wire      [7:0] n5039;
wire            n504;
wire      [7:0] n5040;
wire            n5041;
wire            n5042;
wire            n5043;
wire            n5044;
wire            n5045;
wire            n5046;
wire            n5047;
wire      [7:0] n5048;
wire            n5049;
wire            n5050;
wire      [7:0] n5051;
wire            n5052;
wire      [7:0] n5053;
wire            n5054;
wire      [7:0] n5055;
wire      [7:0] n5056;
wire      [7:0] n5057;
wire      [7:0] n5058;
wire      [7:0] n5059;
wire            n506;
wire      [7:0] n5060;
wire            n5061;
wire            n5062;
wire            n5063;
wire            n5064;
wire      [7:0] n5065;
wire            n5066;
wire            n5067;
wire      [7:0] n5068;
wire      [7:0] n5069;
wire      [7:0] n5070;
wire      [7:0] n5071;
wire            n5072;
wire            n5073;
wire      [7:0] n5074;
wire      [7:0] n5075;
wire      [7:0] n5076;
wire            n5077;
wire            n5078;
wire            n5079;
wire            n508;
wire            n5080;
wire            n5081;
wire            n5082;
wire            n5083;
wire      [7:0] n5084;
wire            n5085;
wire            n5086;
wire      [7:0] n5087;
wire            n5088;
wire      [7:0] n5089;
wire            n5090;
wire      [7:0] n5091;
wire      [7:0] n5092;
wire      [7:0] n5093;
wire      [7:0] n5094;
wire      [7:0] n5095;
wire      [7:0] n5096;
wire      [6:0] n5097;
wire            n5098;
wire      [7:0] n5099;
wire      [7:0] n51;
wire            n510;
wire            n5100;
wire            n5101;
wire      [7:0] n5102;
wire      [7:0] n5103;
wire      [7:0] n5104;
wire            n5105;
wire            n5106;
wire            n5107;
wire            n5108;
wire            n5109;
wire            n5110;
wire      [7:0] n5111;
wire            n5112;
wire            n5113;
wire      [7:0] n5114;
wire            n5115;
wire      [7:0] n5116;
wire            n5117;
wire      [7:0] n5118;
wire      [7:0] n5119;
wire            n512;
wire      [7:0] n5120;
wire      [7:0] n5121;
wire      [7:0] n5122;
wire      [7:0] n5123;
wire      [3:0] n5124;
wire      [3:0] n5125;
wire      [7:0] n5126;
wire            n5127;
wire      [6:0] n5128;
wire            n5129;
wire            n5130;
wire            n5131;
wire            n5132;
wire            n5133;
wire            n5134;
wire            n5135;
wire            n5136;
wire            n5137;
wire            n5138;
wire            n5139;
wire            n514;
wire      [7:0] n5140;
wire            n5141;
wire            n5142;
wire      [7:0] n5143;
wire      [7:0] n5144;
wire      [7:0] n5145;
wire            n5146;
wire            n5147;
wire            n5148;
wire            n5149;
wire            n5150;
wire            n5151;
wire            n5152;
wire      [7:0] n5153;
wire            n5154;
wire            n5155;
wire      [7:0] n5156;
wire            n5157;
wire      [7:0] n5158;
wire            n5159;
wire            n516;
wire      [7:0] n5160;
wire      [7:0] n5161;
wire      [7:0] n5162;
wire      [7:0] n5163;
wire      [7:0] n5164;
wire      [7:0] n5165;
wire            n5166;
wire      [6:0] n5167;
wire      [7:0] n5168;
wire            n5169;
wire            n5170;
wire      [7:0] n5171;
wire      [7:0] n5172;
wire      [7:0] n5173;
wire            n5174;
wire            n5175;
wire            n5176;
wire            n5177;
wire            n5178;
wire            n5179;
wire            n518;
wire            n5180;
wire            n5181;
wire            n5182;
wire            n5183;
wire            n5184;
wire            n5185;
wire            n5186;
wire            n5187;
wire            n5188;
wire            n5189;
wire            n5190;
wire            n5191;
wire      [7:0] n5192;
wire            n5193;
wire            n5194;
wire      [7:0] n5195;
wire            n5196;
wire      [7:0] n5197;
wire            n5198;
wire      [7:0] n5199;
wire            n52;
wire            n520;
wire      [7:0] n5200;
wire      [7:0] n5201;
wire      [7:0] n5202;
wire      [7:0] n5203;
wire      [7:0] n5204;
wire      [6:0] n5205;
wire      [7:0] n5206;
wire            n5207;
wire            n5208;
wire      [7:0] n5209;
wire      [7:0] n5210;
wire      [7:0] n5211;
wire            n5212;
wire            n5213;
wire            n5214;
wire            n5215;
wire            n5216;
wire            n5217;
wire            n5218;
wire            n5219;
wire            n522;
wire            n5220;
wire            n5221;
wire            n5222;
wire            n5223;
wire            n5224;
wire            n5225;
wire            n5226;
wire            n5227;
wire            n5228;
wire            n5229;
wire      [7:0] n5230;
wire            n5231;
wire            n5232;
wire      [7:0] n5233;
wire            n5234;
wire      [7:0] n5235;
wire            n5236;
wire      [7:0] n5237;
wire      [7:0] n5238;
wire      [7:0] n5239;
wire            n524;
wire      [7:0] n5240;
wire      [7:0] n5241;
wire      [7:0] n5242;
wire            n5243;
wire            n5244;
wire            n5245;
wire            n5246;
wire      [7:0] n5247;
wire            n5248;
wire            n5249;
wire      [7:0] n5250;
wire      [7:0] n5251;
wire      [7:0] n5252;
wire      [3:0] n5253;
wire      [3:0] n5254;
wire      [7:0] n5255;
wire      [7:0] n5256;
wire            n5257;
wire            n5258;
wire      [3:0] n5259;
wire            n526;
wire      [3:0] n5260;
wire      [7:0] n5261;
wire      [7:0] n5262;
wire            n5263;
wire            n5264;
wire      [7:0] n5265;
wire      [7:0] n5266;
wire      [7:0] n5267;
wire            n5268;
wire            n5269;
wire            n5270;
wire            n5271;
wire            n5272;
wire            n5273;
wire            n5274;
wire      [7:0] n5275;
wire            n5276;
wire            n5277;
wire      [7:0] n5278;
wire            n5279;
wire            n528;
wire      [7:0] n5280;
wire            n5281;
wire      [7:0] n5282;
wire      [7:0] n5283;
wire      [7:0] n5284;
wire      [7:0] n5285;
wire      [7:0] n5286;
wire      [7:0] n5287;
wire            n5288;
wire            n5289;
wire            n5290;
wire            n5291;
wire      [7:0] n5292;
wire            n5293;
wire            n5294;
wire      [7:0] n5295;
wire      [7:0] n5296;
wire      [7:0] n5297;
wire      [7:0] n5298;
wire            n5299;
wire            n530;
wire            n5300;
wire      [7:0] n5301;
wire      [7:0] n5302;
wire      [7:0] n5303;
wire            n5304;
wire            n5305;
wire      [7:0] n5306;
wire      [7:0] n5307;
wire            n5308;
wire            n5309;
wire            n5310;
wire            n5311;
wire            n5312;
wire      [7:0] n5313;
wire            n5314;
wire            n5315;
wire      [7:0] n5316;
wire            n5317;
wire      [7:0] n5318;
wire            n5319;
wire            n532;
wire      [7:0] n5320;
wire      [7:0] n5321;
wire      [7:0] n5322;
wire      [7:0] n5323;
wire      [7:0] n5324;
wire      [7:0] n5325;
wire            n5326;
wire      [1:0] n5327;
wire            n5328;
wire            n5329;
wire            n5330;
wire            n5331;
wire      [7:0] n5332;
wire            n5333;
wire            n5334;
wire      [7:0] n5335;
wire      [7:0] n5336;
wire      [7:0] n5337;
wire            n5338;
wire      [1:0] n5339;
wire            n534;
wire      [1:0] n5340;
wire      [2:0] n5341;
wire      [3:0] n5342;
wire      [2:0] n5343;
wire      [3:0] n5344;
wire      [3:0] n5345;
wire      [3:0] n5346;
wire      [4:0] n5347;
wire      [3:0] n5348;
wire      [4:0] n5349;
wire      [4:0] n5350;
wire            n5351;
wire            n5352;
wire            n5353;
wire            n5354;
wire            n5355;
wire            n5356;
wire            n5357;
wire            n5358;
wire            n5359;
wire            n536;
wire            n5360;
wire            n5361;
wire      [4:0] n5362;
wire      [4:0] n5363;
wire            n5364;
wire      [3:0] n5365;
wire      [3:0] n5366;
wire            n5367;
wire      [1:0] n5368;
wire      [1:0] n5369;
wire            n5370;
wire      [7:0] n5371;
wire      [7:0] n5372;
wire            n5373;
wire            n5374;
wire      [2:0] n5375;
wire      [3:0] n5376;
wire      [3:0] n5377;
wire      [7:0] n5378;
wire            n5379;
wire            n538;
wire            n5380;
wire      [7:0] n5381;
wire      [7:0] n5382;
wire      [7:0] n5383;
wire            n5384;
wire            n5385;
wire      [7:0] n5386;
wire            n5387;
wire            n5388;
wire      [7:0] n5389;
wire            n5390;
wire            n5391;
wire      [7:0] n5392;
wire            n5393;
wire            n5394;
wire      [7:0] n5395;
wire            n5396;
wire            n5397;
wire      [7:0] n5398;
wire            n5399;
wire            n54;
wire            n540;
wire            n5400;
wire      [7:0] n5401;
wire            n5402;
wire            n5403;
wire      [7:0] n5404;
wire            n5405;
wire            n5406;
wire      [7:0] n5407;
wire            n5408;
wire            n5409;
wire      [7:0] n5410;
wire            n5411;
wire            n5412;
wire      [7:0] n5413;
wire            n5414;
wire            n5415;
wire      [7:0] n5416;
wire            n5417;
wire            n5418;
wire      [7:0] n5419;
wire            n542;
wire            n5420;
wire            n5421;
wire      [7:0] n5422;
wire            n5423;
wire            n5424;
wire      [7:0] n5425;
wire            n5426;
wire            n5427;
wire      [7:0] n5428;
wire            n5429;
wire            n5430;
wire            n5431;
wire      [7:0] n5432;
wire            n5433;
wire      [7:0] n5434;
wire      [7:0] n5435;
wire      [7:0] n5436;
wire      [7:0] n5437;
wire            n5438;
wire            n5439;
wire            n544;
wire            n5440;
wire      [7:0] n5441;
wire            n5442;
wire      [7:0] n5443;
wire      [7:0] n5444;
wire      [7:0] n5445;
wire      [7:0] n5446;
wire            n5447;
wire            n5448;
wire      [7:0] n5449;
wire            n5450;
wire      [7:0] n5451;
wire            n5452;
wire      [7:0] n5453;
wire      [7:0] n5454;
wire      [7:0] n5455;
wire      [7:0] n5456;
wire            n5457;
wire            n5458;
wire            n5459;
wire            n546;
wire      [7:0] n5460;
wire            n5461;
wire      [7:0] n5462;
wire      [7:0] n5463;
wire      [7:0] n5464;
wire      [7:0] n5465;
wire            n5466;
wire            n5467;
wire            n5468;
wire            n5469;
wire            n5470;
wire            n5471;
wire            n5472;
wire      [7:0] n5473;
wire            n5474;
wire            n5475;
wire      [7:0] n5476;
wire            n5477;
wire      [7:0] n5478;
wire            n5479;
wire            n548;
wire      [7:0] n5480;
wire      [7:0] n5481;
wire      [7:0] n5482;
wire      [7:0] n5483;
wire      [7:0] n5484;
wire      [7:0] n5485;
wire            n5486;
wire      [7:0] n5487;
wire            n5488;
wire      [7:0] n5489;
wire      [7:0] n5490;
wire      [7:0] n5491;
wire      [7:0] n5492;
wire            n5493;
wire            n5494;
wire            n5495;
wire            n5496;
wire            n5497;
wire            n5498;
wire            n5499;
wire            n55;
wire            n550;
wire      [7:0] n5500;
wire            n5501;
wire            n5502;
wire      [7:0] n5503;
wire            n5504;
wire      [7:0] n5505;
wire            n5506;
wire      [7:0] n5507;
wire      [7:0] n5508;
wire      [7:0] n5509;
wire      [7:0] n5510;
wire      [7:0] n5511;
wire      [7:0] n5512;
wire            n5513;
wire      [7:0] n5514;
wire            n5515;
wire      [7:0] n5516;
wire      [7:0] n5517;
wire      [7:0] n5518;
wire      [7:0] n5519;
wire            n552;
wire            n5520;
wire            n5521;
wire            n5522;
wire      [7:0] n5523;
wire            n5524;
wire      [7:0] n5525;
wire      [7:0] n5526;
wire      [7:0] n5527;
wire      [7:0] n5528;
wire            n5529;
wire            n5530;
wire            n5531;
wire      [7:0] n5532;
wire            n5533;
wire      [7:0] n5534;
wire      [7:0] n5535;
wire      [7:0] n5536;
wire      [7:0] n5537;
wire            n5538;
wire            n5539;
wire            n554;
wire            n5540;
wire      [7:0] n5541;
wire            n5542;
wire      [7:0] n5543;
wire      [7:0] n5544;
wire      [7:0] n5545;
wire      [7:0] n5546;
wire            n5547;
wire            n5548;
wire            n5549;
wire      [7:0] n5550;
wire            n5551;
wire      [7:0] n5552;
wire      [7:0] n5553;
wire      [7:0] n5554;
wire      [7:0] n5555;
wire            n5556;
wire            n5557;
wire            n5558;
wire      [7:0] n5559;
wire            n556;
wire            n5560;
wire      [7:0] n5561;
wire      [7:0] n5562;
wire      [7:0] n5563;
wire      [7:0] n5564;
wire            n5565;
wire            n5566;
wire            n5567;
wire      [7:0] n5568;
wire            n5569;
wire      [7:0] n5570;
wire      [7:0] n5571;
wire      [7:0] n5572;
wire      [7:0] n5573;
wire            n5574;
wire            n5575;
wire            n5576;
wire      [7:0] n5577;
wire            n5578;
wire      [7:0] n5579;
wire            n558;
wire      [7:0] n5580;
wire      [7:0] n5581;
wire      [7:0] n5582;
wire            n5583;
wire            n5584;
wire            n5585;
wire      [7:0] n5586;
wire            n5587;
wire      [7:0] n5588;
wire      [7:0] n5589;
wire      [7:0] n5590;
wire      [7:0] n5591;
wire            n5592;
wire            n5593;
wire            n5594;
wire      [7:0] n5595;
wire      [7:0] n5596;
wire            n5597;
wire            n5598;
wire            n5599;
wire      [2:0] n56;
wire            n560;
wire      [7:0] n5600;
wire      [7:0] n5601;
wire            n5602;
wire            n5603;
wire            n5604;
wire      [7:0] n5605;
wire      [7:0] n5606;
wire            n5607;
wire            n5608;
wire            n5609;
wire      [7:0] n5610;
wire      [7:0] n5611;
wire            n5612;
wire            n5613;
wire            n5614;
wire      [7:0] n5615;
wire      [7:0] n5616;
wire            n5617;
wire            n5618;
wire            n5619;
wire            n562;
wire      [7:0] n5620;
wire      [7:0] n5621;
wire            n5622;
wire            n5623;
wire            n5624;
wire      [7:0] n5625;
wire      [7:0] n5626;
wire            n5627;
wire            n5628;
wire            n5629;
wire      [7:0] n5630;
wire      [7:0] n5631;
wire            n5632;
wire            n5633;
wire            n5634;
wire      [7:0] n5635;
wire      [7:0] n5636;
wire            n5637;
wire            n5638;
wire            n5639;
wire            n564;
wire      [7:0] n5640;
wire      [7:0] n5641;
wire            n5642;
wire            n5643;
wire            n5644;
wire      [7:0] n5645;
wire      [7:0] n5646;
wire            n5647;
wire            n5648;
wire            n5649;
wire      [7:0] n5650;
wire      [7:0] n5651;
wire            n5652;
wire            n5653;
wire            n5654;
wire      [7:0] n5655;
wire      [7:0] n5656;
wire            n5657;
wire            n5658;
wire            n5659;
wire            n566;
wire      [7:0] n5660;
wire      [7:0] n5661;
wire            n5662;
wire            n5663;
wire            n5664;
wire      [7:0] n5665;
wire      [7:0] n5666;
wire            n5667;
wire            n5668;
wire            n5669;
wire      [7:0] n5670;
wire      [7:0] n5671;
wire            n5672;
wire            n5673;
wire            n5674;
wire      [7:0] n5675;
wire      [7:0] n5676;
wire            n5677;
wire            n5678;
wire            n5679;
wire            n568;
wire      [7:0] n5680;
wire      [7:0] n5681;
wire            n5682;
wire            n5683;
wire            n5684;
wire      [7:0] n5685;
wire      [7:0] n5686;
wire            n5687;
wire            n5688;
wire            n5689;
wire      [7:0] n5690;
wire      [7:0] n5691;
wire            n5692;
wire            n5693;
wire            n5694;
wire      [7:0] n5695;
wire      [7:0] n5696;
wire            n5697;
wire            n5698;
wire            n5699;
wire      [2:0] n57;
wire            n570;
wire      [7:0] n5700;
wire      [7:0] n5701;
wire            n5702;
wire            n5703;
wire            n5704;
wire      [7:0] n5705;
wire      [7:0] n5706;
wire            n5707;
wire            n5708;
wire            n5709;
wire      [7:0] n5710;
wire      [7:0] n5711;
wire            n5712;
wire            n5713;
wire            n5714;
wire      [7:0] n5715;
wire      [7:0] n5716;
wire            n5717;
wire            n5718;
wire            n5719;
wire            n572;
wire      [7:0] n5720;
wire      [7:0] n5721;
wire            n5722;
wire            n5723;
wire            n5724;
wire      [7:0] n5725;
wire      [7:0] n5726;
wire            n5727;
wire            n5728;
wire            n5729;
wire      [7:0] n5730;
wire      [7:0] n5731;
wire            n5732;
wire            n5733;
wire            n5734;
wire      [7:0] n5735;
wire      [7:0] n5736;
wire            n5737;
wire            n5738;
wire            n5739;
wire            n574;
wire      [7:0] n5740;
wire      [7:0] n5741;
wire            n5742;
wire            n5743;
wire      [7:0] n5744;
wire            n5745;
wire            n5746;
wire      [7:0] n5747;
wire            n5748;
wire            n5749;
wire      [7:0] n5750;
wire            n5751;
wire            n5752;
wire      [7:0] n5753;
wire            n5754;
wire            n5755;
wire      [7:0] n5756;
wire            n5757;
wire            n5758;
wire      [7:0] n5759;
wire            n576;
wire            n5760;
wire            n5761;
wire      [7:0] n5762;
wire            n5763;
wire            n5764;
wire      [7:0] n5765;
wire            n5766;
wire            n5767;
wire      [7:0] n5768;
wire            n5769;
wire            n5770;
wire      [7:0] n5771;
wire            n5772;
wire            n5773;
wire      [7:0] n5774;
wire            n5775;
wire            n5776;
wire      [7:0] n5777;
wire            n5778;
wire            n5779;
wire            n578;
wire      [7:0] n5780;
wire            n5781;
wire            n5782;
wire      [7:0] n5783;
wire            n5784;
wire            n5785;
wire      [7:0] n5786;
wire            n5787;
wire            n5788;
wire      [7:0] n5789;
wire      [7:0] n579;
wire            n5790;
wire            n5791;
wire      [7:0] n5792;
wire            n5793;
wire            n5794;
wire      [7:0] n5795;
wire            n5796;
wire            n5797;
wire      [7:0] n5798;
wire            n5799;
wire      [2:0] n58;
wire      [7:0] n580;
wire            n5800;
wire      [7:0] n5801;
wire            n5802;
wire            n5803;
wire      [7:0] n5804;
wire            n5805;
wire            n5806;
wire      [7:0] n5807;
wire            n5808;
wire            n5809;
wire      [7:0] n581;
wire      [7:0] n5810;
wire            n5811;
wire            n5812;
wire      [7:0] n5813;
wire            n5814;
wire            n5815;
wire      [7:0] n5816;
wire            n5817;
wire            n5818;
wire      [7:0] n5819;
wire      [7:0] n582;
wire            n5820;
wire            n5821;
wire      [7:0] n5822;
wire            n5823;
wire            n5824;
wire      [7:0] n5825;
wire            n5826;
wire            n5827;
wire      [7:0] n5828;
wire            n5829;
wire      [7:0] n583;
wire            n5830;
wire      [7:0] n5831;
wire            n5832;
wire            n5833;
wire      [7:0] n5834;
wire            n5835;
wire            n5836;
wire      [7:0] n5837;
wire            n5838;
wire            n5839;
wire      [7:0] n584;
wire      [7:0] n5840;
wire            n5841;
wire            n5842;
wire      [7:0] n5843;
wire            n5844;
wire            n5845;
wire      [7:0] n5846;
wire            n5847;
wire            n5848;
wire      [7:0] n5849;
wire      [7:0] n585;
wire            n5850;
wire            n5851;
wire      [7:0] n5852;
wire            n5853;
wire            n5854;
wire      [7:0] n5855;
wire            n5856;
wire            n5857;
wire      [7:0] n5858;
wire            n5859;
wire      [7:0] n586;
wire            n5860;
wire      [7:0] n5861;
wire            n5862;
wire            n5863;
wire      [7:0] n5864;
wire            n5865;
wire            n5866;
wire      [7:0] n5867;
wire            n5868;
wire            n5869;
wire      [7:0] n587;
wire      [7:0] n5870;
wire            n5871;
wire            n5872;
wire      [7:0] n5873;
wire            n5874;
wire            n5875;
wire      [7:0] n5876;
wire            n5877;
wire            n5878;
wire      [7:0] n5879;
wire      [7:0] n588;
wire            n5880;
wire            n5881;
wire      [7:0] n5882;
wire            n5883;
wire            n5884;
wire      [7:0] n5885;
wire            n5886;
wire            n5887;
wire      [7:0] n5888;
wire            n5889;
wire      [7:0] n589;
wire            n5890;
wire      [7:0] n5891;
wire            n5892;
wire            n5893;
wire      [7:0] n5894;
wire            n5895;
wire            n5896;
wire      [7:0] n5897;
wire            n5898;
wire            n5899;
wire      [2:0] n59;
wire      [7:0] n590;
wire      [7:0] n5900;
wire            n5901;
wire            n5902;
wire      [7:0] n5903;
wire            n5904;
wire            n5905;
wire      [7:0] n5906;
wire            n5907;
wire            n5908;
wire      [7:0] n5909;
wire      [7:0] n591;
wire            n5910;
wire            n5911;
wire      [7:0] n5912;
wire            n5913;
wire            n5914;
wire      [7:0] n5915;
wire            n5916;
wire            n5917;
wire      [7:0] n5918;
wire            n5919;
wire      [7:0] n592;
wire            n5920;
wire      [7:0] n5921;
wire            n5922;
wire            n5923;
wire      [7:0] n5924;
wire            n5925;
wire            n5926;
wire      [7:0] n5927;
wire            n5928;
wire            n5929;
wire      [7:0] n593;
wire      [7:0] n5930;
wire            n5931;
wire            n5932;
wire      [7:0] n5933;
wire            n5934;
wire            n5935;
wire      [7:0] n5936;
wire            n5937;
wire            n5938;
wire      [7:0] n5939;
wire      [7:0] n594;
wire            n5940;
wire            n5941;
wire      [7:0] n5942;
wire            n5943;
wire            n5944;
wire      [7:0] n5945;
wire            n5946;
wire            n5947;
wire      [7:0] n5948;
wire            n5949;
wire      [7:0] n595;
wire            n5950;
wire      [7:0] n5951;
wire            n5952;
wire            n5953;
wire      [7:0] n5954;
wire            n5955;
wire            n5956;
wire      [7:0] n5957;
wire            n5958;
wire            n5959;
wire      [7:0] n596;
wire      [7:0] n5960;
wire            n5961;
wire            n5962;
wire      [7:0] n5963;
wire            n5964;
wire            n5965;
wire      [7:0] n5966;
wire            n5967;
wire            n5968;
wire      [7:0] n5969;
wire      [7:0] n597;
wire            n5970;
wire            n5971;
wire      [7:0] n5972;
wire            n5973;
wire            n5974;
wire      [7:0] n5975;
wire            n5976;
wire            n5977;
wire      [7:0] n5978;
wire            n5979;
wire      [7:0] n598;
wire            n5980;
wire      [7:0] n5981;
wire            n5982;
wire            n5983;
wire      [7:0] n5984;
wire            n5985;
wire            n5986;
wire      [7:0] n5987;
wire            n5988;
wire            n5989;
wire      [7:0] n599;
wire      [7:0] n5990;
wire            n5991;
wire            n5992;
wire      [7:0] n5993;
wire            n5994;
wire            n5995;
wire      [7:0] n5996;
wire            n5997;
wire            n5998;
wire      [7:0] n5999;
wire      [2:0] n60;
wire      [7:0] n600;
wire            n6000;
wire            n6001;
wire      [7:0] n6002;
wire            n6003;
wire            n6004;
wire      [7:0] n6005;
wire            n6006;
wire            n6007;
wire      [7:0] n6008;
wire            n6009;
wire      [7:0] n601;
wire            n6010;
wire      [7:0] n6011;
wire            n6012;
wire            n6013;
wire      [7:0] n6014;
wire            n6015;
wire            n6016;
wire      [7:0] n6017;
wire            n6018;
wire            n6019;
wire      [7:0] n602;
wire      [7:0] n6020;
wire            n6021;
wire            n6022;
wire      [7:0] n6023;
wire            n6024;
wire            n6025;
wire      [7:0] n6026;
wire            n6027;
wire            n6028;
wire      [7:0] n6029;
wire      [7:0] n603;
wire            n6030;
wire            n6031;
wire      [7:0] n6032;
wire            n6033;
wire            n6034;
wire      [7:0] n6035;
wire            n6036;
wire            n6037;
wire      [7:0] n6038;
wire            n6039;
wire      [7:0] n604;
wire            n6040;
wire      [7:0] n6041;
wire            n6042;
wire            n6043;
wire      [7:0] n6044;
wire            n6045;
wire            n6046;
wire      [7:0] n6047;
wire            n6048;
wire            n6049;
wire      [7:0] n605;
wire      [7:0] n6050;
wire            n6051;
wire            n6052;
wire      [7:0] n6053;
wire            n6054;
wire            n6055;
wire      [7:0] n6056;
wire            n6057;
wire            n6058;
wire      [7:0] n6059;
wire      [7:0] n606;
wire            n6060;
wire            n6061;
wire      [7:0] n6062;
wire            n6063;
wire            n6064;
wire      [7:0] n6065;
wire            n6066;
wire            n6067;
wire      [7:0] n6068;
wire            n6069;
wire      [7:0] n607;
wire            n6070;
wire      [7:0] n6071;
wire            n6072;
wire            n6073;
wire      [7:0] n6074;
wire            n6075;
wire            n6076;
wire      [7:0] n6077;
wire            n6078;
wire            n6079;
wire      [7:0] n608;
wire      [7:0] n6080;
wire            n6081;
wire            n6082;
wire      [7:0] n6083;
wire            n6084;
wire            n6085;
wire      [7:0] n6086;
wire            n6087;
wire            n6088;
wire      [7:0] n6089;
wire      [7:0] n609;
wire            n6090;
wire            n6091;
wire      [7:0] n6092;
wire            n6093;
wire            n6094;
wire      [7:0] n6095;
wire            n6096;
wire            n6097;
wire      [7:0] n6098;
wire            n6099;
wire            n61;
wire      [7:0] n610;
wire            n6100;
wire      [7:0] n6101;
wire            n6102;
wire            n6103;
wire      [7:0] n6104;
wire            n6105;
wire            n6106;
wire      [7:0] n6107;
wire            n6108;
wire            n6109;
wire      [7:0] n611;
wire      [7:0] n6110;
wire            n6111;
wire            n6112;
wire      [7:0] n6113;
wire            n6114;
wire            n6115;
wire      [7:0] n6116;
wire            n6117;
wire            n6118;
wire      [7:0] n6119;
wire      [7:0] n612;
wire            n6120;
wire            n6121;
wire      [7:0] n6122;
wire            n6123;
wire            n6124;
wire      [7:0] n6125;
wire            n6126;
wire            n6127;
wire      [7:0] n6128;
wire            n6129;
wire      [7:0] n613;
wire            n6130;
wire      [7:0] n6131;
wire            n6132;
wire            n6133;
wire      [7:0] n6134;
wire            n6135;
wire            n6136;
wire      [7:0] n6137;
wire            n6138;
wire            n6139;
wire      [7:0] n614;
wire      [7:0] n6140;
wire            n6141;
wire            n6142;
wire      [7:0] n6143;
wire            n6144;
wire            n6145;
wire      [7:0] n6146;
wire            n6147;
wire            n6148;
wire      [7:0] n6149;
wire      [7:0] n615;
wire            n6150;
wire            n6151;
wire      [7:0] n6152;
wire            n6153;
wire            n6154;
wire      [7:0] n6155;
wire            n6156;
wire            n6157;
wire      [7:0] n6158;
wire            n6159;
wire      [7:0] n616;
wire            n6160;
wire      [7:0] n6161;
wire            n6162;
wire            n6163;
wire      [7:0] n6164;
wire            n6165;
wire            n6166;
wire      [7:0] n6167;
wire            n6168;
wire            n6169;
wire      [7:0] n617;
wire      [7:0] n6170;
wire            n6171;
wire            n6172;
wire      [7:0] n6173;
wire            n6174;
wire            n6175;
wire      [7:0] n6176;
wire            n6177;
wire            n6178;
wire      [7:0] n6179;
wire      [7:0] n618;
wire            n6180;
wire            n6181;
wire      [7:0] n6182;
wire            n6183;
wire            n6184;
wire      [7:0] n6185;
wire            n6186;
wire            n6187;
wire      [7:0] n6188;
wire            n6189;
wire      [7:0] n619;
wire            n6190;
wire      [7:0] n6191;
wire            n6192;
wire            n6193;
wire      [7:0] n6194;
wire            n6195;
wire            n6196;
wire      [7:0] n6197;
wire            n6198;
wire            n6199;
wire            n62;
wire      [7:0] n620;
wire      [7:0] n6200;
wire            n6201;
wire            n6202;
wire      [7:0] n6203;
wire            n6204;
wire            n6205;
wire      [7:0] n6206;
wire            n6207;
wire            n6208;
wire      [7:0] n6209;
wire      [7:0] n621;
wire            n6210;
wire            n6211;
wire      [7:0] n6212;
wire            n6213;
wire            n6214;
wire      [7:0] n6215;
wire            n6216;
wire            n6217;
wire      [7:0] n6218;
wire            n6219;
wire      [7:0] n622;
wire            n6220;
wire      [7:0] n6221;
wire            n6222;
wire            n6223;
wire      [7:0] n6224;
wire            n6225;
wire            n6226;
wire      [7:0] n6227;
wire            n6228;
wire            n6229;
wire      [7:0] n623;
wire      [7:0] n6230;
wire            n6231;
wire            n6232;
wire      [7:0] n6233;
wire            n6234;
wire            n6235;
wire      [7:0] n6236;
wire            n6237;
wire            n6238;
wire      [7:0] n6239;
wire      [7:0] n624;
wire            n6240;
wire            n6241;
wire      [7:0] n6242;
wire            n6243;
wire            n6244;
wire      [7:0] n6245;
wire            n6246;
wire            n6247;
wire      [7:0] n6248;
wire            n6249;
wire      [7:0] n625;
wire            n6250;
wire      [7:0] n6251;
wire            n6252;
wire            n6253;
wire      [7:0] n6254;
wire            n6255;
wire            n6256;
wire      [7:0] n6257;
wire            n6258;
wire            n6259;
wire      [7:0] n626;
wire      [7:0] n6260;
wire            n6261;
wire            n6262;
wire      [7:0] n6263;
wire            n6264;
wire            n6265;
wire      [7:0] n6266;
wire            n6267;
wire            n6268;
wire      [7:0] n6269;
wire      [7:0] n627;
wire            n6270;
wire            n6271;
wire      [7:0] n6272;
wire            n6273;
wire            n6274;
wire      [7:0] n6275;
wire            n6276;
wire            n6277;
wire      [7:0] n6278;
wire            n6279;
wire      [7:0] n628;
wire            n6280;
wire      [7:0] n6281;
wire            n6282;
wire            n6283;
wire      [7:0] n6284;
wire            n6285;
wire            n6286;
wire      [7:0] n6287;
wire            n6288;
wire            n6289;
wire      [7:0] n629;
wire      [7:0] n6290;
wire            n6291;
wire            n6292;
wire      [7:0] n6293;
wire            n6294;
wire            n6295;
wire      [7:0] n6296;
wire            n6297;
wire            n6298;
wire      [7:0] n6299;
wire      [3:0] n63;
wire      [7:0] n630;
wire            n6300;
wire            n6301;
wire      [7:0] n6302;
wire            n6303;
wire            n6304;
wire      [7:0] n6305;
wire            n6306;
wire            n6307;
wire      [7:0] n6308;
wire            n6309;
wire      [7:0] n631;
wire            n6310;
wire      [7:0] n6311;
wire            n6312;
wire            n6313;
wire      [7:0] n6314;
wire            n6315;
wire            n6316;
wire      [7:0] n6317;
wire            n6318;
wire            n6319;
wire      [7:0] n632;
wire      [7:0] n6320;
wire            n6321;
wire            n6322;
wire      [7:0] n6323;
wire            n6324;
wire            n6325;
wire      [7:0] n6326;
wire            n6327;
wire            n6328;
wire            n6329;
wire      [7:0] n633;
wire            n6330;
wire            n6331;
wire      [7:0] n6332;
wire            n6333;
wire            n6334;
wire            n6335;
wire            n6336;
wire            n6337;
wire      [7:0] n6338;
wire            n6339;
wire      [7:0] n634;
wire            n6340;
wire            n6341;
wire            n6342;
wire            n6343;
wire      [7:0] n6344;
wire            n6345;
wire            n6346;
wire            n6347;
wire            n6348;
wire            n6349;
wire      [7:0] n635;
wire      [7:0] n6350;
wire            n6351;
wire            n6352;
wire            n6353;
wire            n6354;
wire            n6355;
wire      [7:0] n6356;
wire            n6357;
wire            n6358;
wire            n6359;
wire      [7:0] n636;
wire            n6360;
wire            n6361;
wire      [7:0] n6362;
wire            n6363;
wire            n6364;
wire            n6365;
wire            n6366;
wire            n6367;
wire      [7:0] n6368;
wire            n6369;
wire      [7:0] n637;
wire            n6370;
wire            n6371;
wire            n6372;
wire            n6373;
wire      [7:0] n6374;
wire            n6375;
wire            n6376;
wire            n6377;
wire            n6378;
wire            n6379;
wire      [7:0] n638;
wire      [7:0] n6380;
wire            n6381;
wire            n6382;
wire            n6383;
wire            n6384;
wire            n6385;
wire      [7:0] n6386;
wire            n6387;
wire            n6388;
wire            n6389;
wire      [7:0] n639;
wire            n6390;
wire            n6391;
wire      [7:0] n6392;
wire            n6393;
wire            n6394;
wire            n6395;
wire            n6396;
wire            n6397;
wire      [7:0] n6398;
wire            n6399;
wire      [4:0] n64;
wire      [7:0] n640;
wire            n6400;
wire            n6401;
wire            n6402;
wire            n6403;
wire      [7:0] n6404;
wire            n6405;
wire            n6406;
wire            n6407;
wire            n6408;
wire            n6409;
wire      [7:0] n641;
wire      [7:0] n6410;
wire            n6411;
wire            n6412;
wire            n6413;
wire            n6414;
wire            n6415;
wire      [7:0] n6416;
wire            n6417;
wire            n6418;
wire            n6419;
wire      [7:0] n642;
wire            n6420;
wire            n6421;
wire      [7:0] n6422;
wire            n6423;
wire            n6424;
wire            n6425;
wire            n6426;
wire            n6427;
wire      [7:0] n6428;
wire            n6429;
wire      [7:0] n643;
wire            n6430;
wire            n6431;
wire            n6432;
wire            n6433;
wire      [7:0] n6434;
wire            n6435;
wire            n6436;
wire            n6437;
wire            n6438;
wire            n6439;
wire      [7:0] n644;
wire      [7:0] n6440;
wire            n6441;
wire            n6442;
wire            n6443;
wire            n6444;
wire            n6445;
wire      [7:0] n6446;
wire            n6447;
wire            n6448;
wire            n6449;
wire      [7:0] n645;
wire            n6450;
wire            n6451;
wire      [7:0] n6452;
wire            n6453;
wire            n6454;
wire            n6455;
wire            n6456;
wire            n6457;
wire      [7:0] n6458;
wire            n6459;
wire      [7:0] n646;
wire            n6460;
wire            n6461;
wire            n6462;
wire            n6463;
wire      [7:0] n6464;
wire            n6465;
wire            n6466;
wire            n6467;
wire            n6468;
wire            n6469;
wire      [7:0] n647;
wire      [7:0] n6470;
wire            n6471;
wire            n6472;
wire            n6473;
wire            n6474;
wire            n6475;
wire      [7:0] n6476;
wire            n6477;
wire            n6478;
wire            n6479;
wire      [7:0] n648;
wire            n6480;
wire            n6481;
wire      [7:0] n6482;
wire            n6483;
wire            n6484;
wire            n6485;
wire            n6486;
wire            n6487;
wire      [7:0] n6488;
wire            n6489;
wire      [7:0] n649;
wire            n6490;
wire            n6491;
wire            n6492;
wire            n6493;
wire      [7:0] n6494;
wire            n6495;
wire            n6496;
wire            n6497;
wire            n6498;
wire            n6499;
wire      [7:0] n65;
wire      [7:0] n650;
wire      [7:0] n6500;
wire            n6501;
wire            n6502;
wire            n6503;
wire            n6504;
wire            n6505;
wire      [7:0] n6506;
wire            n6507;
wire            n6508;
wire            n6509;
wire      [7:0] n651;
wire            n6510;
wire            n6511;
wire      [7:0] n6512;
wire            n6513;
wire            n6514;
wire            n6515;
wire            n6516;
wire            n6517;
wire      [7:0] n6518;
wire            n6519;
wire      [7:0] n652;
wire            n6520;
wire            n6521;
wire            n6522;
wire            n6523;
wire      [7:0] n6524;
wire            n6525;
wire            n6526;
wire            n6527;
wire            n6528;
wire            n6529;
wire      [7:0] n653;
wire      [7:0] n6530;
wire            n6531;
wire            n6532;
wire            n6533;
wire            n6534;
wire            n6535;
wire      [7:0] n6536;
wire            n6537;
wire            n6538;
wire            n6539;
wire      [7:0] n654;
wire            n6540;
wire            n6541;
wire      [7:0] n6542;
wire            n6543;
wire            n6544;
wire            n6545;
wire            n6546;
wire            n6547;
wire      [7:0] n6548;
wire            n6549;
wire      [7:0] n655;
wire            n6550;
wire            n6551;
wire            n6552;
wire            n6553;
wire      [7:0] n6554;
wire            n6555;
wire            n6556;
wire            n6557;
wire            n6558;
wire            n6559;
wire      [7:0] n656;
wire      [7:0] n6560;
wire            n6561;
wire            n6562;
wire            n6563;
wire            n6564;
wire            n6565;
wire      [7:0] n6566;
wire            n6567;
wire            n6568;
wire            n6569;
wire      [7:0] n657;
wire            n6570;
wire            n6571;
wire      [7:0] n6572;
wire            n6573;
wire            n6574;
wire            n6575;
wire            n6576;
wire            n6577;
wire      [7:0] n6578;
wire            n6579;
wire      [7:0] n658;
wire            n6580;
wire            n6581;
wire            n6582;
wire            n6583;
wire      [7:0] n6584;
wire            n6585;
wire            n6586;
wire            n6587;
wire            n6588;
wire            n6589;
wire      [7:0] n659;
wire      [7:0] n6590;
wire            n6591;
wire            n6592;
wire            n6593;
wire            n6594;
wire            n6595;
wire      [7:0] n6596;
wire            n6597;
wire            n6598;
wire            n6599;
wire      [3:0] n66;
wire      [7:0] n660;
wire            n6600;
wire            n6601;
wire      [7:0] n6602;
wire            n6603;
wire            n6604;
wire            n6605;
wire            n6606;
wire            n6607;
wire      [7:0] n6608;
wire            n6609;
wire      [7:0] n661;
wire            n6610;
wire            n6611;
wire            n6612;
wire            n6613;
wire      [7:0] n6614;
wire            n6615;
wire            n6616;
wire            n6617;
wire            n6618;
wire            n6619;
wire      [7:0] n662;
wire      [7:0] n6620;
wire            n6621;
wire            n6622;
wire            n6623;
wire            n6624;
wire            n6625;
wire      [7:0] n6626;
wire            n6627;
wire            n6628;
wire            n6629;
wire      [7:0] n663;
wire            n6630;
wire            n6631;
wire      [7:0] n6632;
wire            n6633;
wire            n6634;
wire            n6635;
wire            n6636;
wire            n6637;
wire      [7:0] n6638;
wire            n6639;
wire      [7:0] n664;
wire            n6640;
wire            n6641;
wire            n6642;
wire            n6643;
wire      [7:0] n6644;
wire            n6645;
wire            n6646;
wire            n6647;
wire            n6648;
wire            n6649;
wire      [7:0] n665;
wire      [7:0] n6650;
wire            n6651;
wire            n6652;
wire            n6653;
wire            n6654;
wire            n6655;
wire      [7:0] n6656;
wire            n6657;
wire            n6658;
wire            n6659;
wire      [7:0] n666;
wire            n6660;
wire            n6661;
wire      [7:0] n6662;
wire            n6663;
wire            n6664;
wire            n6665;
wire            n6666;
wire            n6667;
wire      [7:0] n6668;
wire            n6669;
wire      [7:0] n667;
wire            n6670;
wire            n6671;
wire            n6672;
wire            n6673;
wire      [7:0] n6674;
wire            n6675;
wire            n6676;
wire            n6677;
wire            n6678;
wire            n6679;
wire      [7:0] n668;
wire      [7:0] n6680;
wire            n6681;
wire            n6682;
wire            n6683;
wire            n6684;
wire            n6685;
wire      [7:0] n6686;
wire            n6687;
wire            n6688;
wire            n6689;
wire      [7:0] n669;
wire            n6690;
wire            n6691;
wire      [7:0] n6692;
wire            n6693;
wire            n6694;
wire            n6695;
wire            n6696;
wire            n6697;
wire      [7:0] n6698;
wire            n6699;
wire      [7:0] n67;
wire      [7:0] n670;
wire            n6700;
wire            n6701;
wire            n6702;
wire            n6703;
wire      [7:0] n6704;
wire            n6705;
wire            n6706;
wire            n6707;
wire            n6708;
wire            n6709;
wire      [7:0] n671;
wire      [7:0] n6710;
wire            n6711;
wire            n6712;
wire            n6713;
wire            n6714;
wire            n6715;
wire      [7:0] n6716;
wire            n6717;
wire            n6718;
wire            n6719;
wire      [7:0] n672;
wire            n6720;
wire            n6721;
wire      [7:0] n6722;
wire            n6723;
wire            n6724;
wire            n6725;
wire            n6726;
wire            n6727;
wire      [7:0] n6728;
wire            n6729;
wire      [7:0] n673;
wire            n6730;
wire            n6731;
wire            n6732;
wire            n6733;
wire      [7:0] n6734;
wire            n6735;
wire            n6736;
wire            n6737;
wire            n6738;
wire            n6739;
wire      [7:0] n674;
wire      [7:0] n6740;
wire            n6741;
wire            n6742;
wire            n6743;
wire            n6744;
wire            n6745;
wire      [7:0] n6746;
wire            n6747;
wire            n6748;
wire            n6749;
wire      [7:0] n675;
wire            n6750;
wire            n6751;
wire      [7:0] n6752;
wire            n6753;
wire            n6754;
wire            n6755;
wire            n6756;
wire            n6757;
wire      [7:0] n6758;
wire            n6759;
wire      [7:0] n676;
wire            n6760;
wire            n6761;
wire            n6762;
wire            n6763;
wire      [7:0] n6764;
wire            n6765;
wire            n6766;
wire            n6767;
wire            n6768;
wire            n6769;
wire      [7:0] n677;
wire      [7:0] n6770;
wire            n6771;
wire            n6772;
wire            n6773;
wire            n6774;
wire            n6775;
wire      [7:0] n6776;
wire            n6777;
wire            n6778;
wire            n6779;
wire      [7:0] n678;
wire            n6780;
wire            n6781;
wire      [7:0] n6782;
wire            n6783;
wire            n6784;
wire            n6785;
wire            n6786;
wire            n6787;
wire      [7:0] n6788;
wire            n6789;
wire      [7:0] n679;
wire            n6790;
wire            n6791;
wire            n6792;
wire            n6793;
wire      [7:0] n6794;
wire            n6795;
wire            n6796;
wire            n6797;
wire            n6798;
wire            n6799;
wire      [7:0] n68;
wire      [7:0] n680;
wire      [7:0] n6800;
wire            n6801;
wire            n6802;
wire            n6803;
wire            n6804;
wire            n6805;
wire      [7:0] n6806;
wire            n6807;
wire            n6808;
wire            n6809;
wire      [7:0] n681;
wire            n6810;
wire            n6811;
wire      [7:0] n6812;
wire            n6813;
wire            n6814;
wire            n6815;
wire            n6816;
wire            n6817;
wire      [7:0] n6818;
wire            n6819;
wire      [7:0] n682;
wire            n6820;
wire            n6821;
wire            n6822;
wire            n6823;
wire      [7:0] n6824;
wire            n6825;
wire            n6826;
wire            n6827;
wire            n6828;
wire            n6829;
wire      [7:0] n683;
wire      [7:0] n6830;
wire            n6831;
wire            n6832;
wire            n6833;
wire            n6834;
wire            n6835;
wire      [7:0] n6836;
wire            n6837;
wire            n6838;
wire            n6839;
wire      [7:0] n684;
wire            n6840;
wire            n6841;
wire      [7:0] n6842;
wire            n6843;
wire            n6844;
wire            n6845;
wire            n6846;
wire            n6847;
wire      [7:0] n6848;
wire            n6849;
wire      [7:0] n685;
wire            n6850;
wire            n6851;
wire            n6852;
wire            n6853;
wire      [7:0] n6854;
wire            n6855;
wire            n6856;
wire            n6857;
wire            n6858;
wire            n6859;
wire      [7:0] n686;
wire      [7:0] n6860;
wire            n6861;
wire            n6862;
wire            n6863;
wire            n6864;
wire            n6865;
wire      [7:0] n6866;
wire            n6867;
wire            n6868;
wire            n6869;
wire      [7:0] n687;
wire            n6870;
wire            n6871;
wire      [7:0] n6872;
wire            n6873;
wire            n6874;
wire            n6875;
wire            n6876;
wire            n6877;
wire      [7:0] n6878;
wire            n6879;
wire      [7:0] n688;
wire            n6880;
wire            n6881;
wire            n6882;
wire            n6883;
wire      [7:0] n6884;
wire            n6885;
wire            n6886;
wire            n6887;
wire            n6888;
wire            n6889;
wire      [7:0] n689;
wire      [7:0] n6890;
wire            n6891;
wire            n6892;
wire            n6893;
wire            n6894;
wire            n6895;
wire      [7:0] n6896;
wire            n6897;
wire            n6898;
wire            n6899;
wire      [7:0] n690;
wire            n6900;
wire            n6901;
wire      [7:0] n6902;
wire            n6903;
wire            n6904;
wire            n6905;
wire            n6906;
wire            n6907;
wire      [7:0] n6908;
wire            n6909;
wire      [7:0] n691;
wire            n6910;
wire            n6911;
wire            n6912;
wire            n6913;
wire      [7:0] n6914;
wire            n6915;
wire            n6916;
wire            n6917;
wire            n6918;
wire            n6919;
wire      [7:0] n692;
wire      [7:0] n6920;
wire            n6921;
wire            n6922;
wire            n6923;
wire            n6924;
wire            n6925;
wire      [7:0] n6926;
wire            n6927;
wire            n6928;
wire            n6929;
wire      [7:0] n693;
wire            n6930;
wire            n6931;
wire      [7:0] n6932;
wire            n6933;
wire            n6934;
wire            n6935;
wire            n6936;
wire            n6937;
wire      [7:0] n6938;
wire            n6939;
wire      [7:0] n694;
wire            n6940;
wire            n6941;
wire            n6942;
wire            n6943;
wire      [7:0] n6944;
wire            n6945;
wire            n6946;
wire            n6947;
wire            n6948;
wire            n6949;
wire      [7:0] n695;
wire      [7:0] n6950;
wire            n6951;
wire            n6952;
wire            n6953;
wire            n6954;
wire            n6955;
wire      [7:0] n6956;
wire            n6957;
wire            n6958;
wire            n6959;
wire      [7:0] n696;
wire            n6960;
wire            n6961;
wire      [7:0] n6962;
wire            n6963;
wire            n6964;
wire            n6965;
wire            n6966;
wire            n6967;
wire      [7:0] n6968;
wire            n6969;
wire      [7:0] n697;
wire            n6970;
wire            n6971;
wire            n6972;
wire            n6973;
wire      [7:0] n6974;
wire            n6975;
wire            n6976;
wire            n6977;
wire            n6978;
wire            n6979;
wire      [7:0] n698;
wire      [7:0] n6980;
wire            n6981;
wire            n6982;
wire            n6983;
wire            n6984;
wire            n6985;
wire      [7:0] n6986;
wire            n6987;
wire            n6988;
wire            n6989;
wire      [7:0] n699;
wire            n6990;
wire            n6991;
wire      [7:0] n6992;
wire            n6993;
wire            n6994;
wire            n6995;
wire            n6996;
wire            n6997;
wire      [7:0] n6998;
wire            n6999;
wire            n7;
wire            n70;
wire      [7:0] n700;
wire            n7000;
wire            n7001;
wire            n7002;
wire            n7003;
wire      [7:0] n7004;
wire            n7005;
wire            n7006;
wire            n7007;
wire            n7008;
wire            n7009;
wire      [7:0] n701;
wire      [7:0] n7010;
wire            n7011;
wire            n7012;
wire            n7013;
wire            n7014;
wire            n7015;
wire      [7:0] n7016;
wire            n7017;
wire            n7018;
wire            n7019;
wire      [7:0] n702;
wire            n7020;
wire            n7021;
wire      [7:0] n7022;
wire            n7023;
wire            n7024;
wire            n7025;
wire            n7026;
wire            n7027;
wire      [7:0] n7028;
wire            n7029;
wire      [7:0] n703;
wire            n7030;
wire            n7031;
wire            n7032;
wire            n7033;
wire      [7:0] n7034;
wire            n7035;
wire            n7036;
wire            n7037;
wire            n7038;
wire            n7039;
wire      [7:0] n704;
wire      [7:0] n7040;
wire            n7041;
wire            n7042;
wire            n7043;
wire            n7044;
wire            n7045;
wire      [7:0] n7046;
wire            n7047;
wire            n7048;
wire            n7049;
wire      [7:0] n705;
wire            n7050;
wire            n7051;
wire      [7:0] n7052;
wire            n7053;
wire            n7054;
wire            n7055;
wire            n7056;
wire            n7057;
wire      [7:0] n7058;
wire            n7059;
wire      [7:0] n706;
wire            n7060;
wire            n7061;
wire            n7062;
wire            n7063;
wire      [7:0] n7064;
wire            n7065;
wire            n7066;
wire            n7067;
wire            n7068;
wire            n7069;
wire      [7:0] n707;
wire      [7:0] n7070;
wire            n7071;
wire            n7072;
wire            n7073;
wire            n7074;
wire            n7075;
wire      [7:0] n7076;
wire            n7077;
wire            n7078;
wire            n7079;
wire      [7:0] n708;
wire            n7080;
wire            n7081;
wire      [7:0] n7082;
wire            n7083;
wire            n7084;
wire            n7085;
wire            n7086;
wire            n7087;
wire      [7:0] n7088;
wire            n7089;
wire      [7:0] n709;
wire            n7090;
wire            n7091;
wire            n7092;
wire            n7093;
wire      [7:0] n7094;
wire            n7095;
wire            n7096;
wire            n7097;
wire            n7098;
wire            n7099;
wire      [7:0] n710;
wire      [7:0] n7100;
wire            n7101;
wire            n7102;
wire            n7103;
wire            n7104;
wire            n7105;
wire      [7:0] n7106;
wire            n7107;
wire            n7108;
wire            n7109;
wire      [7:0] n711;
wire            n7110;
wire            n7111;
wire      [7:0] n7112;
wire            n7113;
wire            n7114;
wire            n7115;
wire            n7116;
wire            n7117;
wire      [7:0] n7118;
wire            n7119;
wire      [7:0] n712;
wire            n7120;
wire            n7121;
wire            n7122;
wire            n7123;
wire      [7:0] n7124;
wire            n7125;
wire            n7126;
wire            n7127;
wire            n7128;
wire            n7129;
wire      [7:0] n713;
wire      [7:0] n7130;
wire            n7131;
wire            n7132;
wire            n7133;
wire            n7134;
wire            n7135;
wire      [7:0] n7136;
wire            n7137;
wire            n7138;
wire            n7139;
wire      [7:0] n714;
wire            n7140;
wire            n7141;
wire      [7:0] n7142;
wire            n7143;
wire            n7144;
wire            n7145;
wire            n7146;
wire            n7147;
wire      [7:0] n7148;
wire            n7149;
wire      [7:0] n715;
wire            n7150;
wire            n7151;
wire            n7152;
wire            n7153;
wire      [7:0] n7154;
wire            n7155;
wire            n7156;
wire            n7157;
wire            n7158;
wire            n7159;
wire      [7:0] n716;
wire      [7:0] n7160;
wire            n7161;
wire            n7162;
wire            n7163;
wire            n7164;
wire            n7165;
wire      [7:0] n7166;
wire            n7167;
wire            n7168;
wire            n7169;
wire      [7:0] n717;
wire            n7170;
wire            n7171;
wire      [7:0] n7172;
wire            n7173;
wire            n7174;
wire            n7175;
wire            n7176;
wire            n7177;
wire      [7:0] n7178;
wire            n7179;
wire      [7:0] n718;
wire            n7180;
wire            n7181;
wire            n7182;
wire            n7183;
wire      [7:0] n7184;
wire            n7185;
wire            n7186;
wire            n7187;
wire            n7188;
wire            n7189;
wire      [7:0] n719;
wire      [7:0] n7190;
wire            n7191;
wire            n7192;
wire            n7193;
wire            n7194;
wire            n7195;
wire      [7:0] n7196;
wire            n7197;
wire            n7198;
wire            n7199;
wire            n72;
wire      [7:0] n720;
wire            n7200;
wire            n7201;
wire      [7:0] n7202;
wire            n7203;
wire            n7204;
wire            n7205;
wire            n7206;
wire            n7207;
wire      [7:0] n7208;
wire            n7209;
wire      [7:0] n721;
wire            n7210;
wire            n7211;
wire            n7212;
wire            n7213;
wire      [7:0] n7214;
wire            n7215;
wire            n7216;
wire            n7217;
wire            n7218;
wire            n7219;
wire      [7:0] n722;
wire      [7:0] n7220;
wire            n7221;
wire            n7222;
wire            n7223;
wire            n7224;
wire            n7225;
wire      [7:0] n7226;
wire            n7227;
wire            n7228;
wire            n7229;
wire      [7:0] n723;
wire            n7230;
wire            n7231;
wire      [7:0] n7232;
wire            n7233;
wire            n7234;
wire            n7235;
wire            n7236;
wire            n7237;
wire      [7:0] n7238;
wire            n7239;
wire      [7:0] n724;
wire            n7240;
wire            n7241;
wire            n7242;
wire            n7243;
wire      [7:0] n7244;
wire            n7245;
wire            n7246;
wire            n7247;
wire            n7248;
wire            n7249;
wire      [7:0] n725;
wire      [7:0] n7250;
wire            n7251;
wire            n7252;
wire            n7253;
wire            n7254;
wire            n7255;
wire      [7:0] n7256;
wire            n7257;
wire            n7258;
wire            n7259;
wire      [7:0] n726;
wire            n7260;
wire            n7261;
wire      [7:0] n7262;
wire            n7263;
wire            n7264;
wire            n7265;
wire            n7266;
wire            n7267;
wire      [7:0] n7268;
wire            n7269;
wire      [7:0] n727;
wire            n7270;
wire            n7271;
wire            n7272;
wire            n7273;
wire      [7:0] n7274;
wire            n7275;
wire            n7276;
wire            n7277;
wire            n7278;
wire            n7279;
wire      [7:0] n728;
wire      [7:0] n7280;
wire            n7281;
wire            n7282;
wire            n7283;
wire            n7284;
wire            n7285;
wire      [7:0] n7286;
wire            n7287;
wire            n7288;
wire            n7289;
wire      [7:0] n729;
wire            n7290;
wire            n7291;
wire      [7:0] n7292;
wire            n7293;
wire            n7294;
wire            n7295;
wire            n7296;
wire            n7297;
wire      [7:0] n7298;
wire            n7299;
wire      [7:0] n730;
wire            n7300;
wire            n7301;
wire            n7302;
wire            n7303;
wire      [7:0] n7304;
wire            n7305;
wire            n7306;
wire            n7307;
wire            n7308;
wire            n7309;
wire      [7:0] n731;
wire      [7:0] n7310;
wire            n7311;
wire            n7312;
wire            n7313;
wire            n7314;
wire            n7315;
wire      [7:0] n7316;
wire            n7317;
wire            n7318;
wire            n7319;
wire      [7:0] n732;
wire            n7320;
wire            n7321;
wire      [7:0] n7322;
wire            n7323;
wire            n7324;
wire            n7325;
wire            n7326;
wire            n7327;
wire      [7:0] n7328;
wire            n7329;
wire      [7:0] n733;
wire            n7330;
wire            n7331;
wire            n7332;
wire            n7333;
wire      [7:0] n7334;
wire            n7335;
wire            n7336;
wire            n7337;
wire            n7338;
wire            n7339;
wire      [7:0] n734;
wire      [7:0] n7340;
wire            n7341;
wire            n7342;
wire            n7343;
wire            n7344;
wire            n7345;
wire      [7:0] n7346;
wire            n7347;
wire            n7348;
wire            n7349;
wire      [7:0] n735;
wire            n7350;
wire            n7351;
wire      [7:0] n7352;
wire            n7353;
wire            n7354;
wire            n7355;
wire            n7356;
wire            n7357;
wire      [7:0] n7358;
wire            n7359;
wire      [7:0] n736;
wire            n7360;
wire            n7361;
wire            n7362;
wire            n7363;
wire      [7:0] n7364;
wire            n7365;
wire            n7366;
wire            n7367;
wire            n7368;
wire            n7369;
wire      [7:0] n737;
wire      [7:0] n7370;
wire            n7371;
wire            n7372;
wire            n7373;
wire            n7374;
wire            n7375;
wire      [7:0] n7376;
wire            n7377;
wire            n7378;
wire            n7379;
wire      [7:0] n738;
wire            n7380;
wire            n7381;
wire      [7:0] n7382;
wire            n7383;
wire            n7384;
wire            n7385;
wire            n7386;
wire            n7387;
wire      [7:0] n7388;
wire            n7389;
wire      [7:0] n739;
wire            n7390;
wire            n7391;
wire            n7392;
wire            n7393;
wire      [7:0] n7394;
wire            n7395;
wire            n7396;
wire            n7397;
wire            n7398;
wire            n7399;
wire            n74;
wire      [7:0] n740;
wire      [7:0] n7400;
wire            n7401;
wire            n7402;
wire            n7403;
wire            n7404;
wire            n7405;
wire      [7:0] n7406;
wire            n7407;
wire            n7408;
wire            n7409;
wire      [7:0] n741;
wire            n7410;
wire            n7411;
wire      [7:0] n7412;
wire            n7413;
wire            n7414;
wire            n7415;
wire            n7416;
wire            n7417;
wire      [7:0] n7418;
wire            n7419;
wire      [7:0] n742;
wire            n7420;
wire            n7421;
wire            n7422;
wire            n7423;
wire      [7:0] n7424;
wire            n7425;
wire            n7426;
wire            n7427;
wire            n7428;
wire            n7429;
wire      [7:0] n743;
wire      [7:0] n7430;
wire            n7431;
wire            n7432;
wire            n7433;
wire            n7434;
wire            n7435;
wire      [7:0] n7436;
wire            n7437;
wire            n7438;
wire            n7439;
wire      [7:0] n744;
wire            n7440;
wire            n7441;
wire      [7:0] n7442;
wire            n7443;
wire            n7444;
wire            n7445;
wire            n7446;
wire            n7447;
wire      [7:0] n7448;
wire            n7449;
wire      [7:0] n745;
wire            n7450;
wire            n7451;
wire            n7452;
wire            n7453;
wire      [7:0] n7454;
wire            n7455;
wire            n7456;
wire            n7457;
wire            n7458;
wire            n7459;
wire      [7:0] n746;
wire      [7:0] n7460;
wire            n7461;
wire            n7462;
wire            n7463;
wire            n7464;
wire            n7465;
wire      [7:0] n7466;
wire            n7467;
wire            n7468;
wire            n7469;
wire      [7:0] n747;
wire            n7470;
wire            n7471;
wire      [7:0] n7472;
wire            n7473;
wire            n7474;
wire            n7475;
wire            n7476;
wire            n7477;
wire      [7:0] n7478;
wire            n7479;
wire      [7:0] n748;
wire            n7480;
wire            n7481;
wire            n7482;
wire            n7483;
wire      [7:0] n7484;
wire            n7485;
wire            n7486;
wire            n7487;
wire            n7488;
wire            n7489;
wire      [7:0] n749;
wire      [7:0] n7490;
wire            n7491;
wire            n7492;
wire            n7493;
wire            n7494;
wire            n7495;
wire      [7:0] n7496;
wire            n7497;
wire            n7498;
wire            n7499;
wire      [7:0] n750;
wire            n7500;
wire            n7501;
wire      [7:0] n7502;
wire            n7503;
wire            n7504;
wire            n7505;
wire            n7506;
wire            n7507;
wire      [7:0] n7508;
wire            n7509;
wire      [7:0] n751;
wire            n7510;
wire            n7511;
wire            n7512;
wire            n7513;
wire      [7:0] n7514;
wire            n7515;
wire            n7516;
wire            n7517;
wire            n7518;
wire            n7519;
wire      [7:0] n752;
wire      [7:0] n7520;
wire            n7521;
wire            n7522;
wire            n7523;
wire            n7524;
wire            n7525;
wire      [7:0] n7526;
wire            n7527;
wire            n7528;
wire            n7529;
wire      [7:0] n753;
wire            n7530;
wire            n7531;
wire      [7:0] n7532;
wire            n7533;
wire            n7534;
wire            n7535;
wire            n7536;
wire            n7537;
wire      [7:0] n7538;
wire            n7539;
wire      [7:0] n754;
wire            n7540;
wire            n7541;
wire            n7542;
wire            n7543;
wire      [7:0] n7544;
wire            n7545;
wire            n7546;
wire            n7547;
wire            n7548;
wire            n7549;
wire      [7:0] n755;
wire      [7:0] n7550;
wire            n7551;
wire            n7552;
wire            n7553;
wire            n7554;
wire            n7555;
wire      [7:0] n7556;
wire            n7557;
wire            n7558;
wire            n7559;
wire      [7:0] n756;
wire            n7560;
wire            n7561;
wire      [7:0] n7562;
wire            n7563;
wire            n7564;
wire            n7565;
wire            n7566;
wire            n7567;
wire      [7:0] n7568;
wire            n7569;
wire      [7:0] n757;
wire            n7570;
wire            n7571;
wire            n7572;
wire            n7573;
wire      [7:0] n7574;
wire            n7575;
wire            n7576;
wire            n7577;
wire            n7578;
wire            n7579;
wire      [7:0] n758;
wire      [7:0] n7580;
wire            n7581;
wire            n7582;
wire            n7583;
wire            n7584;
wire            n7585;
wire      [7:0] n7586;
wire            n7587;
wire            n7588;
wire            n7589;
wire      [7:0] n759;
wire            n7590;
wire            n7591;
wire      [7:0] n7592;
wire            n7593;
wire            n7594;
wire            n7595;
wire            n7596;
wire            n7597;
wire      [7:0] n7598;
wire            n7599;
wire            n76;
wire      [7:0] n760;
wire            n7600;
wire            n7601;
wire            n7602;
wire            n7603;
wire      [7:0] n7604;
wire            n7605;
wire            n7606;
wire            n7607;
wire            n7608;
wire            n7609;
wire      [7:0] n761;
wire      [7:0] n7610;
wire            n7611;
wire            n7612;
wire            n7613;
wire            n7614;
wire            n7615;
wire      [7:0] n7616;
wire            n7617;
wire            n7618;
wire            n7619;
wire      [7:0] n762;
wire            n7620;
wire            n7621;
wire      [7:0] n7622;
wire            n7623;
wire            n7624;
wire            n7625;
wire            n7626;
wire            n7627;
wire      [7:0] n7628;
wire            n7629;
wire      [7:0] n763;
wire            n7630;
wire            n7631;
wire            n7632;
wire            n7633;
wire      [7:0] n7634;
wire            n7635;
wire            n7636;
wire            n7637;
wire            n7638;
wire            n7639;
wire      [7:0] n764;
wire      [7:0] n7640;
wire            n7641;
wire            n7642;
wire            n7643;
wire            n7644;
wire            n7645;
wire      [7:0] n7646;
wire            n7647;
wire            n7648;
wire            n7649;
wire      [7:0] n765;
wire            n7650;
wire            n7651;
wire      [7:0] n7652;
wire            n7653;
wire            n7654;
wire            n7655;
wire            n7656;
wire            n7657;
wire      [7:0] n7658;
wire            n7659;
wire      [7:0] n766;
wire            n7660;
wire            n7661;
wire            n7662;
wire            n7663;
wire      [7:0] n7664;
wire            n7665;
wire            n7666;
wire            n7667;
wire            n7668;
wire            n7669;
wire      [7:0] n767;
wire      [7:0] n7670;
wire            n7671;
wire            n7672;
wire            n7673;
wire            n7674;
wire            n7675;
wire      [7:0] n7676;
wire            n7677;
wire            n7678;
wire            n7679;
wire      [7:0] n768;
wire            n7680;
wire            n7681;
wire      [7:0] n7682;
wire            n7683;
wire            n7684;
wire            n7685;
wire            n7686;
wire            n7687;
wire      [7:0] n7688;
wire            n7689;
wire      [7:0] n769;
wire            n7690;
wire            n7691;
wire            n7692;
wire            n7693;
wire      [7:0] n7694;
wire            n7695;
wire            n7696;
wire            n7697;
wire            n7698;
wire            n7699;
wire      [7:0] n770;
wire      [7:0] n7700;
wire            n7701;
wire            n7702;
wire            n7703;
wire            n7704;
wire            n7705;
wire      [7:0] n7706;
wire            n7707;
wire            n7708;
wire            n7709;
wire      [7:0] n771;
wire            n7710;
wire            n7711;
wire      [7:0] n7712;
wire            n7713;
wire            n7714;
wire            n7715;
wire            n7716;
wire            n7717;
wire      [7:0] n7718;
wire            n7719;
wire      [7:0] n772;
wire            n7720;
wire            n7721;
wire            n7722;
wire            n7723;
wire      [7:0] n7724;
wire            n7725;
wire            n7726;
wire            n7727;
wire            n7728;
wire            n7729;
wire      [7:0] n773;
wire      [7:0] n7730;
wire            n7731;
wire            n7732;
wire            n7733;
wire            n7734;
wire            n7735;
wire      [7:0] n7736;
wire            n7737;
wire            n7738;
wire            n7739;
wire      [7:0] n774;
wire            n7740;
wire            n7741;
wire      [7:0] n7742;
wire            n7743;
wire            n7744;
wire            n7745;
wire            n7746;
wire            n7747;
wire      [7:0] n7748;
wire            n7749;
wire      [7:0] n775;
wire            n7750;
wire            n7751;
wire            n7752;
wire            n7753;
wire      [7:0] n7754;
wire            n7755;
wire            n7756;
wire            n7757;
wire            n7758;
wire            n7759;
wire      [7:0] n776;
wire      [7:0] n7760;
wire            n7761;
wire            n7762;
wire            n7763;
wire            n7764;
wire            n7765;
wire      [7:0] n7766;
wire            n7767;
wire            n7768;
wire            n7769;
wire      [7:0] n777;
wire            n7770;
wire            n7771;
wire      [7:0] n7772;
wire            n7773;
wire            n7774;
wire            n7775;
wire            n7776;
wire            n7777;
wire      [7:0] n7778;
wire            n7779;
wire      [7:0] n778;
wire            n7780;
wire            n7781;
wire            n7782;
wire            n7783;
wire      [7:0] n7784;
wire            n7785;
wire            n7786;
wire            n7787;
wire            n7788;
wire            n7789;
wire      [7:0] n779;
wire      [7:0] n7790;
wire            n7791;
wire            n7792;
wire            n7793;
wire            n7794;
wire            n7795;
wire      [7:0] n7796;
wire            n7797;
wire            n7798;
wire            n7799;
wire            n78;
wire      [7:0] n780;
wire            n7800;
wire            n7801;
wire      [7:0] n7802;
wire            n7803;
wire            n7804;
wire            n7805;
wire            n7806;
wire            n7807;
wire      [7:0] n7808;
wire            n7809;
wire      [7:0] n781;
wire            n7810;
wire            n7811;
wire            n7812;
wire            n7813;
wire      [7:0] n7814;
wire            n7815;
wire            n7816;
wire            n7817;
wire            n7818;
wire            n7819;
wire      [7:0] n782;
wire      [7:0] n7820;
wire            n7821;
wire            n7822;
wire            n7823;
wire            n7824;
wire            n7825;
wire      [7:0] n7826;
wire            n7827;
wire            n7828;
wire            n7829;
wire      [7:0] n783;
wire            n7830;
wire            n7831;
wire      [7:0] n7832;
wire            n7833;
wire            n7834;
wire            n7835;
wire            n7836;
wire            n7837;
wire      [7:0] n7838;
wire            n7839;
wire      [7:0] n784;
wire            n7840;
wire            n7841;
wire            n7842;
wire            n7843;
wire      [7:0] n7844;
wire            n7845;
wire            n7846;
wire            n7847;
wire            n7848;
wire            n7849;
wire      [7:0] n785;
wire      [7:0] n7850;
wire            n7851;
wire            n7852;
wire            n7853;
wire            n7854;
wire            n7855;
wire      [7:0] n7856;
wire            n7857;
wire            n7858;
wire            n7859;
wire      [7:0] n786;
wire            n7860;
wire            n7861;
wire      [7:0] n7862;
wire            n7863;
wire            n7864;
wire            n7865;
wire            n7866;
wire            n7867;
wire      [7:0] n7868;
wire            n7869;
wire      [7:0] n787;
wire            n7870;
wire            n7871;
wire            n7872;
wire            n7873;
wire      [7:0] n7874;
wire            n7875;
wire            n7876;
wire            n7877;
wire            n7878;
wire            n7879;
wire      [7:0] n788;
wire      [7:0] n7880;
wire            n7881;
wire            n7882;
wire            n7883;
wire            n7884;
wire            n7885;
wire      [7:0] n7886;
wire            n7887;
wire            n7888;
wire            n7889;
wire      [7:0] n789;
wire            n7890;
wire            n7891;
wire      [7:0] n7892;
wire            n7893;
wire            n7894;
wire            n7895;
wire            n7896;
wire            n7897;
wire      [7:0] n7898;
wire            n7899;
wire      [7:0] n790;
wire            n7900;
wire            n7901;
wire            n7902;
wire            n7903;
wire      [7:0] n7904;
wire            n7905;
wire            n7906;
wire            n7907;
wire            n7908;
wire            n7909;
wire      [7:0] n791;
wire      [7:0] n7910;
wire            n7911;
wire            n7912;
wire            n7913;
wire            n7914;
wire            n7915;
wire      [7:0] n7916;
wire            n7917;
wire            n7918;
wire            n7919;
wire      [7:0] n792;
wire            n7920;
wire            n7921;
wire      [7:0] n7922;
wire            n7923;
wire            n7924;
wire            n7925;
wire            n7926;
wire            n7927;
wire      [7:0] n7928;
wire            n7929;
wire      [7:0] n793;
wire            n7930;
wire            n7931;
wire            n7932;
wire            n7933;
wire      [7:0] n7934;
wire            n7935;
wire            n7936;
wire            n7937;
wire            n7938;
wire            n7939;
wire      [7:0] n794;
wire      [7:0] n7940;
wire            n7941;
wire            n7942;
wire            n7943;
wire            n7944;
wire            n7945;
wire      [7:0] n7946;
wire            n7947;
wire            n7948;
wire            n7949;
wire      [7:0] n795;
wire            n7950;
wire            n7951;
wire      [7:0] n7952;
wire            n7953;
wire            n7954;
wire            n7955;
wire            n7956;
wire            n7957;
wire      [7:0] n7958;
wire            n7959;
wire      [7:0] n796;
wire            n7960;
wire            n7961;
wire            n7962;
wire            n7963;
wire      [7:0] n7964;
wire            n7965;
wire            n7966;
wire            n7967;
wire            n7968;
wire            n7969;
wire      [7:0] n797;
wire      [7:0] n7970;
wire            n7971;
wire            n7972;
wire            n7973;
wire            n7974;
wire            n7975;
wire      [7:0] n7976;
wire            n7977;
wire            n7978;
wire            n7979;
wire      [7:0] n798;
wire            n7980;
wire            n7981;
wire      [7:0] n7982;
wire            n7983;
wire            n7984;
wire            n7985;
wire            n7986;
wire            n7987;
wire      [7:0] n7988;
wire            n7989;
wire      [7:0] n799;
wire            n7990;
wire            n7991;
wire            n7992;
wire            n7993;
wire      [7:0] n7994;
wire            n7995;
wire            n7996;
wire            n7997;
wire            n7998;
wire            n7999;
wire            n80;
wire      [7:0] n800;
wire      [7:0] n8000;
wire            n8001;
wire            n8002;
wire            n8003;
wire            n8004;
wire            n8005;
wire      [7:0] n8006;
wire            n8007;
wire            n8008;
wire            n8009;
wire      [7:0] n801;
wire            n8010;
wire            n8011;
wire      [7:0] n8012;
wire            n8013;
wire            n8014;
wire            n8015;
wire            n8016;
wire            n8017;
wire      [7:0] n8018;
wire            n8019;
wire      [7:0] n802;
wire            n8020;
wire            n8021;
wire            n8022;
wire            n8023;
wire      [7:0] n8024;
wire            n8025;
wire            n8026;
wire            n8027;
wire            n8028;
wire            n8029;
wire      [7:0] n803;
wire      [7:0] n8030;
wire            n8031;
wire            n8032;
wire            n8033;
wire            n8034;
wire            n8035;
wire      [7:0] n8036;
wire            n8037;
wire            n8038;
wire            n8039;
wire      [7:0] n804;
wire            n8040;
wire            n8041;
wire      [7:0] n8042;
wire            n8043;
wire            n8044;
wire            n8045;
wire            n8046;
wire            n8047;
wire      [7:0] n8048;
wire            n8049;
wire      [7:0] n805;
wire            n8050;
wire            n8051;
wire            n8052;
wire            n8053;
wire      [7:0] n8054;
wire            n8055;
wire            n8056;
wire            n8057;
wire            n8058;
wire            n8059;
wire      [7:0] n806;
wire      [7:0] n8060;
wire            n8061;
wire            n8062;
wire            n8063;
wire            n8064;
wire            n8065;
wire      [7:0] n8066;
wire            n8067;
wire            n8068;
wire            n8069;
wire      [7:0] n807;
wire            n8070;
wire            n8071;
wire      [7:0] n8072;
wire            n8073;
wire            n8074;
wire            n8075;
wire            n8076;
wire            n8077;
wire      [7:0] n8078;
wire            n8079;
wire      [7:0] n808;
wire            n8080;
wire            n8081;
wire            n8082;
wire            n8083;
wire      [7:0] n8084;
wire            n8085;
wire            n8086;
wire            n8087;
wire            n8088;
wire            n8089;
wire      [7:0] n809;
wire      [7:0] n8090;
wire            n8091;
wire            n8092;
wire            n8093;
wire            n8094;
wire            n8095;
wire      [7:0] n8096;
wire            n8097;
wire            n8098;
wire            n8099;
wire      [7:0] n810;
wire            n8100;
wire            n8101;
wire      [7:0] n8102;
wire            n8103;
wire            n8104;
wire            n8105;
wire            n8106;
wire            n8107;
wire      [7:0] n8108;
wire            n8109;
wire      [7:0] n811;
wire            n8110;
wire            n8111;
wire            n8112;
wire            n8113;
wire      [7:0] n8114;
wire            n8115;
wire            n8116;
wire            n8117;
wire            n8118;
wire            n8119;
wire      [7:0] n812;
wire      [7:0] n8120;
wire            n8121;
wire            n8122;
wire            n8123;
wire            n8124;
wire            n8125;
wire      [7:0] n8126;
wire            n8127;
wire            n8128;
wire            n8129;
wire      [7:0] n813;
wire            n8130;
wire            n8131;
wire      [7:0] n8132;
wire            n8133;
wire            n8134;
wire            n8135;
wire            n8136;
wire            n8137;
wire      [7:0] n8138;
wire            n8139;
wire      [7:0] n814;
wire            n8140;
wire            n8141;
wire            n8142;
wire            n8143;
wire      [7:0] n8144;
wire            n8145;
wire            n8146;
wire            n8147;
wire            n8148;
wire            n8149;
wire      [7:0] n815;
wire      [7:0] n8150;
wire            n8151;
wire            n8152;
wire            n8153;
wire            n8154;
wire            n8155;
wire      [7:0] n8156;
wire            n8157;
wire            n8158;
wire            n8159;
wire      [7:0] n816;
wire            n8160;
wire            n8161;
wire      [7:0] n8162;
wire            n8163;
wire            n8164;
wire            n8165;
wire            n8166;
wire            n8167;
wire      [7:0] n8168;
wire            n8169;
wire      [7:0] n817;
wire            n8170;
wire            n8171;
wire            n8172;
wire            n8173;
wire      [7:0] n8174;
wire            n8175;
wire            n8176;
wire            n8177;
wire            n8178;
wire            n8179;
wire      [7:0] n818;
wire      [7:0] n8180;
wire            n8181;
wire            n8182;
wire            n8183;
wire            n8184;
wire            n8185;
wire      [7:0] n8186;
wire            n8187;
wire            n8188;
wire            n8189;
wire      [7:0] n819;
wire            n8190;
wire            n8191;
wire      [7:0] n8192;
wire            n8193;
wire            n8194;
wire            n8195;
wire            n8196;
wire            n8197;
wire      [7:0] n8198;
wire            n8199;
wire            n82;
wire      [7:0] n820;
wire            n8200;
wire            n8201;
wire            n8202;
wire            n8203;
wire      [7:0] n8204;
wire            n8205;
wire            n8206;
wire            n8207;
wire            n8208;
wire            n8209;
wire      [7:0] n821;
wire      [7:0] n8210;
wire            n8211;
wire            n8212;
wire            n8213;
wire            n8214;
wire            n8215;
wire      [7:0] n8216;
wire            n8217;
wire            n8218;
wire            n8219;
wire      [7:0] n822;
wire            n8220;
wire            n8221;
wire      [7:0] n8222;
wire            n8223;
wire            n8224;
wire            n8225;
wire            n8226;
wire            n8227;
wire      [7:0] n8228;
wire            n8229;
wire      [7:0] n823;
wire            n8230;
wire            n8231;
wire            n8232;
wire            n8233;
wire      [7:0] n8234;
wire            n8235;
wire            n8236;
wire            n8237;
wire            n8238;
wire            n8239;
wire      [7:0] n824;
wire      [7:0] n8240;
wire            n8241;
wire            n8242;
wire            n8243;
wire            n8244;
wire            n8245;
wire      [7:0] n8246;
wire            n8247;
wire            n8248;
wire            n8249;
wire      [7:0] n825;
wire            n8250;
wire            n8251;
wire      [7:0] n8252;
wire            n8253;
wire            n8254;
wire            n8255;
wire            n8256;
wire            n8257;
wire      [7:0] n8258;
wire            n8259;
wire      [7:0] n826;
wire            n8260;
wire            n8261;
wire            n8262;
wire            n8263;
wire      [7:0] n8264;
wire            n8265;
wire            n8266;
wire            n8267;
wire            n8268;
wire            n8269;
wire      [7:0] n827;
wire      [7:0] n8270;
wire            n8271;
wire            n8272;
wire            n8273;
wire            n8274;
wire            n8275;
wire      [7:0] n8276;
wire            n8277;
wire            n8278;
wire            n8279;
wire      [7:0] n828;
wire            n8280;
wire            n8281;
wire      [7:0] n8282;
wire            n8283;
wire            n8284;
wire            n8285;
wire            n8286;
wire            n8287;
wire      [7:0] n8288;
wire            n8289;
wire      [7:0] n829;
wire            n8290;
wire            n8291;
wire            n8292;
wire            n8293;
wire      [7:0] n8294;
wire            n8295;
wire            n8296;
wire            n8297;
wire            n8298;
wire            n8299;
wire      [7:0] n830;
wire      [7:0] n8300;
wire            n8301;
wire            n8302;
wire            n8303;
wire            n8304;
wire            n8305;
wire      [7:0] n8306;
wire            n8307;
wire            n8308;
wire            n8309;
wire      [7:0] n831;
wire            n8310;
wire            n8311;
wire      [7:0] n8312;
wire            n8313;
wire            n8314;
wire            n8315;
wire            n8316;
wire            n8317;
wire      [7:0] n8318;
wire            n8319;
wire      [7:0] n832;
wire            n8320;
wire            n8321;
wire            n8322;
wire            n8323;
wire      [7:0] n8324;
wire            n8325;
wire            n8326;
wire            n8327;
wire            n8328;
wire            n8329;
wire      [7:0] n833;
wire      [7:0] n8330;
wire            n8331;
wire            n8332;
wire            n8333;
wire            n8334;
wire            n8335;
wire      [7:0] n8336;
wire            n8337;
wire            n8338;
wire            n8339;
wire            n834;
wire            n8340;
wire            n8341;
wire      [7:0] n8342;
wire            n8343;
wire            n8344;
wire            n8345;
wire            n8346;
wire            n8347;
wire      [7:0] n8348;
wire            n8349;
wire            n835;
wire            n8350;
wire            n8351;
wire            n8352;
wire            n8353;
wire      [7:0] n8354;
wire            n8355;
wire            n8356;
wire            n8357;
wire            n8358;
wire            n8359;
wire            n836;
wire      [7:0] n8360;
wire            n8361;
wire            n8362;
wire            n8363;
wire            n8364;
wire            n8365;
wire      [7:0] n8366;
wire            n8367;
wire            n8368;
wire            n8369;
wire            n837;
wire            n8370;
wire            n8371;
wire      [7:0] n8372;
wire            n8373;
wire            n8374;
wire            n8375;
wire            n8376;
wire            n8377;
wire      [7:0] n8378;
wire            n8379;
wire            n838;
wire            n8380;
wire            n8381;
wire            n8382;
wire            n8383;
wire      [7:0] n8384;
wire            n8385;
wire            n8386;
wire            n8387;
wire            n8388;
wire            n8389;
wire            n839;
wire      [7:0] n8390;
wire            n8391;
wire            n8392;
wire            n8393;
wire            n8394;
wire            n8395;
wire      [7:0] n8396;
wire            n8397;
wire            n8398;
wire            n8399;
wire            n84;
wire            n840;
wire            n8400;
wire            n8401;
wire      [7:0] n8402;
wire            n8403;
wire            n8404;
wire            n8405;
wire            n8406;
wire            n8407;
wire      [7:0] n8408;
wire            n8409;
wire            n841;
wire            n8410;
wire            n8411;
wire            n8412;
wire            n8413;
wire      [7:0] n8414;
wire            n8415;
wire            n8416;
wire            n8417;
wire            n8418;
wire            n8419;
wire            n842;
wire      [7:0] n8420;
wire            n8421;
wire            n8422;
wire            n8423;
wire            n8424;
wire            n8425;
wire      [7:0] n8426;
wire            n8427;
wire            n8428;
wire            n8429;
wire            n843;
wire            n8430;
wire            n8431;
wire      [7:0] n8432;
wire            n8433;
wire            n8434;
wire            n8435;
wire            n8436;
wire            n8437;
wire      [7:0] n8438;
wire            n8439;
wire            n844;
wire            n8440;
wire            n8441;
wire            n8442;
wire            n8443;
wire      [7:0] n8444;
wire            n8445;
wire            n8446;
wire            n8447;
wire            n8448;
wire            n8449;
wire            n845;
wire      [7:0] n8450;
wire            n8451;
wire            n8452;
wire            n8453;
wire            n8454;
wire            n8455;
wire      [7:0] n8456;
wire            n8457;
wire            n8458;
wire            n8459;
wire            n846;
wire            n8460;
wire            n8461;
wire      [7:0] n8462;
wire            n8463;
wire            n8464;
wire            n8465;
wire            n8466;
wire            n8467;
wire      [7:0] n8468;
wire            n8469;
wire            n847;
wire            n8470;
wire            n8471;
wire            n8472;
wire            n8473;
wire      [7:0] n8474;
wire            n8475;
wire            n8476;
wire            n8477;
wire            n8478;
wire            n8479;
wire            n848;
wire      [7:0] n8480;
wire            n8481;
wire            n8482;
wire            n8483;
wire            n8484;
wire            n8485;
wire      [7:0] n8486;
wire            n8487;
wire            n8488;
wire            n8489;
wire            n849;
wire            n8490;
wire            n8491;
wire      [7:0] n8492;
wire            n8493;
wire            n8494;
wire            n8495;
wire            n8496;
wire            n8497;
wire      [7:0] n8498;
wire            n8499;
wire            n850;
wire            n8500;
wire            n8501;
wire            n8502;
wire            n8503;
wire      [7:0] n8504;
wire            n8505;
wire            n8506;
wire            n8507;
wire            n8508;
wire            n8509;
wire            n851;
wire      [7:0] n8510;
wire            n8511;
wire            n8512;
wire            n8513;
wire            n8514;
wire            n8515;
wire      [7:0] n8516;
wire            n8517;
wire            n8518;
wire            n8519;
wire            n852;
wire            n8520;
wire            n8521;
wire      [7:0] n8522;
wire            n8523;
wire            n8524;
wire            n8525;
wire            n8526;
wire            n8527;
wire      [7:0] n8528;
wire            n8529;
wire            n853;
wire            n8530;
wire            n8531;
wire            n8532;
wire            n8533;
wire      [7:0] n8534;
wire            n8535;
wire            n8536;
wire            n8537;
wire            n8538;
wire            n8539;
wire            n854;
wire      [7:0] n8540;
wire            n8541;
wire            n8542;
wire            n8543;
wire            n8544;
wire            n8545;
wire      [7:0] n8546;
wire            n8547;
wire            n8548;
wire            n8549;
wire            n855;
wire            n8550;
wire            n8551;
wire      [7:0] n8552;
wire            n8553;
wire            n8554;
wire            n8555;
wire            n8556;
wire            n8557;
wire      [7:0] n8558;
wire            n8559;
wire            n856;
wire            n8560;
wire            n8561;
wire            n8562;
wire            n8563;
wire      [7:0] n8564;
wire            n8565;
wire            n8566;
wire            n8567;
wire            n8568;
wire            n8569;
wire            n857;
wire      [7:0] n8570;
wire            n8571;
wire            n8572;
wire            n8573;
wire            n8574;
wire            n8575;
wire      [7:0] n8576;
wire            n8577;
wire            n8578;
wire            n8579;
wire            n858;
wire            n8580;
wire            n8581;
wire      [7:0] n8582;
wire            n8583;
wire            n8584;
wire            n8585;
wire            n8586;
wire            n8587;
wire      [7:0] n8588;
wire            n8589;
wire            n859;
wire            n8590;
wire            n8591;
wire            n8592;
wire            n8593;
wire      [7:0] n8594;
wire            n8595;
wire            n8596;
wire            n8597;
wire            n8598;
wire            n8599;
wire            n86;
wire            n860;
wire      [7:0] n8600;
wire            n8601;
wire            n8602;
wire            n8603;
wire            n8604;
wire            n8605;
wire      [7:0] n8606;
wire            n8607;
wire            n8608;
wire            n8609;
wire            n861;
wire            n8610;
wire            n8611;
wire      [7:0] n8612;
wire            n8613;
wire            n8614;
wire            n8615;
wire            n8616;
wire            n8617;
wire      [7:0] n8618;
wire            n8619;
wire            n862;
wire            n8620;
wire            n8621;
wire            n8622;
wire            n8623;
wire      [7:0] n8624;
wire            n8625;
wire            n8626;
wire            n8627;
wire            n8628;
wire            n8629;
wire            n863;
wire      [7:0] n8630;
wire            n8631;
wire            n8632;
wire            n8633;
wire            n8634;
wire            n8635;
wire      [7:0] n8636;
wire            n8637;
wire            n8638;
wire            n8639;
wire            n864;
wire            n8640;
wire            n8641;
wire      [7:0] n8642;
wire            n8643;
wire            n8644;
wire            n8645;
wire            n8646;
wire            n8647;
wire      [7:0] n8648;
wire            n8649;
wire            n865;
wire            n8650;
wire            n8651;
wire            n8652;
wire            n8653;
wire      [7:0] n8654;
wire            n8655;
wire            n8656;
wire            n8657;
wire            n8658;
wire            n8659;
wire            n866;
wire      [7:0] n8660;
wire            n8661;
wire            n8662;
wire            n8663;
wire            n8664;
wire            n8665;
wire      [7:0] n8666;
wire            n8667;
wire            n8668;
wire            n8669;
wire            n867;
wire            n8670;
wire            n8671;
wire      [7:0] n8672;
wire            n8673;
wire            n8674;
wire            n8675;
wire            n8676;
wire            n8677;
wire      [7:0] n8678;
wire            n8679;
wire            n868;
wire            n8680;
wire            n8681;
wire            n8682;
wire            n8683;
wire      [7:0] n8684;
wire            n8685;
wire            n8686;
wire            n8687;
wire            n8688;
wire            n8689;
wire            n869;
wire      [7:0] n8690;
wire            n8691;
wire            n8692;
wire            n8693;
wire            n8694;
wire            n8695;
wire      [7:0] n8696;
wire            n8697;
wire            n8698;
wire            n8699;
wire            n870;
wire            n8700;
wire            n8701;
wire      [7:0] n8702;
wire            n8703;
wire            n8704;
wire            n8705;
wire            n8706;
wire            n8707;
wire      [7:0] n8708;
wire            n8709;
wire            n871;
wire            n8710;
wire            n8711;
wire            n8712;
wire            n8713;
wire      [7:0] n8714;
wire            n8715;
wire            n8716;
wire            n8717;
wire            n8718;
wire            n8719;
wire            n872;
wire      [7:0] n8720;
wire            n8721;
wire            n8722;
wire            n8723;
wire            n8724;
wire            n8725;
wire      [7:0] n8726;
wire            n8727;
wire            n8728;
wire            n8729;
wire            n873;
wire            n8730;
wire            n8731;
wire      [7:0] n8732;
wire            n8733;
wire            n8734;
wire            n8735;
wire            n8736;
wire            n8737;
wire      [7:0] n8738;
wire            n8739;
wire            n874;
wire            n8740;
wire            n8741;
wire            n8742;
wire            n8743;
wire      [7:0] n8744;
wire            n8745;
wire            n8746;
wire            n8747;
wire            n8748;
wire            n8749;
wire            n875;
wire      [7:0] n8750;
wire            n8751;
wire            n8752;
wire            n8753;
wire            n8754;
wire            n8755;
wire      [7:0] n8756;
wire            n8757;
wire            n8758;
wire            n8759;
wire            n876;
wire            n8760;
wire            n8761;
wire      [7:0] n8762;
wire            n8763;
wire            n8764;
wire            n8765;
wire            n8766;
wire            n8767;
wire      [7:0] n8768;
wire            n8769;
wire            n877;
wire            n8770;
wire            n8771;
wire            n8772;
wire            n8773;
wire      [7:0] n8774;
wire            n8775;
wire            n8776;
wire            n8777;
wire            n8778;
wire            n8779;
wire            n878;
wire      [7:0] n8780;
wire            n8781;
wire            n8782;
wire            n8783;
wire            n8784;
wire            n8785;
wire      [7:0] n8786;
wire            n8787;
wire            n8788;
wire            n8789;
wire            n879;
wire            n8790;
wire            n8791;
wire      [7:0] n8792;
wire            n8793;
wire            n8794;
wire            n8795;
wire            n8796;
wire            n8797;
wire      [7:0] n8798;
wire            n8799;
wire            n88;
wire            n880;
wire            n8800;
wire            n8801;
wire            n8802;
wire            n8803;
wire      [7:0] n8804;
wire            n8805;
wire            n8806;
wire            n8807;
wire            n8808;
wire            n8809;
wire            n881;
wire      [7:0] n8810;
wire            n8811;
wire            n8812;
wire            n8813;
wire            n8814;
wire            n8815;
wire      [7:0] n8816;
wire            n8817;
wire            n8818;
wire            n8819;
wire            n882;
wire            n8820;
wire            n8821;
wire      [7:0] n8822;
wire            n8823;
wire            n8824;
wire            n8825;
wire            n8826;
wire            n8827;
wire      [7:0] n8828;
wire            n8829;
wire            n883;
wire            n8830;
wire            n8831;
wire            n8832;
wire            n8833;
wire      [7:0] n8834;
wire            n8835;
wire            n8836;
wire            n8837;
wire            n8838;
wire            n8839;
wire            n884;
wire      [7:0] n8840;
wire            n8841;
wire            n8842;
wire            n8843;
wire            n8844;
wire            n8845;
wire      [7:0] n8846;
wire            n8847;
wire            n8848;
wire            n8849;
wire            n885;
wire            n8850;
wire            n8851;
wire      [7:0] n8852;
wire            n8853;
wire            n8854;
wire            n8855;
wire            n8856;
wire            n8857;
wire      [7:0] n8858;
wire            n8859;
wire            n886;
wire            n8860;
wire            n8861;
wire            n8862;
wire            n8863;
wire      [7:0] n8864;
wire            n8865;
wire            n8866;
wire            n8867;
wire            n8868;
wire            n8869;
wire            n887;
wire      [7:0] n8870;
wire            n8871;
wire            n8872;
wire            n8873;
wire            n8874;
wire            n8875;
wire      [7:0] n8876;
wire            n8877;
wire            n8878;
wire            n8879;
wire            n888;
wire            n8880;
wire            n8881;
wire      [7:0] n8882;
wire            n8883;
wire            n8884;
wire            n8885;
wire            n8886;
wire            n8887;
wire      [7:0] n8888;
wire            n8889;
wire            n889;
wire            n8890;
wire            n8891;
wire            n8892;
wire            n8893;
wire      [7:0] n8894;
wire            n8895;
wire            n8896;
wire            n8897;
wire            n8898;
wire            n8899;
wire            n890;
wire      [7:0] n8900;
wire            n8901;
wire            n8902;
wire            n8903;
wire            n8904;
wire            n8905;
wire      [7:0] n8906;
wire            n8907;
wire            n8908;
wire            n8909;
wire            n891;
wire            n8910;
wire            n8911;
wire      [7:0] n8912;
wire            n8913;
wire            n8914;
wire            n8915;
wire            n8916;
wire            n8917;
wire      [7:0] n8918;
wire            n8919;
wire            n892;
wire            n8920;
wire            n8921;
wire            n8922;
wire            n8923;
wire      [7:0] n8924;
wire            n8925;
wire            n8926;
wire            n8927;
wire            n8928;
wire            n8929;
wire            n893;
wire      [7:0] n8930;
wire            n8931;
wire            n8932;
wire            n8933;
wire            n8934;
wire            n8935;
wire      [7:0] n8936;
wire            n8937;
wire            n8938;
wire            n8939;
wire            n894;
wire            n8940;
wire            n8941;
wire      [7:0] n8942;
wire            n8943;
wire            n8944;
wire            n8945;
wire            n8946;
wire            n8947;
wire      [7:0] n8948;
wire            n8949;
wire            n895;
wire            n8950;
wire            n8951;
wire            n8952;
wire            n8953;
wire      [7:0] n8954;
wire            n8955;
wire            n8956;
wire            n8957;
wire            n8958;
wire            n8959;
wire            n896;
wire      [7:0] n8960;
wire            n8961;
wire            n8962;
wire            n8963;
wire            n8964;
wire            n8965;
wire      [7:0] n8966;
wire            n8967;
wire            n8968;
wire            n8969;
wire            n897;
wire            n8970;
wire            n8971;
wire      [7:0] n8972;
wire            n8973;
wire            n8974;
wire            n8975;
wire            n8976;
wire            n8977;
wire      [7:0] n8978;
wire            n8979;
wire            n898;
wire            n8980;
wire            n8981;
wire            n8982;
wire            n8983;
wire      [7:0] n8984;
wire            n8985;
wire            n8986;
wire            n8987;
wire            n8988;
wire            n8989;
wire            n899;
wire      [7:0] n8990;
wire            n8991;
wire            n8992;
wire            n8993;
wire            n8994;
wire            n8995;
wire      [7:0] n8996;
wire            n8997;
wire            n8998;
wire            n8999;
wire            n9;
wire            n90;
wire            n900;
wire            n9000;
wire            n9001;
wire      [7:0] n9002;
wire            n9003;
wire            n9004;
wire            n9005;
wire            n9006;
wire            n9007;
wire      [7:0] n9008;
wire            n9009;
wire            n901;
wire            n9010;
wire            n9011;
wire            n9012;
wire            n9013;
wire      [7:0] n9014;
wire            n9015;
wire            n9016;
wire            n9017;
wire            n9018;
wire            n9019;
wire            n902;
wire      [7:0] n9020;
wire            n9021;
wire            n9022;
wire            n9023;
wire            n9024;
wire            n9025;
wire      [7:0] n9026;
wire            n9027;
wire            n9028;
wire            n9029;
wire            n903;
wire            n9030;
wire            n9031;
wire      [7:0] n9032;
wire            n9033;
wire            n9034;
wire            n9035;
wire            n9036;
wire            n9037;
wire      [7:0] n9038;
wire            n9039;
wire            n904;
wire            n9040;
wire            n9041;
wire            n9042;
wire            n9043;
wire      [7:0] n9044;
wire            n9045;
wire            n9046;
wire            n9047;
wire            n9048;
wire            n9049;
wire            n905;
wire      [7:0] n9050;
wire            n9051;
wire            n9052;
wire            n9053;
wire            n9054;
wire            n9055;
wire      [7:0] n9056;
wire            n9057;
wire            n9058;
wire            n9059;
wire            n906;
wire            n9060;
wire            n9061;
wire      [7:0] n9062;
wire            n9063;
wire            n9064;
wire            n9065;
wire            n9066;
wire            n9067;
wire      [7:0] n9068;
wire            n9069;
wire            n907;
wire            n9070;
wire            n9071;
wire            n9072;
wire            n9073;
wire      [7:0] n9074;
wire            n9075;
wire            n9076;
wire            n9077;
wire            n9078;
wire            n9079;
wire            n908;
wire      [7:0] n9080;
wire            n9081;
wire            n9082;
wire            n9083;
wire            n9084;
wire            n9085;
wire      [7:0] n9086;
wire            n9087;
wire            n9088;
wire            n9089;
wire            n909;
wire            n9090;
wire            n9091;
wire      [7:0] n9092;
wire            n9093;
wire            n9094;
wire            n9095;
wire            n9096;
wire            n9097;
wire      [7:0] n9098;
wire            n9099;
wire            n910;
wire            n9100;
wire            n9101;
wire            n9102;
wire            n9103;
wire      [7:0] n9104;
wire            n9105;
wire            n9106;
wire            n9107;
wire            n9108;
wire            n9109;
wire            n911;
wire      [7:0] n9110;
wire            n9111;
wire            n9112;
wire            n9113;
wire            n9114;
wire            n9115;
wire      [7:0] n9116;
wire            n9117;
wire            n9118;
wire            n9119;
wire            n912;
wire            n9120;
wire            n9121;
wire      [7:0] n9122;
wire            n9123;
wire            n9124;
wire            n9125;
wire            n9126;
wire            n9127;
wire      [7:0] n9128;
wire            n9129;
wire            n913;
wire            n9130;
wire            n9131;
wire            n9132;
wire            n9133;
wire      [7:0] n9134;
wire            n9135;
wire            n9136;
wire            n9137;
wire            n9138;
wire            n9139;
wire            n914;
wire      [7:0] n9140;
wire            n9141;
wire            n9142;
wire            n9143;
wire            n9144;
wire            n9145;
wire      [7:0] n9146;
wire            n9147;
wire            n9148;
wire            n9149;
wire            n915;
wire            n9150;
wire            n9151;
wire      [7:0] n9152;
wire            n9153;
wire            n9154;
wire            n9155;
wire            n9156;
wire            n9157;
wire      [7:0] n9158;
wire            n9159;
wire            n916;
wire            n9160;
wire            n9161;
wire            n9162;
wire            n9163;
wire      [7:0] n9164;
wire            n9165;
wire            n9166;
wire            n9167;
wire            n9168;
wire            n9169;
wire            n917;
wire      [7:0] n9170;
wire            n9171;
wire            n9172;
wire            n9173;
wire            n9174;
wire            n9175;
wire      [7:0] n9176;
wire            n9177;
wire            n9178;
wire            n9179;
wire            n918;
wire            n9180;
wire            n9181;
wire      [7:0] n9182;
wire            n9183;
wire            n9184;
wire            n9185;
wire            n9186;
wire            n9187;
wire      [7:0] n9188;
wire            n9189;
wire            n919;
wire            n9190;
wire            n9191;
wire            n9192;
wire            n9193;
wire      [7:0] n9194;
wire            n9195;
wire            n9196;
wire            n9197;
wire            n9198;
wire            n9199;
wire            n92;
wire            n920;
wire      [7:0] n9200;
wire            n9201;
wire            n9202;
wire            n9203;
wire            n9204;
wire            n9205;
wire      [7:0] n9206;
wire            n9207;
wire            n9208;
wire            n9209;
wire            n921;
wire            n9210;
wire            n9211;
wire      [7:0] n9212;
wire            n9213;
wire            n9214;
wire            n9215;
wire            n9216;
wire            n9217;
wire      [7:0] n9218;
wire            n9219;
wire            n922;
wire            n9220;
wire            n9221;
wire            n9222;
wire            n9223;
wire      [7:0] n9224;
wire            n9225;
wire            n9226;
wire            n9227;
wire            n9228;
wire            n9229;
wire            n923;
wire      [7:0] n9230;
wire            n9231;
wire            n9232;
wire            n9233;
wire            n9234;
wire            n9235;
wire      [7:0] n9236;
wire            n9237;
wire            n9238;
wire            n9239;
wire            n924;
wire            n9240;
wire            n9241;
wire      [7:0] n9242;
wire            n9243;
wire            n9244;
wire            n9245;
wire            n9246;
wire            n9247;
wire      [7:0] n9248;
wire            n9249;
wire            n925;
wire            n9250;
wire            n9251;
wire            n9252;
wire            n9253;
wire      [7:0] n9254;
wire            n9255;
wire            n9256;
wire            n9257;
wire            n9258;
wire            n9259;
wire            n926;
wire      [7:0] n9260;
wire            n9261;
wire            n9262;
wire            n9263;
wire            n9264;
wire            n9265;
wire      [7:0] n9266;
wire            n9267;
wire            n9268;
wire            n9269;
wire            n927;
wire            n9270;
wire            n9271;
wire      [7:0] n9272;
wire            n9273;
wire            n9274;
wire            n9275;
wire            n9276;
wire            n9277;
wire      [7:0] n9278;
wire            n9279;
wire            n928;
wire            n9280;
wire            n9281;
wire            n9282;
wire            n9283;
wire      [7:0] n9284;
wire            n9285;
wire            n9286;
wire            n9287;
wire            n9288;
wire            n9289;
wire            n929;
wire      [7:0] n9290;
wire            n9291;
wire            n9292;
wire            n9293;
wire            n9294;
wire            n9295;
wire      [7:0] n9296;
wire            n9297;
wire            n9298;
wire            n9299;
wire            n930;
wire            n9300;
wire            n9301;
wire      [7:0] n9302;
wire            n9303;
wire            n9304;
wire            n9305;
wire            n9306;
wire            n9307;
wire      [7:0] n9308;
wire            n9309;
wire            n931;
wire            n9310;
wire            n9311;
wire            n9312;
wire            n9313;
wire      [7:0] n9314;
wire            n9315;
wire            n9316;
wire            n9317;
wire            n9318;
wire            n9319;
wire            n932;
wire      [7:0] n9320;
wire            n9321;
wire            n9322;
wire            n9323;
wire            n9324;
wire            n9325;
wire      [7:0] n9326;
wire            n9327;
wire            n9328;
wire            n9329;
wire            n933;
wire            n9330;
wire            n9331;
wire      [7:0] n9332;
wire            n9333;
wire            n9334;
wire            n9335;
wire            n9336;
wire            n9337;
wire      [7:0] n9338;
wire            n9339;
wire            n934;
wire            n9340;
wire            n9341;
wire            n9342;
wire            n9343;
wire      [7:0] n9344;
wire            n9345;
wire            n9346;
wire            n9347;
wire            n9348;
wire            n9349;
wire            n935;
wire      [7:0] n9350;
wire            n9351;
wire            n9352;
wire            n9353;
wire            n9354;
wire            n9355;
wire      [7:0] n9356;
wire            n9357;
wire            n9358;
wire            n9359;
wire            n936;
wire            n9360;
wire            n9361;
wire      [7:0] n9362;
wire            n9363;
wire            n9364;
wire            n9365;
wire            n9366;
wire            n9367;
wire      [7:0] n9368;
wire            n9369;
wire            n937;
wire            n9370;
wire            n9371;
wire            n9372;
wire            n9373;
wire      [7:0] n9374;
wire            n9375;
wire            n9376;
wire            n9377;
wire            n9378;
wire            n9379;
wire            n938;
wire      [7:0] n9380;
wire            n9381;
wire            n9382;
wire            n9383;
wire            n9384;
wire            n9385;
wire      [7:0] n9386;
wire            n9387;
wire            n9388;
wire            n9389;
wire            n939;
wire            n9390;
wire            n9391;
wire      [7:0] n9392;
wire            n9393;
wire            n9394;
wire            n9395;
wire            n9396;
wire            n9397;
wire      [7:0] n9398;
wire            n9399;
wire            n94;
wire            n940;
wire            n9400;
wire            n9401;
wire            n9402;
wire            n9403;
wire      [7:0] n9404;
wire            n9405;
wire            n9406;
wire            n9407;
wire            n9408;
wire            n9409;
wire            n941;
wire      [7:0] n9410;
wire            n9411;
wire            n9412;
wire            n9413;
wire            n9414;
wire            n9415;
wire      [7:0] n9416;
wire            n9417;
wire            n9418;
wire            n9419;
wire            n942;
wire            n9420;
wire            n9421;
wire      [7:0] n9422;
wire            n9423;
wire            n9424;
wire            n9425;
wire            n9426;
wire            n9427;
wire      [7:0] n9428;
wire            n9429;
wire            n943;
wire            n9430;
wire            n9431;
wire            n9432;
wire            n9433;
wire      [7:0] n9434;
wire            n9435;
wire            n9436;
wire            n9437;
wire            n9438;
wire            n9439;
wire            n944;
wire      [7:0] n9440;
wire            n9441;
wire            n9442;
wire            n9443;
wire            n9444;
wire            n9445;
wire      [7:0] n9446;
wire            n9447;
wire            n9448;
wire            n9449;
wire            n945;
wire            n9450;
wire            n9451;
wire      [7:0] n9452;
wire            n9453;
wire            n9454;
wire            n9455;
wire            n9456;
wire            n9457;
wire      [7:0] n9458;
wire            n9459;
wire            n946;
wire            n9460;
wire            n9461;
wire            n9462;
wire            n9463;
wire      [7:0] n9464;
wire            n9465;
wire            n9466;
wire            n9467;
wire            n9468;
wire            n9469;
wire            n947;
wire      [7:0] n9470;
wire            n9471;
wire            n9472;
wire            n9473;
wire            n9474;
wire            n9475;
wire      [7:0] n9476;
wire            n9477;
wire            n9478;
wire            n9479;
wire            n948;
wire            n9480;
wire            n9481;
wire      [7:0] n9482;
wire            n9483;
wire            n9484;
wire            n9485;
wire            n9486;
wire            n9487;
wire      [7:0] n9488;
wire            n9489;
wire            n949;
wire            n9490;
wire            n9491;
wire            n9492;
wire            n9493;
wire      [7:0] n9494;
wire            n9495;
wire            n9496;
wire            n9497;
wire            n9498;
wire            n9499;
wire            n950;
wire      [7:0] n9500;
wire            n9501;
wire            n9502;
wire            n9503;
wire            n9504;
wire            n9505;
wire      [7:0] n9506;
wire            n9507;
wire            n9508;
wire            n9509;
wire            n951;
wire            n9510;
wire            n9511;
wire      [7:0] n9512;
wire            n9513;
wire            n9514;
wire            n9515;
wire            n9516;
wire            n9517;
wire      [7:0] n9518;
wire            n9519;
wire            n952;
wire            n9520;
wire            n9521;
wire            n9522;
wire            n9523;
wire      [7:0] n9524;
wire            n9525;
wire            n9526;
wire            n9527;
wire            n9528;
wire            n9529;
wire            n953;
wire      [7:0] n9530;
wire            n9531;
wire            n9532;
wire            n9533;
wire            n9534;
wire            n9535;
wire      [7:0] n9536;
wire            n9537;
wire            n9538;
wire            n9539;
wire            n954;
wire            n9540;
wire            n9541;
wire      [7:0] n9542;
wire            n9543;
wire            n9544;
wire            n9545;
wire            n9546;
wire            n9547;
wire      [7:0] n9548;
wire            n9549;
wire            n955;
wire            n9550;
wire            n9551;
wire            n9552;
wire            n9553;
wire      [7:0] n9554;
wire            n9555;
wire            n9556;
wire            n9557;
wire            n9558;
wire            n9559;
wire            n956;
wire      [7:0] n9560;
wire            n9561;
wire            n9562;
wire            n9563;
wire            n9564;
wire            n9565;
wire      [7:0] n9566;
wire            n9567;
wire            n9568;
wire            n9569;
wire            n957;
wire            n9570;
wire            n9571;
wire      [7:0] n9572;
wire            n9573;
wire            n9574;
wire            n9575;
wire            n9576;
wire            n9577;
wire      [7:0] n9578;
wire            n9579;
wire            n958;
wire            n9580;
wire            n9581;
wire            n9582;
wire            n9583;
wire      [7:0] n9584;
wire            n9585;
wire            n9586;
wire            n9587;
wire            n9588;
wire            n9589;
wire            n959;
wire      [7:0] n9590;
wire            n9591;
wire            n9592;
wire            n9593;
wire            n9594;
wire            n9595;
wire      [7:0] n9596;
wire            n9597;
wire            n9598;
wire            n9599;
wire            n96;
wire            n960;
wire            n9600;
wire            n9601;
wire      [7:0] n9602;
wire            n9603;
wire            n9604;
wire            n9605;
wire            n9606;
wire            n9607;
wire      [7:0] n9608;
wire            n9609;
wire            n961;
wire            n9610;
wire            n9611;
wire            n9612;
wire            n9613;
wire      [7:0] n9614;
wire            n9615;
wire            n9616;
wire            n9617;
wire            n9618;
wire            n9619;
wire            n962;
wire      [7:0] n9620;
wire            n9621;
wire            n9622;
wire            n9623;
wire            n9624;
wire            n9625;
wire      [7:0] n9626;
wire            n9627;
wire            n9628;
wire            n9629;
wire            n963;
wire            n9630;
wire            n9631;
wire      [7:0] n9632;
wire            n9633;
wire            n9634;
wire            n9635;
wire            n9636;
wire            n9637;
wire      [7:0] n9638;
wire            n9639;
wire            n964;
wire            n9640;
wire            n9641;
wire            n9642;
wire            n9643;
wire      [7:0] n9644;
wire            n9645;
wire            n9646;
wire            n9647;
wire            n9648;
wire            n9649;
wire            n965;
wire      [7:0] n9650;
wire            n9651;
wire            n9652;
wire            n9653;
wire            n9654;
wire            n9655;
wire      [7:0] n9656;
wire            n9657;
wire            n9658;
wire            n9659;
wire            n966;
wire            n9660;
wire            n9661;
wire      [7:0] n9662;
wire            n9663;
wire            n9664;
wire            n9665;
wire            n9666;
wire            n9667;
wire      [7:0] n9668;
wire            n9669;
wire            n967;
wire            n9670;
wire            n9671;
wire            n9672;
wire            n9673;
wire      [7:0] n9674;
wire            n9675;
wire            n9676;
wire            n9677;
wire            n9678;
wire            n9679;
wire            n968;
wire      [7:0] n9680;
wire            n9681;
wire            n9682;
wire            n9683;
wire            n9684;
wire            n9685;
wire      [7:0] n9686;
wire            n9687;
wire            n9688;
wire            n9689;
wire            n969;
wire            n9690;
wire            n9691;
wire      [7:0] n9692;
wire            n9693;
wire            n9694;
wire            n9695;
wire            n9696;
wire            n9697;
wire      [7:0] n9698;
wire            n9699;
wire            n970;
wire            n9700;
wire            n9701;
wire            n9702;
wire            n9703;
wire      [7:0] n9704;
wire            n9705;
wire            n9706;
wire            n9707;
wire            n9708;
wire            n9709;
wire            n971;
wire      [7:0] n9710;
wire            n9711;
wire            n9712;
wire            n9713;
wire            n9714;
wire            n9715;
wire      [7:0] n9716;
wire            n9717;
wire            n9718;
wire            n9719;
wire            n972;
wire            n9720;
wire            n9721;
wire      [7:0] n9722;
wire            n9723;
wire            n9724;
wire            n9725;
wire            n9726;
wire            n9727;
wire      [7:0] n9728;
wire            n9729;
wire            n973;
wire            n9730;
wire            n9731;
wire            n9732;
wire            n9733;
wire      [7:0] n9734;
wire            n9735;
wire            n9736;
wire            n9737;
wire            n9738;
wire            n9739;
wire            n974;
wire      [7:0] n9740;
wire            n9741;
wire            n9742;
wire            n9743;
wire            n9744;
wire            n9745;
wire      [7:0] n9746;
wire            n9747;
wire            n9748;
wire            n9749;
wire            n975;
wire            n9750;
wire            n9751;
wire      [7:0] n9752;
wire            n9753;
wire            n9754;
wire            n9755;
wire            n9756;
wire            n9757;
wire      [7:0] n9758;
wire            n9759;
wire            n976;
wire            n9760;
wire            n9761;
wire            n9762;
wire            n9763;
wire      [7:0] n9764;
wire            n9765;
wire            n9766;
wire            n9767;
wire            n9768;
wire            n9769;
wire            n977;
wire      [7:0] n9770;
wire            n9771;
wire            n9772;
wire            n9773;
wire            n9774;
wire            n9775;
wire      [7:0] n9776;
wire            n9777;
wire            n9778;
wire            n9779;
wire            n978;
wire            n9780;
wire            n9781;
wire      [7:0] n9782;
wire            n9783;
wire            n9784;
wire            n9785;
wire            n9786;
wire            n9787;
wire      [7:0] n9788;
wire            n9789;
wire            n979;
wire            n9790;
wire            n9791;
wire            n9792;
wire            n9793;
wire      [7:0] n9794;
wire            n9795;
wire            n9796;
wire            n9797;
wire            n9798;
wire            n9799;
wire            n98;
wire            n980;
wire      [7:0] n9800;
wire            n9801;
wire            n9802;
wire            n9803;
wire            n9804;
wire            n9805;
wire      [7:0] n9806;
wire            n9807;
wire            n9808;
wire            n9809;
wire            n981;
wire            n9810;
wire            n9811;
wire      [7:0] n9812;
wire            n9813;
wire            n9814;
wire            n9815;
wire            n9816;
wire            n9817;
wire      [7:0] n9818;
wire            n9819;
wire            n982;
wire            n9820;
wire            n9821;
wire            n9822;
wire            n9823;
wire      [7:0] n9824;
wire            n9825;
wire            n9826;
wire            n9827;
wire            n9828;
wire            n9829;
wire            n983;
wire      [7:0] n9830;
wire            n9831;
wire            n9832;
wire            n9833;
wire            n9834;
wire            n9835;
wire      [7:0] n9836;
wire            n9837;
wire            n9838;
wire            n9839;
wire            n984;
wire            n9840;
wire            n9841;
wire      [7:0] n9842;
wire            n9843;
wire            n9844;
wire            n9845;
wire            n9846;
wire            n9847;
wire      [7:0] n9848;
wire            n9849;
wire            n985;
wire            n9850;
wire            n9851;
wire            n9852;
wire            n9853;
wire      [7:0] n9854;
wire            n9855;
wire            n9856;
wire            n9857;
wire            n9858;
wire            n9859;
wire            n986;
wire      [7:0] n9860;
wire            n9861;
wire            n9862;
wire            n9863;
wire            n9864;
wire            n9865;
wire      [7:0] n9866;
wire            n9867;
wire            n9868;
wire            n9869;
wire            n987;
wire            n9870;
wire            n9871;
wire      [7:0] n9872;
wire            n9873;
wire            n9874;
wire            n9875;
wire            n9876;
wire            n9877;
wire      [7:0] n9878;
wire            n9879;
wire            n988;
wire            n9880;
wire            n9881;
wire            n9882;
wire            n9883;
wire      [7:0] n9884;
wire            n9885;
wire            n9886;
wire            n9887;
wire            n9888;
wire            n9889;
wire            n989;
wire      [7:0] n9890;
wire            n9891;
wire            n9892;
wire            n9893;
wire            n9894;
wire            n9895;
wire      [7:0] n9896;
wire            n9897;
wire            n9898;
wire            n9899;
wire            n990;
wire            n9900;
wire            n9901;
wire      [7:0] n9902;
wire            n9903;
wire            n9904;
wire            n9905;
wire            n9906;
wire            n9907;
wire      [7:0] n9908;
wire            n9909;
wire            n991;
wire            n9910;
wire            n9911;
wire            n9912;
wire            n9913;
wire      [7:0] n9914;
wire            n9915;
wire            n9916;
wire            n9917;
wire            n9918;
wire            n9919;
wire            n992;
wire      [7:0] n9920;
wire            n9921;
wire            n9922;
wire            n9923;
wire            n9924;
wire            n9925;
wire      [7:0] n9926;
wire            n9927;
wire            n9928;
wire            n9929;
wire            n993;
wire            n9930;
wire            n9931;
wire      [7:0] n9932;
wire            n9933;
wire            n9934;
wire            n9935;
wire            n9936;
wire            n9937;
wire      [7:0] n9938;
wire            n9939;
wire            n994;
wire            n9940;
wire            n9941;
wire            n9942;
wire            n9943;
wire      [7:0] n9944;
wire            n9945;
wire            n9946;
wire            n9947;
wire            n9948;
wire            n9949;
wire            n995;
wire      [7:0] n9950;
wire            n9951;
wire            n9952;
wire            n9953;
wire            n9954;
wire            n9955;
wire      [7:0] n9956;
wire            n9957;
wire            n9958;
wire            n9959;
wire            n996;
wire            n9960;
wire            n9961;
wire      [7:0] n9962;
wire            n9963;
wire            n9964;
wire            n9965;
wire            n9966;
wire            n9967;
wire      [7:0] n9968;
wire            n9969;
wire            n997;
wire            n9970;
wire            n9971;
wire            n9972;
wire            n9973;
wire      [7:0] n9974;
wire            n9975;
wire            n9976;
wire            n9977;
wire            n9978;
wire            n9979;
wire            n998;
wire      [7:0] n9980;
wire            n9981;
wire            n9982;
wire            n9983;
wire            n9984;
wire            n9985;
wire      [7:0] n9986;
wire            n9987;
wire            n9988;
wire            n9989;
wire            n999;
wire            n9990;
wire            n9991;
wire      [7:0] n9992;
wire            n9993;
wire            n9994;
wire            n9995;
wire            n9996;
wire            n9997;
wire      [7:0] n9998;
wire            n9999;
wire      [7:0] nondet_des1_func_n3936;
wire            nondet_desCy_func_n3988;
wire      [7:0] nondet_des_acc_func_n3499;
wire      [7:0] nondet_div_des1_n4958;
wire      [7:0] nondet_div_des2_n4955;
wire      [7:0] nondet_mul_des1_n4947;
wire      [7:0] nondet_mul_des2_n4944;
wire      [7:0] nondet_psw_next_func_n3704;
wire      [7:0] op2;
wire      [7:0] op3;
wire            p;
wire     [15:0] pc;
wire      [1:0] psw_set;
wire      [2:0] ram_rd_sel;
wire      [2:0] ram_wr_sel;
wire      [7:0] rd_addr;
wire            rst;
wire      [2:0] src_sel1;
wire      [1:0] src_sel2;
wire            src_sel3;
wire            wr;
wire      [7:0] wr_addr;
wire            wr_ind;
wire      [1:0] wr_sfr;
assign __ILA_DATAPATH_valid__ = 1'b1 ;
assign bv_4_7_n0 = 4'h7 ;
assign n1 =  ( alu_op ) == ( bv_4_7_n0 )  ;
assign __ILA_DATAPATH_decode_of_alu_and__ = n1 ;
assign __ILA_DATAPATH_acc_decode__[0] = __ILA_DATAPATH_decode_of_alu_and__ ;
assign bv_4_14_n2 = 4'he ;
assign n3 =  ( alu_op ) == ( bv_4_14_n2 )  ;
assign __ILA_DATAPATH_decode_of_alu_inc__ = n3 ;
assign __ILA_DATAPATH_acc_decode__[1] = __ILA_DATAPATH_decode_of_alu_inc__ ;
assign bv_4_6_n4 = 4'h6 ;
assign n5 =  ( alu_op ) == ( bv_4_6_n4 )  ;
assign __ILA_DATAPATH_decode_of_alu_not__ = n5 ;
assign __ILA_DATAPATH_acc_decode__[2] = __ILA_DATAPATH_decode_of_alu_not__ ;
assign bv_4_5_n6 = 4'h5 ;
assign n7 =  ( alu_op ) == ( bv_4_5_n6 )  ;
assign __ILA_DATAPATH_decode_of_alu_da__ = n7 ;
assign __ILA_DATAPATH_acc_decode__[3] = __ILA_DATAPATH_decode_of_alu_da__ ;
assign bv_4_3_n8 = 4'h3 ;
assign n9 =  ( alu_op ) == ( bv_4_3_n8 )  ;
assign __ILA_DATAPATH_decode_of_alu_mul__ = n9 ;
assign __ILA_DATAPATH_acc_decode__[4] = __ILA_DATAPATH_decode_of_alu_mul__ ;
assign bv_4_4_n10 = 4'h4 ;
assign n11 =  ( alu_op ) == ( bv_4_4_n10 )  ;
assign __ILA_DATAPATH_decode_of_alu_div__ = n11 ;
assign __ILA_DATAPATH_acc_decode__[5] = __ILA_DATAPATH_decode_of_alu_div__ ;
assign bv_4_2_n12 = 4'h2 ;
assign n13 =  ( alu_op ) == ( bv_4_2_n12 )  ;
assign __ILA_DATAPATH_decode_of_alu_sub__ = n13 ;
assign __ILA_DATAPATH_acc_decode__[6] = __ILA_DATAPATH_decode_of_alu_sub__ ;
assign bv_4_9_n14 = 4'h9 ;
assign n15 =  ( alu_op ) == ( bv_4_9_n14 )  ;
assign __ILA_DATAPATH_decode_of_alu_or__ = n15 ;
assign __ILA_DATAPATH_acc_decode__[7] = __ILA_DATAPATH_decode_of_alu_or__ ;
assign bv_4_10_n16 = 4'ha ;
assign n17 =  ( alu_op ) == ( bv_4_10_n16 )  ;
assign __ILA_DATAPATH_decode_of_alu_rl__ = n17 ;
assign __ILA_DATAPATH_acc_decode__[8] = __ILA_DATAPATH_decode_of_alu_rl__ ;
assign bv_4_11_n18 = 4'hb ;
assign n19 =  ( alu_op ) == ( bv_4_11_n18 )  ;
assign __ILA_DATAPATH_decode_of_alu_rlc__ = n19 ;
assign __ILA_DATAPATH_acc_decode__[9] = __ILA_DATAPATH_decode_of_alu_rlc__ ;
assign bv_4_12_n20 = 4'hc ;
assign n21 =  ( alu_op ) == ( bv_4_12_n20 )  ;
assign __ILA_DATAPATH_decode_of_alu_rr__ = n21 ;
assign __ILA_DATAPATH_acc_decode__[10] = __ILA_DATAPATH_decode_of_alu_rr__ ;
assign bv_4_13_n22 = 4'hd ;
assign n23 =  ( alu_op ) == ( bv_4_13_n22 )  ;
assign __ILA_DATAPATH_decode_of_alu_rrc__ = n23 ;
assign __ILA_DATAPATH_acc_decode__[11] = __ILA_DATAPATH_decode_of_alu_rrc__ ;
assign bv_4_15_n24 = 4'hf ;
assign n25 =  ( alu_op ) == ( bv_4_15_n24 )  ;
assign __ILA_DATAPATH_decode_of_alu_xch__ = n25 ;
assign __ILA_DATAPATH_acc_decode__[12] = __ILA_DATAPATH_decode_of_alu_xch__ ;
assign bv_4_8_n26 = 4'h8 ;
assign n27 =  ( alu_op ) == ( bv_4_8_n26 )  ;
assign __ILA_DATAPATH_decode_of_alu_xor__ = n27 ;
assign __ILA_DATAPATH_acc_decode__[13] = __ILA_DATAPATH_decode_of_alu_xor__ ;
assign bv_4_1_n28 = 4'h1 ;
assign n29 =  ( alu_op ) == ( bv_4_1_n28 )  ;
assign __ILA_DATAPATH_decode_of_alu_add__ = n29 ;
assign __ILA_DATAPATH_acc_decode__[14] = __ILA_DATAPATH_decode_of_alu_add__ ;
assign bv_4_0_n30 = 4'h0 ;
assign n31 =  ( alu_op ) == ( bv_4_0_n30 )  ;
assign __ILA_DATAPATH_decode_of_read_data__ = n31 ;
assign __ILA_DATAPATH_acc_decode__[15] = __ILA_DATAPATH_decode_of_read_data__ ;
assign n32 =  ( wr ) == ( 1'b0 )  ;
assign __ILA_DATAPATH_decode_of_no_wr__ = n32 ;
assign __ILA_DATAPATH_acc_decode__[16] = __ILA_DATAPATH_decode_of_no_wr__ ;
assign n33 = wr_addr[7:7] ;
assign bv_1_1_n34 = 1'h1 ;
assign n35 =  ( n33 ) == ( bv_1_1_n34 )  ;
assign n36 =  ( wr_ind ) == ( 1'b0 )  ;
assign n37 =  ( n35 ) & (n36 )  ;
assign n38 =  ( wr ) & (n37 )  ;
assign __ILA_DATAPATH_decode_of_wr_sfr__ = n38 ;
assign __ILA_DATAPATH_acc_decode__[17] = __ILA_DATAPATH_decode_of_wr_sfr__ ;
assign n39 =  ( wr ) & (wr_ind )  ;
assign __ILA_DATAPATH_decode_of_wr_ram__ = n39 ;
assign __ILA_DATAPATH_acc_decode__[18] = __ILA_DATAPATH_decode_of_wr_ram__ ;
assign n40 =  ( wr_ind ) == ( 1'b0 )  ;
assign n41 =  ( wr ) & (n40 )  ;
assign n42 = wr_addr[7:7] ;
assign n43 =  ( n42 ) == ( bv_1_1_n34 )  ;
assign n44 = wr_addr[6:3] ;
assign n45 =  { ( bv_1_1_n34 ) , ( n44 ) }  ;
assign bv_3_0_n46 = 3'h0 ;
assign n47 =  { ( n45 ) , ( bv_3_0_n46 ) }  ;
assign n48 = wr_addr[6:3] ;
assign n49 =  { ( bv_4_2_n12 ) , ( n48 ) }  ;
assign n50 =  ( n43 ) ? ( n47 ) : ( n49 ) ;
assign n51 =  ( bit_addr_r ) ? ( n50 ) : ( wr_addr ) ;
assign n52 = n51[7:7] ;
assign bv_1_0_n53 = 1'h0 ;
assign n54 =  ( n52 ) == ( bv_1_0_n53 )  ;
assign n55 =  ( n41 ) & (n54 )  ;
assign __ILA_DATAPATH_decode_of_wr_sfr_ram__ = n55 ;
assign __ILA_DATAPATH_acc_decode__[19] = __ILA_DATAPATH_decode_of_wr_sfr_ram__ ;
assign n56 = rd_addr[2:0] ;
assign n57 = rd_addr[2:0] ;
assign n58 = rd_addr[2:0] ;
assign n59 = rd_addr[2:0] ;
assign n60 = rd_addr[2:0] ;
assign n61 = rd_addr[7:7] ;
assign n62 =  ( n61 ) == ( bv_1_1_n34 )  ;
assign n63 = rd_addr[6:3] ;
assign n64 =  { ( bv_1_1_n34 ) , ( n63 ) }  ;
assign n65 =  { ( n64 ) , ( bv_3_0_n46 ) }  ;
assign n66 = rd_addr[6:3] ;
assign n67 =  { ( bv_4_2_n12 ) , ( n66 ) }  ;
assign n68 =  ( n62 ) ? ( n65 ) : ( n67 ) ;
assign bv_8_0_n69 = 8'h0 ;
assign n70 =  ( n68 ) == ( bv_8_0_n69 )  ;
assign bv_8_1_n71 = 8'h1 ;
assign n72 =  ( n68 ) == ( bv_8_1_n71 )  ;
assign bv_8_2_n73 = 8'h2 ;
assign n74 =  ( n68 ) == ( bv_8_2_n73 )  ;
assign bv_8_3_n75 = 8'h3 ;
assign n76 =  ( n68 ) == ( bv_8_3_n75 )  ;
assign bv_8_4_n77 = 8'h4 ;
assign n78 =  ( n68 ) == ( bv_8_4_n77 )  ;
assign bv_8_5_n79 = 8'h5 ;
assign n80 =  ( n68 ) == ( bv_8_5_n79 )  ;
assign bv_8_6_n81 = 8'h6 ;
assign n82 =  ( n68 ) == ( bv_8_6_n81 )  ;
assign bv_8_7_n83 = 8'h7 ;
assign n84 =  ( n68 ) == ( bv_8_7_n83 )  ;
assign bv_8_8_n85 = 8'h8 ;
assign n86 =  ( n68 ) == ( bv_8_8_n85 )  ;
assign bv_8_9_n87 = 8'h9 ;
assign n88 =  ( n68 ) == ( bv_8_9_n87 )  ;
assign bv_8_10_n89 = 8'ha ;
assign n90 =  ( n68 ) == ( bv_8_10_n89 )  ;
assign bv_8_11_n91 = 8'hb ;
assign n92 =  ( n68 ) == ( bv_8_11_n91 )  ;
assign bv_8_12_n93 = 8'hc ;
assign n94 =  ( n68 ) == ( bv_8_12_n93 )  ;
assign bv_8_13_n95 = 8'hd ;
assign n96 =  ( n68 ) == ( bv_8_13_n95 )  ;
assign bv_8_14_n97 = 8'he ;
assign n98 =  ( n68 ) == ( bv_8_14_n97 )  ;
assign bv_8_15_n99 = 8'hf ;
assign n100 =  ( n68 ) == ( bv_8_15_n99 )  ;
assign bv_8_16_n101 = 8'h10 ;
assign n102 =  ( n68 ) == ( bv_8_16_n101 )  ;
assign bv_8_17_n103 = 8'h11 ;
assign n104 =  ( n68 ) == ( bv_8_17_n103 )  ;
assign bv_8_18_n105 = 8'h12 ;
assign n106 =  ( n68 ) == ( bv_8_18_n105 )  ;
assign bv_8_19_n107 = 8'h13 ;
assign n108 =  ( n68 ) == ( bv_8_19_n107 )  ;
assign bv_8_20_n109 = 8'h14 ;
assign n110 =  ( n68 ) == ( bv_8_20_n109 )  ;
assign bv_8_21_n111 = 8'h15 ;
assign n112 =  ( n68 ) == ( bv_8_21_n111 )  ;
assign bv_8_22_n113 = 8'h16 ;
assign n114 =  ( n68 ) == ( bv_8_22_n113 )  ;
assign bv_8_23_n115 = 8'h17 ;
assign n116 =  ( n68 ) == ( bv_8_23_n115 )  ;
assign bv_8_24_n117 = 8'h18 ;
assign n118 =  ( n68 ) == ( bv_8_24_n117 )  ;
assign bv_8_25_n119 = 8'h19 ;
assign n120 =  ( n68 ) == ( bv_8_25_n119 )  ;
assign bv_8_26_n121 = 8'h1a ;
assign n122 =  ( n68 ) == ( bv_8_26_n121 )  ;
assign bv_8_27_n123 = 8'h1b ;
assign n124 =  ( n68 ) == ( bv_8_27_n123 )  ;
assign bv_8_28_n125 = 8'h1c ;
assign n126 =  ( n68 ) == ( bv_8_28_n125 )  ;
assign bv_8_29_n127 = 8'h1d ;
assign n128 =  ( n68 ) == ( bv_8_29_n127 )  ;
assign bv_8_30_n129 = 8'h1e ;
assign n130 =  ( n68 ) == ( bv_8_30_n129 )  ;
assign bv_8_31_n131 = 8'h1f ;
assign n132 =  ( n68 ) == ( bv_8_31_n131 )  ;
assign bv_8_32_n133 = 8'h20 ;
assign n134 =  ( n68 ) == ( bv_8_32_n133 )  ;
assign bv_8_33_n135 = 8'h21 ;
assign n136 =  ( n68 ) == ( bv_8_33_n135 )  ;
assign bv_8_34_n137 = 8'h22 ;
assign n138 =  ( n68 ) == ( bv_8_34_n137 )  ;
assign bv_8_35_n139 = 8'h23 ;
assign n140 =  ( n68 ) == ( bv_8_35_n139 )  ;
assign bv_8_36_n141 = 8'h24 ;
assign n142 =  ( n68 ) == ( bv_8_36_n141 )  ;
assign bv_8_37_n143 = 8'h25 ;
assign n144 =  ( n68 ) == ( bv_8_37_n143 )  ;
assign bv_8_38_n145 = 8'h26 ;
assign n146 =  ( n68 ) == ( bv_8_38_n145 )  ;
assign bv_8_39_n147 = 8'h27 ;
assign n148 =  ( n68 ) == ( bv_8_39_n147 )  ;
assign bv_8_40_n149 = 8'h28 ;
assign n150 =  ( n68 ) == ( bv_8_40_n149 )  ;
assign bv_8_41_n151 = 8'h29 ;
assign n152 =  ( n68 ) == ( bv_8_41_n151 )  ;
assign bv_8_42_n153 = 8'h2a ;
assign n154 =  ( n68 ) == ( bv_8_42_n153 )  ;
assign bv_8_43_n155 = 8'h2b ;
assign n156 =  ( n68 ) == ( bv_8_43_n155 )  ;
assign bv_8_44_n157 = 8'h2c ;
assign n158 =  ( n68 ) == ( bv_8_44_n157 )  ;
assign bv_8_45_n159 = 8'h2d ;
assign n160 =  ( n68 ) == ( bv_8_45_n159 )  ;
assign bv_8_46_n161 = 8'h2e ;
assign n162 =  ( n68 ) == ( bv_8_46_n161 )  ;
assign bv_8_47_n163 = 8'h2f ;
assign n164 =  ( n68 ) == ( bv_8_47_n163 )  ;
assign bv_8_48_n165 = 8'h30 ;
assign n166 =  ( n68 ) == ( bv_8_48_n165 )  ;
assign bv_8_49_n167 = 8'h31 ;
assign n168 =  ( n68 ) == ( bv_8_49_n167 )  ;
assign bv_8_50_n169 = 8'h32 ;
assign n170 =  ( n68 ) == ( bv_8_50_n169 )  ;
assign bv_8_51_n171 = 8'h33 ;
assign n172 =  ( n68 ) == ( bv_8_51_n171 )  ;
assign bv_8_52_n173 = 8'h34 ;
assign n174 =  ( n68 ) == ( bv_8_52_n173 )  ;
assign bv_8_53_n175 = 8'h35 ;
assign n176 =  ( n68 ) == ( bv_8_53_n175 )  ;
assign bv_8_54_n177 = 8'h36 ;
assign n178 =  ( n68 ) == ( bv_8_54_n177 )  ;
assign bv_8_55_n179 = 8'h37 ;
assign n180 =  ( n68 ) == ( bv_8_55_n179 )  ;
assign bv_8_56_n181 = 8'h38 ;
assign n182 =  ( n68 ) == ( bv_8_56_n181 )  ;
assign bv_8_57_n183 = 8'h39 ;
assign n184 =  ( n68 ) == ( bv_8_57_n183 )  ;
assign bv_8_58_n185 = 8'h3a ;
assign n186 =  ( n68 ) == ( bv_8_58_n185 )  ;
assign bv_8_59_n187 = 8'h3b ;
assign n188 =  ( n68 ) == ( bv_8_59_n187 )  ;
assign bv_8_60_n189 = 8'h3c ;
assign n190 =  ( n68 ) == ( bv_8_60_n189 )  ;
assign bv_8_61_n191 = 8'h3d ;
assign n192 =  ( n68 ) == ( bv_8_61_n191 )  ;
assign bv_8_62_n193 = 8'h3e ;
assign n194 =  ( n68 ) == ( bv_8_62_n193 )  ;
assign bv_8_63_n195 = 8'h3f ;
assign n196 =  ( n68 ) == ( bv_8_63_n195 )  ;
assign bv_8_64_n197 = 8'h40 ;
assign n198 =  ( n68 ) == ( bv_8_64_n197 )  ;
assign bv_8_65_n199 = 8'h41 ;
assign n200 =  ( n68 ) == ( bv_8_65_n199 )  ;
assign bv_8_66_n201 = 8'h42 ;
assign n202 =  ( n68 ) == ( bv_8_66_n201 )  ;
assign bv_8_67_n203 = 8'h43 ;
assign n204 =  ( n68 ) == ( bv_8_67_n203 )  ;
assign bv_8_68_n205 = 8'h44 ;
assign n206 =  ( n68 ) == ( bv_8_68_n205 )  ;
assign bv_8_69_n207 = 8'h45 ;
assign n208 =  ( n68 ) == ( bv_8_69_n207 )  ;
assign bv_8_70_n209 = 8'h46 ;
assign n210 =  ( n68 ) == ( bv_8_70_n209 )  ;
assign bv_8_71_n211 = 8'h47 ;
assign n212 =  ( n68 ) == ( bv_8_71_n211 )  ;
assign bv_8_72_n213 = 8'h48 ;
assign n214 =  ( n68 ) == ( bv_8_72_n213 )  ;
assign bv_8_73_n215 = 8'h49 ;
assign n216 =  ( n68 ) == ( bv_8_73_n215 )  ;
assign bv_8_74_n217 = 8'h4a ;
assign n218 =  ( n68 ) == ( bv_8_74_n217 )  ;
assign bv_8_75_n219 = 8'h4b ;
assign n220 =  ( n68 ) == ( bv_8_75_n219 )  ;
assign bv_8_76_n221 = 8'h4c ;
assign n222 =  ( n68 ) == ( bv_8_76_n221 )  ;
assign bv_8_77_n223 = 8'h4d ;
assign n224 =  ( n68 ) == ( bv_8_77_n223 )  ;
assign bv_8_78_n225 = 8'h4e ;
assign n226 =  ( n68 ) == ( bv_8_78_n225 )  ;
assign bv_8_79_n227 = 8'h4f ;
assign n228 =  ( n68 ) == ( bv_8_79_n227 )  ;
assign bv_8_80_n229 = 8'h50 ;
assign n230 =  ( n68 ) == ( bv_8_80_n229 )  ;
assign bv_8_81_n231 = 8'h51 ;
assign n232 =  ( n68 ) == ( bv_8_81_n231 )  ;
assign bv_8_82_n233 = 8'h52 ;
assign n234 =  ( n68 ) == ( bv_8_82_n233 )  ;
assign bv_8_83_n235 = 8'h53 ;
assign n236 =  ( n68 ) == ( bv_8_83_n235 )  ;
assign bv_8_84_n237 = 8'h54 ;
assign n238 =  ( n68 ) == ( bv_8_84_n237 )  ;
assign bv_8_85_n239 = 8'h55 ;
assign n240 =  ( n68 ) == ( bv_8_85_n239 )  ;
assign bv_8_86_n241 = 8'h56 ;
assign n242 =  ( n68 ) == ( bv_8_86_n241 )  ;
assign bv_8_87_n243 = 8'h57 ;
assign n244 =  ( n68 ) == ( bv_8_87_n243 )  ;
assign bv_8_88_n245 = 8'h58 ;
assign n246 =  ( n68 ) == ( bv_8_88_n245 )  ;
assign bv_8_89_n247 = 8'h59 ;
assign n248 =  ( n68 ) == ( bv_8_89_n247 )  ;
assign bv_8_90_n249 = 8'h5a ;
assign n250 =  ( n68 ) == ( bv_8_90_n249 )  ;
assign bv_8_91_n251 = 8'h5b ;
assign n252 =  ( n68 ) == ( bv_8_91_n251 )  ;
assign bv_8_92_n253 = 8'h5c ;
assign n254 =  ( n68 ) == ( bv_8_92_n253 )  ;
assign bv_8_93_n255 = 8'h5d ;
assign n256 =  ( n68 ) == ( bv_8_93_n255 )  ;
assign bv_8_94_n257 = 8'h5e ;
assign n258 =  ( n68 ) == ( bv_8_94_n257 )  ;
assign bv_8_95_n259 = 8'h5f ;
assign n260 =  ( n68 ) == ( bv_8_95_n259 )  ;
assign bv_8_96_n261 = 8'h60 ;
assign n262 =  ( n68 ) == ( bv_8_96_n261 )  ;
assign bv_8_97_n263 = 8'h61 ;
assign n264 =  ( n68 ) == ( bv_8_97_n263 )  ;
assign bv_8_98_n265 = 8'h62 ;
assign n266 =  ( n68 ) == ( bv_8_98_n265 )  ;
assign bv_8_99_n267 = 8'h63 ;
assign n268 =  ( n68 ) == ( bv_8_99_n267 )  ;
assign bv_8_100_n269 = 8'h64 ;
assign n270 =  ( n68 ) == ( bv_8_100_n269 )  ;
assign bv_8_101_n271 = 8'h65 ;
assign n272 =  ( n68 ) == ( bv_8_101_n271 )  ;
assign bv_8_102_n273 = 8'h66 ;
assign n274 =  ( n68 ) == ( bv_8_102_n273 )  ;
assign bv_8_103_n275 = 8'h67 ;
assign n276 =  ( n68 ) == ( bv_8_103_n275 )  ;
assign bv_8_104_n277 = 8'h68 ;
assign n278 =  ( n68 ) == ( bv_8_104_n277 )  ;
assign bv_8_105_n279 = 8'h69 ;
assign n280 =  ( n68 ) == ( bv_8_105_n279 )  ;
assign bv_8_106_n281 = 8'h6a ;
assign n282 =  ( n68 ) == ( bv_8_106_n281 )  ;
assign bv_8_107_n283 = 8'h6b ;
assign n284 =  ( n68 ) == ( bv_8_107_n283 )  ;
assign bv_8_108_n285 = 8'h6c ;
assign n286 =  ( n68 ) == ( bv_8_108_n285 )  ;
assign bv_8_109_n287 = 8'h6d ;
assign n288 =  ( n68 ) == ( bv_8_109_n287 )  ;
assign bv_8_110_n289 = 8'h6e ;
assign n290 =  ( n68 ) == ( bv_8_110_n289 )  ;
assign bv_8_111_n291 = 8'h6f ;
assign n292 =  ( n68 ) == ( bv_8_111_n291 )  ;
assign bv_8_112_n293 = 8'h70 ;
assign n294 =  ( n68 ) == ( bv_8_112_n293 )  ;
assign bv_8_113_n295 = 8'h71 ;
assign n296 =  ( n68 ) == ( bv_8_113_n295 )  ;
assign bv_8_114_n297 = 8'h72 ;
assign n298 =  ( n68 ) == ( bv_8_114_n297 )  ;
assign bv_8_115_n299 = 8'h73 ;
assign n300 =  ( n68 ) == ( bv_8_115_n299 )  ;
assign bv_8_116_n301 = 8'h74 ;
assign n302 =  ( n68 ) == ( bv_8_116_n301 )  ;
assign bv_8_117_n303 = 8'h75 ;
assign n304 =  ( n68 ) == ( bv_8_117_n303 )  ;
assign bv_8_118_n305 = 8'h76 ;
assign n306 =  ( n68 ) == ( bv_8_118_n305 )  ;
assign bv_8_119_n307 = 8'h77 ;
assign n308 =  ( n68 ) == ( bv_8_119_n307 )  ;
assign bv_8_120_n309 = 8'h78 ;
assign n310 =  ( n68 ) == ( bv_8_120_n309 )  ;
assign bv_8_121_n311 = 8'h79 ;
assign n312 =  ( n68 ) == ( bv_8_121_n311 )  ;
assign bv_8_122_n313 = 8'h7a ;
assign n314 =  ( n68 ) == ( bv_8_122_n313 )  ;
assign bv_8_123_n315 = 8'h7b ;
assign n316 =  ( n68 ) == ( bv_8_123_n315 )  ;
assign bv_8_124_n317 = 8'h7c ;
assign n318 =  ( n68 ) == ( bv_8_124_n317 )  ;
assign bv_8_125_n319 = 8'h7d ;
assign n320 =  ( n68 ) == ( bv_8_125_n319 )  ;
assign bv_8_126_n321 = 8'h7e ;
assign n322 =  ( n68 ) == ( bv_8_126_n321 )  ;
assign bv_8_127_n323 = 8'h7f ;
assign n324 =  ( n68 ) == ( bv_8_127_n323 )  ;
assign bv_8_128_n325 = 8'h80 ;
assign n326 =  ( n68 ) == ( bv_8_128_n325 )  ;
assign bv_8_129_n327 = 8'h81 ;
assign n328 =  ( n68 ) == ( bv_8_129_n327 )  ;
assign bv_8_130_n329 = 8'h82 ;
assign n330 =  ( n68 ) == ( bv_8_130_n329 )  ;
assign bv_8_131_n331 = 8'h83 ;
assign n332 =  ( n68 ) == ( bv_8_131_n331 )  ;
assign bv_8_132_n333 = 8'h84 ;
assign n334 =  ( n68 ) == ( bv_8_132_n333 )  ;
assign bv_8_133_n335 = 8'h85 ;
assign n336 =  ( n68 ) == ( bv_8_133_n335 )  ;
assign bv_8_134_n337 = 8'h86 ;
assign n338 =  ( n68 ) == ( bv_8_134_n337 )  ;
assign bv_8_135_n339 = 8'h87 ;
assign n340 =  ( n68 ) == ( bv_8_135_n339 )  ;
assign bv_8_136_n341 = 8'h88 ;
assign n342 =  ( n68 ) == ( bv_8_136_n341 )  ;
assign bv_8_137_n343 = 8'h89 ;
assign n344 =  ( n68 ) == ( bv_8_137_n343 )  ;
assign bv_8_138_n345 = 8'h8a ;
assign n346 =  ( n68 ) == ( bv_8_138_n345 )  ;
assign bv_8_139_n347 = 8'h8b ;
assign n348 =  ( n68 ) == ( bv_8_139_n347 )  ;
assign bv_8_140_n349 = 8'h8c ;
assign n350 =  ( n68 ) == ( bv_8_140_n349 )  ;
assign bv_8_141_n351 = 8'h8d ;
assign n352 =  ( n68 ) == ( bv_8_141_n351 )  ;
assign bv_8_142_n353 = 8'h8e ;
assign n354 =  ( n68 ) == ( bv_8_142_n353 )  ;
assign bv_8_143_n355 = 8'h8f ;
assign n356 =  ( n68 ) == ( bv_8_143_n355 )  ;
assign bv_8_144_n357 = 8'h90 ;
assign n358 =  ( n68 ) == ( bv_8_144_n357 )  ;
assign bv_8_145_n359 = 8'h91 ;
assign n360 =  ( n68 ) == ( bv_8_145_n359 )  ;
assign bv_8_146_n361 = 8'h92 ;
assign n362 =  ( n68 ) == ( bv_8_146_n361 )  ;
assign bv_8_147_n363 = 8'h93 ;
assign n364 =  ( n68 ) == ( bv_8_147_n363 )  ;
assign bv_8_148_n365 = 8'h94 ;
assign n366 =  ( n68 ) == ( bv_8_148_n365 )  ;
assign bv_8_149_n367 = 8'h95 ;
assign n368 =  ( n68 ) == ( bv_8_149_n367 )  ;
assign bv_8_150_n369 = 8'h96 ;
assign n370 =  ( n68 ) == ( bv_8_150_n369 )  ;
assign bv_8_151_n371 = 8'h97 ;
assign n372 =  ( n68 ) == ( bv_8_151_n371 )  ;
assign bv_8_152_n373 = 8'h98 ;
assign n374 =  ( n68 ) == ( bv_8_152_n373 )  ;
assign bv_8_153_n375 = 8'h99 ;
assign n376 =  ( n68 ) == ( bv_8_153_n375 )  ;
assign bv_8_154_n377 = 8'h9a ;
assign n378 =  ( n68 ) == ( bv_8_154_n377 )  ;
assign bv_8_155_n379 = 8'h9b ;
assign n380 =  ( n68 ) == ( bv_8_155_n379 )  ;
assign bv_8_156_n381 = 8'h9c ;
assign n382 =  ( n68 ) == ( bv_8_156_n381 )  ;
assign bv_8_157_n383 = 8'h9d ;
assign n384 =  ( n68 ) == ( bv_8_157_n383 )  ;
assign bv_8_158_n385 = 8'h9e ;
assign n386 =  ( n68 ) == ( bv_8_158_n385 )  ;
assign bv_8_159_n387 = 8'h9f ;
assign n388 =  ( n68 ) == ( bv_8_159_n387 )  ;
assign bv_8_160_n389 = 8'ha0 ;
assign n390 =  ( n68 ) == ( bv_8_160_n389 )  ;
assign bv_8_161_n391 = 8'ha1 ;
assign n392 =  ( n68 ) == ( bv_8_161_n391 )  ;
assign bv_8_162_n393 = 8'ha2 ;
assign n394 =  ( n68 ) == ( bv_8_162_n393 )  ;
assign bv_8_163_n395 = 8'ha3 ;
assign n396 =  ( n68 ) == ( bv_8_163_n395 )  ;
assign bv_8_164_n397 = 8'ha4 ;
assign n398 =  ( n68 ) == ( bv_8_164_n397 )  ;
assign bv_8_165_n399 = 8'ha5 ;
assign n400 =  ( n68 ) == ( bv_8_165_n399 )  ;
assign bv_8_166_n401 = 8'ha6 ;
assign n402 =  ( n68 ) == ( bv_8_166_n401 )  ;
assign bv_8_167_n403 = 8'ha7 ;
assign n404 =  ( n68 ) == ( bv_8_167_n403 )  ;
assign bv_8_168_n405 = 8'ha8 ;
assign n406 =  ( n68 ) == ( bv_8_168_n405 )  ;
assign bv_8_169_n407 = 8'ha9 ;
assign n408 =  ( n68 ) == ( bv_8_169_n407 )  ;
assign bv_8_170_n409 = 8'haa ;
assign n410 =  ( n68 ) == ( bv_8_170_n409 )  ;
assign bv_8_171_n411 = 8'hab ;
assign n412 =  ( n68 ) == ( bv_8_171_n411 )  ;
assign bv_8_172_n413 = 8'hac ;
assign n414 =  ( n68 ) == ( bv_8_172_n413 )  ;
assign bv_8_173_n415 = 8'had ;
assign n416 =  ( n68 ) == ( bv_8_173_n415 )  ;
assign bv_8_174_n417 = 8'hae ;
assign n418 =  ( n68 ) == ( bv_8_174_n417 )  ;
assign bv_8_175_n419 = 8'haf ;
assign n420 =  ( n68 ) == ( bv_8_175_n419 )  ;
assign bv_8_176_n421 = 8'hb0 ;
assign n422 =  ( n68 ) == ( bv_8_176_n421 )  ;
assign bv_8_177_n423 = 8'hb1 ;
assign n424 =  ( n68 ) == ( bv_8_177_n423 )  ;
assign bv_8_178_n425 = 8'hb2 ;
assign n426 =  ( n68 ) == ( bv_8_178_n425 )  ;
assign bv_8_179_n427 = 8'hb3 ;
assign n428 =  ( n68 ) == ( bv_8_179_n427 )  ;
assign bv_8_180_n429 = 8'hb4 ;
assign n430 =  ( n68 ) == ( bv_8_180_n429 )  ;
assign bv_8_181_n431 = 8'hb5 ;
assign n432 =  ( n68 ) == ( bv_8_181_n431 )  ;
assign bv_8_182_n433 = 8'hb6 ;
assign n434 =  ( n68 ) == ( bv_8_182_n433 )  ;
assign bv_8_183_n435 = 8'hb7 ;
assign n436 =  ( n68 ) == ( bv_8_183_n435 )  ;
assign bv_8_184_n437 = 8'hb8 ;
assign n438 =  ( n68 ) == ( bv_8_184_n437 )  ;
assign bv_8_185_n439 = 8'hb9 ;
assign n440 =  ( n68 ) == ( bv_8_185_n439 )  ;
assign bv_8_186_n441 = 8'hba ;
assign n442 =  ( n68 ) == ( bv_8_186_n441 )  ;
assign bv_8_187_n443 = 8'hbb ;
assign n444 =  ( n68 ) == ( bv_8_187_n443 )  ;
assign bv_8_188_n445 = 8'hbc ;
assign n446 =  ( n68 ) == ( bv_8_188_n445 )  ;
assign bv_8_189_n447 = 8'hbd ;
assign n448 =  ( n68 ) == ( bv_8_189_n447 )  ;
assign bv_8_190_n449 = 8'hbe ;
assign n450 =  ( n68 ) == ( bv_8_190_n449 )  ;
assign bv_8_191_n451 = 8'hbf ;
assign n452 =  ( n68 ) == ( bv_8_191_n451 )  ;
assign bv_8_192_n453 = 8'hc0 ;
assign n454 =  ( n68 ) == ( bv_8_192_n453 )  ;
assign bv_8_193_n455 = 8'hc1 ;
assign n456 =  ( n68 ) == ( bv_8_193_n455 )  ;
assign bv_8_194_n457 = 8'hc2 ;
assign n458 =  ( n68 ) == ( bv_8_194_n457 )  ;
assign bv_8_195_n459 = 8'hc3 ;
assign n460 =  ( n68 ) == ( bv_8_195_n459 )  ;
assign bv_8_196_n461 = 8'hc4 ;
assign n462 =  ( n68 ) == ( bv_8_196_n461 )  ;
assign bv_8_197_n463 = 8'hc5 ;
assign n464 =  ( n68 ) == ( bv_8_197_n463 )  ;
assign bv_8_198_n465 = 8'hc6 ;
assign n466 =  ( n68 ) == ( bv_8_198_n465 )  ;
assign bv_8_199_n467 = 8'hc7 ;
assign n468 =  ( n68 ) == ( bv_8_199_n467 )  ;
assign bv_8_200_n469 = 8'hc8 ;
assign n470 =  ( n68 ) == ( bv_8_200_n469 )  ;
assign bv_8_201_n471 = 8'hc9 ;
assign n472 =  ( n68 ) == ( bv_8_201_n471 )  ;
assign bv_8_202_n473 = 8'hca ;
assign n474 =  ( n68 ) == ( bv_8_202_n473 )  ;
assign bv_8_203_n475 = 8'hcb ;
assign n476 =  ( n68 ) == ( bv_8_203_n475 )  ;
assign bv_8_204_n477 = 8'hcc ;
assign n478 =  ( n68 ) == ( bv_8_204_n477 )  ;
assign bv_8_205_n479 = 8'hcd ;
assign n480 =  ( n68 ) == ( bv_8_205_n479 )  ;
assign bv_8_206_n481 = 8'hce ;
assign n482 =  ( n68 ) == ( bv_8_206_n481 )  ;
assign bv_8_207_n483 = 8'hcf ;
assign n484 =  ( n68 ) == ( bv_8_207_n483 )  ;
assign bv_8_208_n485 = 8'hd0 ;
assign n486 =  ( n68 ) == ( bv_8_208_n485 )  ;
assign bv_8_209_n487 = 8'hd1 ;
assign n488 =  ( n68 ) == ( bv_8_209_n487 )  ;
assign bv_8_210_n489 = 8'hd2 ;
assign n490 =  ( n68 ) == ( bv_8_210_n489 )  ;
assign bv_8_211_n491 = 8'hd3 ;
assign n492 =  ( n68 ) == ( bv_8_211_n491 )  ;
assign bv_8_212_n493 = 8'hd4 ;
assign n494 =  ( n68 ) == ( bv_8_212_n493 )  ;
assign bv_8_213_n495 = 8'hd5 ;
assign n496 =  ( n68 ) == ( bv_8_213_n495 )  ;
assign bv_8_214_n497 = 8'hd6 ;
assign n498 =  ( n68 ) == ( bv_8_214_n497 )  ;
assign bv_8_215_n499 = 8'hd7 ;
assign n500 =  ( n68 ) == ( bv_8_215_n499 )  ;
assign bv_8_216_n501 = 8'hd8 ;
assign n502 =  ( n68 ) == ( bv_8_216_n501 )  ;
assign bv_8_217_n503 = 8'hd9 ;
assign n504 =  ( n68 ) == ( bv_8_217_n503 )  ;
assign bv_8_218_n505 = 8'hda ;
assign n506 =  ( n68 ) == ( bv_8_218_n505 )  ;
assign bv_8_219_n507 = 8'hdb ;
assign n508 =  ( n68 ) == ( bv_8_219_n507 )  ;
assign bv_8_220_n509 = 8'hdc ;
assign n510 =  ( n68 ) == ( bv_8_220_n509 )  ;
assign bv_8_221_n511 = 8'hdd ;
assign n512 =  ( n68 ) == ( bv_8_221_n511 )  ;
assign bv_8_222_n513 = 8'hde ;
assign n514 =  ( n68 ) == ( bv_8_222_n513 )  ;
assign bv_8_223_n515 = 8'hdf ;
assign n516 =  ( n68 ) == ( bv_8_223_n515 )  ;
assign bv_8_224_n517 = 8'he0 ;
assign n518 =  ( n68 ) == ( bv_8_224_n517 )  ;
assign bv_8_225_n519 = 8'he1 ;
assign n520 =  ( n68 ) == ( bv_8_225_n519 )  ;
assign bv_8_226_n521 = 8'he2 ;
assign n522 =  ( n68 ) == ( bv_8_226_n521 )  ;
assign bv_8_227_n523 = 8'he3 ;
assign n524 =  ( n68 ) == ( bv_8_227_n523 )  ;
assign bv_8_228_n525 = 8'he4 ;
assign n526 =  ( n68 ) == ( bv_8_228_n525 )  ;
assign bv_8_229_n527 = 8'he5 ;
assign n528 =  ( n68 ) == ( bv_8_229_n527 )  ;
assign bv_8_230_n529 = 8'he6 ;
assign n530 =  ( n68 ) == ( bv_8_230_n529 )  ;
assign bv_8_231_n531 = 8'he7 ;
assign n532 =  ( n68 ) == ( bv_8_231_n531 )  ;
assign bv_8_232_n533 = 8'he8 ;
assign n534 =  ( n68 ) == ( bv_8_232_n533 )  ;
assign bv_8_233_n535 = 8'he9 ;
assign n536 =  ( n68 ) == ( bv_8_233_n535 )  ;
assign bv_8_234_n537 = 8'hea ;
assign n538 =  ( n68 ) == ( bv_8_234_n537 )  ;
assign bv_8_235_n539 = 8'heb ;
assign n540 =  ( n68 ) == ( bv_8_235_n539 )  ;
assign bv_8_236_n541 = 8'hec ;
assign n542 =  ( n68 ) == ( bv_8_236_n541 )  ;
assign bv_8_237_n543 = 8'hed ;
assign n544 =  ( n68 ) == ( bv_8_237_n543 )  ;
assign bv_8_238_n545 = 8'hee ;
assign n546 =  ( n68 ) == ( bv_8_238_n545 )  ;
assign bv_8_239_n547 = 8'hef ;
assign n548 =  ( n68 ) == ( bv_8_239_n547 )  ;
assign bv_8_240_n549 = 8'hf0 ;
assign n550 =  ( n68 ) == ( bv_8_240_n549 )  ;
assign bv_8_241_n551 = 8'hf1 ;
assign n552 =  ( n68 ) == ( bv_8_241_n551 )  ;
assign bv_8_242_n553 = 8'hf2 ;
assign n554 =  ( n68 ) == ( bv_8_242_n553 )  ;
assign bv_8_243_n555 = 8'hf3 ;
assign n556 =  ( n68 ) == ( bv_8_243_n555 )  ;
assign bv_8_244_n557 = 8'hf4 ;
assign n558 =  ( n68 ) == ( bv_8_244_n557 )  ;
assign bv_8_245_n559 = 8'hf5 ;
assign n560 =  ( n68 ) == ( bv_8_245_n559 )  ;
assign bv_8_246_n561 = 8'hf6 ;
assign n562 =  ( n68 ) == ( bv_8_246_n561 )  ;
assign bv_8_247_n563 = 8'hf7 ;
assign n564 =  ( n68 ) == ( bv_8_247_n563 )  ;
assign bv_8_248_n565 = 8'hf8 ;
assign n566 =  ( n68 ) == ( bv_8_248_n565 )  ;
assign bv_8_249_n567 = 8'hf9 ;
assign n568 =  ( n68 ) == ( bv_8_249_n567 )  ;
assign bv_8_250_n569 = 8'hfa ;
assign n570 =  ( n68 ) == ( bv_8_250_n569 )  ;
assign bv_8_251_n571 = 8'hfb ;
assign n572 =  ( n68 ) == ( bv_8_251_n571 )  ;
assign bv_8_252_n573 = 8'hfc ;
assign n574 =  ( n68 ) == ( bv_8_252_n573 )  ;
assign bv_8_253_n575 = 8'hfd ;
assign n576 =  ( n68 ) == ( bv_8_253_n575 )  ;
assign bv_8_254_n577 = 8'hfe ;
assign n578 =  ( n68 ) == ( bv_8_254_n577 )  ;
assign n579 =  ( n578 ) ? ( iram_254 ) : ( iram_255 ) ;
assign n580 =  ( n576 ) ? ( iram_253 ) : ( n579 ) ;
assign n581 =  ( n574 ) ? ( iram_252 ) : ( n580 ) ;
assign n582 =  ( n572 ) ? ( iram_251 ) : ( n581 ) ;
assign n583 =  ( n570 ) ? ( iram_250 ) : ( n582 ) ;
assign n584 =  ( n568 ) ? ( iram_249 ) : ( n583 ) ;
assign n585 =  ( n566 ) ? ( iram_248 ) : ( n584 ) ;
assign n586 =  ( n564 ) ? ( iram_247 ) : ( n585 ) ;
assign n587 =  ( n562 ) ? ( iram_246 ) : ( n586 ) ;
assign n588 =  ( n560 ) ? ( iram_245 ) : ( n587 ) ;
assign n589 =  ( n558 ) ? ( iram_244 ) : ( n588 ) ;
assign n590 =  ( n556 ) ? ( iram_243 ) : ( n589 ) ;
assign n591 =  ( n554 ) ? ( iram_242 ) : ( n590 ) ;
assign n592 =  ( n552 ) ? ( iram_241 ) : ( n591 ) ;
assign n593 =  ( n550 ) ? ( iram_240 ) : ( n592 ) ;
assign n594 =  ( n548 ) ? ( iram_239 ) : ( n593 ) ;
assign n595 =  ( n546 ) ? ( iram_238 ) : ( n594 ) ;
assign n596 =  ( n544 ) ? ( iram_237 ) : ( n595 ) ;
assign n597 =  ( n542 ) ? ( iram_236 ) : ( n596 ) ;
assign n598 =  ( n540 ) ? ( iram_235 ) : ( n597 ) ;
assign n599 =  ( n538 ) ? ( iram_234 ) : ( n598 ) ;
assign n600 =  ( n536 ) ? ( iram_233 ) : ( n599 ) ;
assign n601 =  ( n534 ) ? ( iram_232 ) : ( n600 ) ;
assign n602 =  ( n532 ) ? ( iram_231 ) : ( n601 ) ;
assign n603 =  ( n530 ) ? ( iram_230 ) : ( n602 ) ;
assign n604 =  ( n528 ) ? ( iram_229 ) : ( n603 ) ;
assign n605 =  ( n526 ) ? ( iram_228 ) : ( n604 ) ;
assign n606 =  ( n524 ) ? ( iram_227 ) : ( n605 ) ;
assign n607 =  ( n522 ) ? ( iram_226 ) : ( n606 ) ;
assign n608 =  ( n520 ) ? ( iram_225 ) : ( n607 ) ;
assign n609 =  ( n518 ) ? ( iram_224 ) : ( n608 ) ;
assign n610 =  ( n516 ) ? ( iram_223 ) : ( n609 ) ;
assign n611 =  ( n514 ) ? ( iram_222 ) : ( n610 ) ;
assign n612 =  ( n512 ) ? ( iram_221 ) : ( n611 ) ;
assign n613 =  ( n510 ) ? ( iram_220 ) : ( n612 ) ;
assign n614 =  ( n508 ) ? ( iram_219 ) : ( n613 ) ;
assign n615 =  ( n506 ) ? ( iram_218 ) : ( n614 ) ;
assign n616 =  ( n504 ) ? ( iram_217 ) : ( n615 ) ;
assign n617 =  ( n502 ) ? ( iram_216 ) : ( n616 ) ;
assign n618 =  ( n500 ) ? ( iram_215 ) : ( n617 ) ;
assign n619 =  ( n498 ) ? ( iram_214 ) : ( n618 ) ;
assign n620 =  ( n496 ) ? ( iram_213 ) : ( n619 ) ;
assign n621 =  ( n494 ) ? ( iram_212 ) : ( n620 ) ;
assign n622 =  ( n492 ) ? ( iram_211 ) : ( n621 ) ;
assign n623 =  ( n490 ) ? ( iram_210 ) : ( n622 ) ;
assign n624 =  ( n488 ) ? ( iram_209 ) : ( n623 ) ;
assign n625 =  ( n486 ) ? ( iram_208 ) : ( n624 ) ;
assign n626 =  ( n484 ) ? ( iram_207 ) : ( n625 ) ;
assign n627 =  ( n482 ) ? ( iram_206 ) : ( n626 ) ;
assign n628 =  ( n480 ) ? ( iram_205 ) : ( n627 ) ;
assign n629 =  ( n478 ) ? ( iram_204 ) : ( n628 ) ;
assign n630 =  ( n476 ) ? ( iram_203 ) : ( n629 ) ;
assign n631 =  ( n474 ) ? ( iram_202 ) : ( n630 ) ;
assign n632 =  ( n472 ) ? ( iram_201 ) : ( n631 ) ;
assign n633 =  ( n470 ) ? ( iram_200 ) : ( n632 ) ;
assign n634 =  ( n468 ) ? ( iram_199 ) : ( n633 ) ;
assign n635 =  ( n466 ) ? ( iram_198 ) : ( n634 ) ;
assign n636 =  ( n464 ) ? ( iram_197 ) : ( n635 ) ;
assign n637 =  ( n462 ) ? ( iram_196 ) : ( n636 ) ;
assign n638 =  ( n460 ) ? ( iram_195 ) : ( n637 ) ;
assign n639 =  ( n458 ) ? ( iram_194 ) : ( n638 ) ;
assign n640 =  ( n456 ) ? ( iram_193 ) : ( n639 ) ;
assign n641 =  ( n454 ) ? ( iram_192 ) : ( n640 ) ;
assign n642 =  ( n452 ) ? ( iram_191 ) : ( n641 ) ;
assign n643 =  ( n450 ) ? ( iram_190 ) : ( n642 ) ;
assign n644 =  ( n448 ) ? ( iram_189 ) : ( n643 ) ;
assign n645 =  ( n446 ) ? ( iram_188 ) : ( n644 ) ;
assign n646 =  ( n444 ) ? ( iram_187 ) : ( n645 ) ;
assign n647 =  ( n442 ) ? ( iram_186 ) : ( n646 ) ;
assign n648 =  ( n440 ) ? ( iram_185 ) : ( n647 ) ;
assign n649 =  ( n438 ) ? ( iram_184 ) : ( n648 ) ;
assign n650 =  ( n436 ) ? ( iram_183 ) : ( n649 ) ;
assign n651 =  ( n434 ) ? ( iram_182 ) : ( n650 ) ;
assign n652 =  ( n432 ) ? ( iram_181 ) : ( n651 ) ;
assign n653 =  ( n430 ) ? ( iram_180 ) : ( n652 ) ;
assign n654 =  ( n428 ) ? ( iram_179 ) : ( n653 ) ;
assign n655 =  ( n426 ) ? ( iram_178 ) : ( n654 ) ;
assign n656 =  ( n424 ) ? ( iram_177 ) : ( n655 ) ;
assign n657 =  ( n422 ) ? ( iram_176 ) : ( n656 ) ;
assign n658 =  ( n420 ) ? ( iram_175 ) : ( n657 ) ;
assign n659 =  ( n418 ) ? ( iram_174 ) : ( n658 ) ;
assign n660 =  ( n416 ) ? ( iram_173 ) : ( n659 ) ;
assign n661 =  ( n414 ) ? ( iram_172 ) : ( n660 ) ;
assign n662 =  ( n412 ) ? ( iram_171 ) : ( n661 ) ;
assign n663 =  ( n410 ) ? ( iram_170 ) : ( n662 ) ;
assign n664 =  ( n408 ) ? ( iram_169 ) : ( n663 ) ;
assign n665 =  ( n406 ) ? ( iram_168 ) : ( n664 ) ;
assign n666 =  ( n404 ) ? ( iram_167 ) : ( n665 ) ;
assign n667 =  ( n402 ) ? ( iram_166 ) : ( n666 ) ;
assign n668 =  ( n400 ) ? ( iram_165 ) : ( n667 ) ;
assign n669 =  ( n398 ) ? ( iram_164 ) : ( n668 ) ;
assign n670 =  ( n396 ) ? ( iram_163 ) : ( n669 ) ;
assign n671 =  ( n394 ) ? ( iram_162 ) : ( n670 ) ;
assign n672 =  ( n392 ) ? ( iram_161 ) : ( n671 ) ;
assign n673 =  ( n390 ) ? ( iram_160 ) : ( n672 ) ;
assign n674 =  ( n388 ) ? ( iram_159 ) : ( n673 ) ;
assign n675 =  ( n386 ) ? ( iram_158 ) : ( n674 ) ;
assign n676 =  ( n384 ) ? ( iram_157 ) : ( n675 ) ;
assign n677 =  ( n382 ) ? ( iram_156 ) : ( n676 ) ;
assign n678 =  ( n380 ) ? ( iram_155 ) : ( n677 ) ;
assign n679 =  ( n378 ) ? ( iram_154 ) : ( n678 ) ;
assign n680 =  ( n376 ) ? ( iram_153 ) : ( n679 ) ;
assign n681 =  ( n374 ) ? ( iram_152 ) : ( n680 ) ;
assign n682 =  ( n372 ) ? ( iram_151 ) : ( n681 ) ;
assign n683 =  ( n370 ) ? ( iram_150 ) : ( n682 ) ;
assign n684 =  ( n368 ) ? ( iram_149 ) : ( n683 ) ;
assign n685 =  ( n366 ) ? ( iram_148 ) : ( n684 ) ;
assign n686 =  ( n364 ) ? ( iram_147 ) : ( n685 ) ;
assign n687 =  ( n362 ) ? ( iram_146 ) : ( n686 ) ;
assign n688 =  ( n360 ) ? ( iram_145 ) : ( n687 ) ;
assign n689 =  ( n358 ) ? ( iram_144 ) : ( n688 ) ;
assign n690 =  ( n356 ) ? ( iram_143 ) : ( n689 ) ;
assign n691 =  ( n354 ) ? ( iram_142 ) : ( n690 ) ;
assign n692 =  ( n352 ) ? ( iram_141 ) : ( n691 ) ;
assign n693 =  ( n350 ) ? ( iram_140 ) : ( n692 ) ;
assign n694 =  ( n348 ) ? ( iram_139 ) : ( n693 ) ;
assign n695 =  ( n346 ) ? ( iram_138 ) : ( n694 ) ;
assign n696 =  ( n344 ) ? ( iram_137 ) : ( n695 ) ;
assign n697 =  ( n342 ) ? ( iram_136 ) : ( n696 ) ;
assign n698 =  ( n340 ) ? ( iram_135 ) : ( n697 ) ;
assign n699 =  ( n338 ) ? ( iram_134 ) : ( n698 ) ;
assign n700 =  ( n336 ) ? ( iram_133 ) : ( n699 ) ;
assign n701 =  ( n334 ) ? ( iram_132 ) : ( n700 ) ;
assign n702 =  ( n332 ) ? ( iram_131 ) : ( n701 ) ;
assign n703 =  ( n330 ) ? ( iram_130 ) : ( n702 ) ;
assign n704 =  ( n328 ) ? ( iram_129 ) : ( n703 ) ;
assign n705 =  ( n326 ) ? ( iram_128 ) : ( n704 ) ;
assign n706 =  ( n324 ) ? ( iram_127 ) : ( n705 ) ;
assign n707 =  ( n322 ) ? ( iram_126 ) : ( n706 ) ;
assign n708 =  ( n320 ) ? ( iram_125 ) : ( n707 ) ;
assign n709 =  ( n318 ) ? ( iram_124 ) : ( n708 ) ;
assign n710 =  ( n316 ) ? ( iram_123 ) : ( n709 ) ;
assign n711 =  ( n314 ) ? ( iram_122 ) : ( n710 ) ;
assign n712 =  ( n312 ) ? ( iram_121 ) : ( n711 ) ;
assign n713 =  ( n310 ) ? ( iram_120 ) : ( n712 ) ;
assign n714 =  ( n308 ) ? ( iram_119 ) : ( n713 ) ;
assign n715 =  ( n306 ) ? ( iram_118 ) : ( n714 ) ;
assign n716 =  ( n304 ) ? ( iram_117 ) : ( n715 ) ;
assign n717 =  ( n302 ) ? ( iram_116 ) : ( n716 ) ;
assign n718 =  ( n300 ) ? ( iram_115 ) : ( n717 ) ;
assign n719 =  ( n298 ) ? ( iram_114 ) : ( n718 ) ;
assign n720 =  ( n296 ) ? ( iram_113 ) : ( n719 ) ;
assign n721 =  ( n294 ) ? ( iram_112 ) : ( n720 ) ;
assign n722 =  ( n292 ) ? ( iram_111 ) : ( n721 ) ;
assign n723 =  ( n290 ) ? ( iram_110 ) : ( n722 ) ;
assign n724 =  ( n288 ) ? ( iram_109 ) : ( n723 ) ;
assign n725 =  ( n286 ) ? ( iram_108 ) : ( n724 ) ;
assign n726 =  ( n284 ) ? ( iram_107 ) : ( n725 ) ;
assign n727 =  ( n282 ) ? ( iram_106 ) : ( n726 ) ;
assign n728 =  ( n280 ) ? ( iram_105 ) : ( n727 ) ;
assign n729 =  ( n278 ) ? ( iram_104 ) : ( n728 ) ;
assign n730 =  ( n276 ) ? ( iram_103 ) : ( n729 ) ;
assign n731 =  ( n274 ) ? ( iram_102 ) : ( n730 ) ;
assign n732 =  ( n272 ) ? ( iram_101 ) : ( n731 ) ;
assign n733 =  ( n270 ) ? ( iram_100 ) : ( n732 ) ;
assign n734 =  ( n268 ) ? ( iram_99 ) : ( n733 ) ;
assign n735 =  ( n266 ) ? ( iram_98 ) : ( n734 ) ;
assign n736 =  ( n264 ) ? ( iram_97 ) : ( n735 ) ;
assign n737 =  ( n262 ) ? ( iram_96 ) : ( n736 ) ;
assign n738 =  ( n260 ) ? ( iram_95 ) : ( n737 ) ;
assign n739 =  ( n258 ) ? ( iram_94 ) : ( n738 ) ;
assign n740 =  ( n256 ) ? ( iram_93 ) : ( n739 ) ;
assign n741 =  ( n254 ) ? ( iram_92 ) : ( n740 ) ;
assign n742 =  ( n252 ) ? ( iram_91 ) : ( n741 ) ;
assign n743 =  ( n250 ) ? ( iram_90 ) : ( n742 ) ;
assign n744 =  ( n248 ) ? ( iram_89 ) : ( n743 ) ;
assign n745 =  ( n246 ) ? ( iram_88 ) : ( n744 ) ;
assign n746 =  ( n244 ) ? ( iram_87 ) : ( n745 ) ;
assign n747 =  ( n242 ) ? ( iram_86 ) : ( n746 ) ;
assign n748 =  ( n240 ) ? ( iram_85 ) : ( n747 ) ;
assign n749 =  ( n238 ) ? ( iram_84 ) : ( n748 ) ;
assign n750 =  ( n236 ) ? ( iram_83 ) : ( n749 ) ;
assign n751 =  ( n234 ) ? ( iram_82 ) : ( n750 ) ;
assign n752 =  ( n232 ) ? ( iram_81 ) : ( n751 ) ;
assign n753 =  ( n230 ) ? ( iram_80 ) : ( n752 ) ;
assign n754 =  ( n228 ) ? ( iram_79 ) : ( n753 ) ;
assign n755 =  ( n226 ) ? ( iram_78 ) : ( n754 ) ;
assign n756 =  ( n224 ) ? ( iram_77 ) : ( n755 ) ;
assign n757 =  ( n222 ) ? ( iram_76 ) : ( n756 ) ;
assign n758 =  ( n220 ) ? ( iram_75 ) : ( n757 ) ;
assign n759 =  ( n218 ) ? ( iram_74 ) : ( n758 ) ;
assign n760 =  ( n216 ) ? ( iram_73 ) : ( n759 ) ;
assign n761 =  ( n214 ) ? ( iram_72 ) : ( n760 ) ;
assign n762 =  ( n212 ) ? ( iram_71 ) : ( n761 ) ;
assign n763 =  ( n210 ) ? ( iram_70 ) : ( n762 ) ;
assign n764 =  ( n208 ) ? ( iram_69 ) : ( n763 ) ;
assign n765 =  ( n206 ) ? ( iram_68 ) : ( n764 ) ;
assign n766 =  ( n204 ) ? ( iram_67 ) : ( n765 ) ;
assign n767 =  ( n202 ) ? ( iram_66 ) : ( n766 ) ;
assign n768 =  ( n200 ) ? ( iram_65 ) : ( n767 ) ;
assign n769 =  ( n198 ) ? ( iram_64 ) : ( n768 ) ;
assign n770 =  ( n196 ) ? ( iram_63 ) : ( n769 ) ;
assign n771 =  ( n194 ) ? ( iram_62 ) : ( n770 ) ;
assign n772 =  ( n192 ) ? ( iram_61 ) : ( n771 ) ;
assign n773 =  ( n190 ) ? ( iram_60 ) : ( n772 ) ;
assign n774 =  ( n188 ) ? ( iram_59 ) : ( n773 ) ;
assign n775 =  ( n186 ) ? ( iram_58 ) : ( n774 ) ;
assign n776 =  ( n184 ) ? ( iram_57 ) : ( n775 ) ;
assign n777 =  ( n182 ) ? ( iram_56 ) : ( n776 ) ;
assign n778 =  ( n180 ) ? ( iram_55 ) : ( n777 ) ;
assign n779 =  ( n178 ) ? ( iram_54 ) : ( n778 ) ;
assign n780 =  ( n176 ) ? ( iram_53 ) : ( n779 ) ;
assign n781 =  ( n174 ) ? ( iram_52 ) : ( n780 ) ;
assign n782 =  ( n172 ) ? ( iram_51 ) : ( n781 ) ;
assign n783 =  ( n170 ) ? ( iram_50 ) : ( n782 ) ;
assign n784 =  ( n168 ) ? ( iram_49 ) : ( n783 ) ;
assign n785 =  ( n166 ) ? ( iram_48 ) : ( n784 ) ;
assign n786 =  ( n164 ) ? ( iram_47 ) : ( n785 ) ;
assign n787 =  ( n162 ) ? ( iram_46 ) : ( n786 ) ;
assign n788 =  ( n160 ) ? ( iram_45 ) : ( n787 ) ;
assign n789 =  ( n158 ) ? ( iram_44 ) : ( n788 ) ;
assign n790 =  ( n156 ) ? ( iram_43 ) : ( n789 ) ;
assign n791 =  ( n154 ) ? ( iram_42 ) : ( n790 ) ;
assign n792 =  ( n152 ) ? ( iram_41 ) : ( n791 ) ;
assign n793 =  ( n150 ) ? ( iram_40 ) : ( n792 ) ;
assign n794 =  ( n148 ) ? ( iram_39 ) : ( n793 ) ;
assign n795 =  ( n146 ) ? ( iram_38 ) : ( n794 ) ;
assign n796 =  ( n144 ) ? ( iram_37 ) : ( n795 ) ;
assign n797 =  ( n142 ) ? ( iram_36 ) : ( n796 ) ;
assign n798 =  ( n140 ) ? ( iram_35 ) : ( n797 ) ;
assign n799 =  ( n138 ) ? ( iram_34 ) : ( n798 ) ;
assign n800 =  ( n136 ) ? ( iram_33 ) : ( n799 ) ;
assign n801 =  ( n134 ) ? ( iram_32 ) : ( n800 ) ;
assign n802 =  ( n132 ) ? ( iram_31 ) : ( n801 ) ;
assign n803 =  ( n130 ) ? ( iram_30 ) : ( n802 ) ;
assign n804 =  ( n128 ) ? ( iram_29 ) : ( n803 ) ;
assign n805 =  ( n126 ) ? ( iram_28 ) : ( n804 ) ;
assign n806 =  ( n124 ) ? ( iram_27 ) : ( n805 ) ;
assign n807 =  ( n122 ) ? ( iram_26 ) : ( n806 ) ;
assign n808 =  ( n120 ) ? ( iram_25 ) : ( n807 ) ;
assign n809 =  ( n118 ) ? ( iram_24 ) : ( n808 ) ;
assign n810 =  ( n116 ) ? ( iram_23 ) : ( n809 ) ;
assign n811 =  ( n114 ) ? ( iram_22 ) : ( n810 ) ;
assign n812 =  ( n112 ) ? ( iram_21 ) : ( n811 ) ;
assign n813 =  ( n110 ) ? ( iram_20 ) : ( n812 ) ;
assign n814 =  ( n108 ) ? ( iram_19 ) : ( n813 ) ;
assign n815 =  ( n106 ) ? ( iram_18 ) : ( n814 ) ;
assign n816 =  ( n104 ) ? ( iram_17 ) : ( n815 ) ;
assign n817 =  ( n102 ) ? ( iram_16 ) : ( n816 ) ;
assign n818 =  ( n100 ) ? ( iram_15 ) : ( n817 ) ;
assign n819 =  ( n98 ) ? ( iram_14 ) : ( n818 ) ;
assign n820 =  ( n96 ) ? ( iram_13 ) : ( n819 ) ;
assign n821 =  ( n94 ) ? ( iram_12 ) : ( n820 ) ;
assign n822 =  ( n92 ) ? ( iram_11 ) : ( n821 ) ;
assign n823 =  ( n90 ) ? ( iram_10 ) : ( n822 ) ;
assign n824 =  ( n88 ) ? ( iram_9 ) : ( n823 ) ;
assign n825 =  ( n86 ) ? ( iram_8 ) : ( n824 ) ;
assign n826 =  ( n84 ) ? ( iram_7 ) : ( n825 ) ;
assign n827 =  ( n82 ) ? ( iram_6 ) : ( n826 ) ;
assign n828 =  ( n80 ) ? ( iram_5 ) : ( n827 ) ;
assign n829 =  ( n78 ) ? ( iram_4 ) : ( n828 ) ;
assign n830 =  ( n76 ) ? ( iram_3 ) : ( n829 ) ;
assign n831 =  ( n74 ) ? ( iram_2 ) : ( n830 ) ;
assign n832 =  ( n72 ) ? ( iram_1 ) : ( n831 ) ;
assign n833 =  ( n70 ) ? ( iram_0 ) : ( n832 ) ;
assign n834 =  ( rd_addr ) == ( bv_8_0_n69 )  ;
assign n835 =  ( rd_addr ) == ( bv_8_1_n71 )  ;
assign n836 =  ( rd_addr ) == ( bv_8_2_n73 )  ;
assign n837 =  ( rd_addr ) == ( bv_8_3_n75 )  ;
assign n838 =  ( rd_addr ) == ( bv_8_4_n77 )  ;
assign n839 =  ( rd_addr ) == ( bv_8_5_n79 )  ;
assign n840 =  ( rd_addr ) == ( bv_8_6_n81 )  ;
assign n841 =  ( rd_addr ) == ( bv_8_7_n83 )  ;
assign n842 =  ( rd_addr ) == ( bv_8_8_n85 )  ;
assign n843 =  ( rd_addr ) == ( bv_8_9_n87 )  ;
assign n844 =  ( rd_addr ) == ( bv_8_10_n89 )  ;
assign n845 =  ( rd_addr ) == ( bv_8_11_n91 )  ;
assign n846 =  ( rd_addr ) == ( bv_8_12_n93 )  ;
assign n847 =  ( rd_addr ) == ( bv_8_13_n95 )  ;
assign n848 =  ( rd_addr ) == ( bv_8_14_n97 )  ;
assign n849 =  ( rd_addr ) == ( bv_8_15_n99 )  ;
assign n850 =  ( rd_addr ) == ( bv_8_16_n101 )  ;
assign n851 =  ( rd_addr ) == ( bv_8_17_n103 )  ;
assign n852 =  ( rd_addr ) == ( bv_8_18_n105 )  ;
assign n853 =  ( rd_addr ) == ( bv_8_19_n107 )  ;
assign n854 =  ( rd_addr ) == ( bv_8_20_n109 )  ;
assign n855 =  ( rd_addr ) == ( bv_8_21_n111 )  ;
assign n856 =  ( rd_addr ) == ( bv_8_22_n113 )  ;
assign n857 =  ( rd_addr ) == ( bv_8_23_n115 )  ;
assign n858 =  ( rd_addr ) == ( bv_8_24_n117 )  ;
assign n859 =  ( rd_addr ) == ( bv_8_25_n119 )  ;
assign n860 =  ( rd_addr ) == ( bv_8_26_n121 )  ;
assign n861 =  ( rd_addr ) == ( bv_8_27_n123 )  ;
assign n862 =  ( rd_addr ) == ( bv_8_28_n125 )  ;
assign n863 =  ( rd_addr ) == ( bv_8_29_n127 )  ;
assign n864 =  ( rd_addr ) == ( bv_8_30_n129 )  ;
assign n865 =  ( rd_addr ) == ( bv_8_31_n131 )  ;
assign n866 =  ( rd_addr ) == ( bv_8_32_n133 )  ;
assign n867 =  ( rd_addr ) == ( bv_8_33_n135 )  ;
assign n868 =  ( rd_addr ) == ( bv_8_34_n137 )  ;
assign n869 =  ( rd_addr ) == ( bv_8_35_n139 )  ;
assign n870 =  ( rd_addr ) == ( bv_8_36_n141 )  ;
assign n871 =  ( rd_addr ) == ( bv_8_37_n143 )  ;
assign n872 =  ( rd_addr ) == ( bv_8_38_n145 )  ;
assign n873 =  ( rd_addr ) == ( bv_8_39_n147 )  ;
assign n874 =  ( rd_addr ) == ( bv_8_40_n149 )  ;
assign n875 =  ( rd_addr ) == ( bv_8_41_n151 )  ;
assign n876 =  ( rd_addr ) == ( bv_8_42_n153 )  ;
assign n877 =  ( rd_addr ) == ( bv_8_43_n155 )  ;
assign n878 =  ( rd_addr ) == ( bv_8_44_n157 )  ;
assign n879 =  ( rd_addr ) == ( bv_8_45_n159 )  ;
assign n880 =  ( rd_addr ) == ( bv_8_46_n161 )  ;
assign n881 =  ( rd_addr ) == ( bv_8_47_n163 )  ;
assign n882 =  ( rd_addr ) == ( bv_8_48_n165 )  ;
assign n883 =  ( rd_addr ) == ( bv_8_49_n167 )  ;
assign n884 =  ( rd_addr ) == ( bv_8_50_n169 )  ;
assign n885 =  ( rd_addr ) == ( bv_8_51_n171 )  ;
assign n886 =  ( rd_addr ) == ( bv_8_52_n173 )  ;
assign n887 =  ( rd_addr ) == ( bv_8_53_n175 )  ;
assign n888 =  ( rd_addr ) == ( bv_8_54_n177 )  ;
assign n889 =  ( rd_addr ) == ( bv_8_55_n179 )  ;
assign n890 =  ( rd_addr ) == ( bv_8_56_n181 )  ;
assign n891 =  ( rd_addr ) == ( bv_8_57_n183 )  ;
assign n892 =  ( rd_addr ) == ( bv_8_58_n185 )  ;
assign n893 =  ( rd_addr ) == ( bv_8_59_n187 )  ;
assign n894 =  ( rd_addr ) == ( bv_8_60_n189 )  ;
assign n895 =  ( rd_addr ) == ( bv_8_61_n191 )  ;
assign n896 =  ( rd_addr ) == ( bv_8_62_n193 )  ;
assign n897 =  ( rd_addr ) == ( bv_8_63_n195 )  ;
assign n898 =  ( rd_addr ) == ( bv_8_64_n197 )  ;
assign n899 =  ( rd_addr ) == ( bv_8_65_n199 )  ;
assign n900 =  ( rd_addr ) == ( bv_8_66_n201 )  ;
assign n901 =  ( rd_addr ) == ( bv_8_67_n203 )  ;
assign n902 =  ( rd_addr ) == ( bv_8_68_n205 )  ;
assign n903 =  ( rd_addr ) == ( bv_8_69_n207 )  ;
assign n904 =  ( rd_addr ) == ( bv_8_70_n209 )  ;
assign n905 =  ( rd_addr ) == ( bv_8_71_n211 )  ;
assign n906 =  ( rd_addr ) == ( bv_8_72_n213 )  ;
assign n907 =  ( rd_addr ) == ( bv_8_73_n215 )  ;
assign n908 =  ( rd_addr ) == ( bv_8_74_n217 )  ;
assign n909 =  ( rd_addr ) == ( bv_8_75_n219 )  ;
assign n910 =  ( rd_addr ) == ( bv_8_76_n221 )  ;
assign n911 =  ( rd_addr ) == ( bv_8_77_n223 )  ;
assign n912 =  ( rd_addr ) == ( bv_8_78_n225 )  ;
assign n913 =  ( rd_addr ) == ( bv_8_79_n227 )  ;
assign n914 =  ( rd_addr ) == ( bv_8_80_n229 )  ;
assign n915 =  ( rd_addr ) == ( bv_8_81_n231 )  ;
assign n916 =  ( rd_addr ) == ( bv_8_82_n233 )  ;
assign n917 =  ( rd_addr ) == ( bv_8_83_n235 )  ;
assign n918 =  ( rd_addr ) == ( bv_8_84_n237 )  ;
assign n919 =  ( rd_addr ) == ( bv_8_85_n239 )  ;
assign n920 =  ( rd_addr ) == ( bv_8_86_n241 )  ;
assign n921 =  ( rd_addr ) == ( bv_8_87_n243 )  ;
assign n922 =  ( rd_addr ) == ( bv_8_88_n245 )  ;
assign n923 =  ( rd_addr ) == ( bv_8_89_n247 )  ;
assign n924 =  ( rd_addr ) == ( bv_8_90_n249 )  ;
assign n925 =  ( rd_addr ) == ( bv_8_91_n251 )  ;
assign n926 =  ( rd_addr ) == ( bv_8_92_n253 )  ;
assign n927 =  ( rd_addr ) == ( bv_8_93_n255 )  ;
assign n928 =  ( rd_addr ) == ( bv_8_94_n257 )  ;
assign n929 =  ( rd_addr ) == ( bv_8_95_n259 )  ;
assign n930 =  ( rd_addr ) == ( bv_8_96_n261 )  ;
assign n931 =  ( rd_addr ) == ( bv_8_97_n263 )  ;
assign n932 =  ( rd_addr ) == ( bv_8_98_n265 )  ;
assign n933 =  ( rd_addr ) == ( bv_8_99_n267 )  ;
assign n934 =  ( rd_addr ) == ( bv_8_100_n269 )  ;
assign n935 =  ( rd_addr ) == ( bv_8_101_n271 )  ;
assign n936 =  ( rd_addr ) == ( bv_8_102_n273 )  ;
assign n937 =  ( rd_addr ) == ( bv_8_103_n275 )  ;
assign n938 =  ( rd_addr ) == ( bv_8_104_n277 )  ;
assign n939 =  ( rd_addr ) == ( bv_8_105_n279 )  ;
assign n940 =  ( rd_addr ) == ( bv_8_106_n281 )  ;
assign n941 =  ( rd_addr ) == ( bv_8_107_n283 )  ;
assign n942 =  ( rd_addr ) == ( bv_8_108_n285 )  ;
assign n943 =  ( rd_addr ) == ( bv_8_109_n287 )  ;
assign n944 =  ( rd_addr ) == ( bv_8_110_n289 )  ;
assign n945 =  ( rd_addr ) == ( bv_8_111_n291 )  ;
assign n946 =  ( rd_addr ) == ( bv_8_112_n293 )  ;
assign n947 =  ( rd_addr ) == ( bv_8_113_n295 )  ;
assign n948 =  ( rd_addr ) == ( bv_8_114_n297 )  ;
assign n949 =  ( rd_addr ) == ( bv_8_115_n299 )  ;
assign n950 =  ( rd_addr ) == ( bv_8_116_n301 )  ;
assign n951 =  ( rd_addr ) == ( bv_8_117_n303 )  ;
assign n952 =  ( rd_addr ) == ( bv_8_118_n305 )  ;
assign n953 =  ( rd_addr ) == ( bv_8_119_n307 )  ;
assign n954 =  ( rd_addr ) == ( bv_8_120_n309 )  ;
assign n955 =  ( rd_addr ) == ( bv_8_121_n311 )  ;
assign n956 =  ( rd_addr ) == ( bv_8_122_n313 )  ;
assign n957 =  ( rd_addr ) == ( bv_8_123_n315 )  ;
assign n958 =  ( rd_addr ) == ( bv_8_124_n317 )  ;
assign n959 =  ( rd_addr ) == ( bv_8_125_n319 )  ;
assign n960 =  ( rd_addr ) == ( bv_8_126_n321 )  ;
assign n961 =  ( rd_addr ) == ( bv_8_127_n323 )  ;
assign n962 =  ( rd_addr ) == ( bv_8_128_n325 )  ;
assign n963 =  ( rd_addr ) == ( bv_8_129_n327 )  ;
assign n964 =  ( rd_addr ) == ( bv_8_130_n329 )  ;
assign n965 =  ( rd_addr ) == ( bv_8_131_n331 )  ;
assign n966 =  ( rd_addr ) == ( bv_8_132_n333 )  ;
assign n967 =  ( rd_addr ) == ( bv_8_133_n335 )  ;
assign n968 =  ( rd_addr ) == ( bv_8_134_n337 )  ;
assign n969 =  ( rd_addr ) == ( bv_8_135_n339 )  ;
assign n970 =  ( rd_addr ) == ( bv_8_136_n341 )  ;
assign n971 =  ( rd_addr ) == ( bv_8_137_n343 )  ;
assign n972 =  ( rd_addr ) == ( bv_8_138_n345 )  ;
assign n973 =  ( rd_addr ) == ( bv_8_139_n347 )  ;
assign n974 =  ( rd_addr ) == ( bv_8_140_n349 )  ;
assign n975 =  ( rd_addr ) == ( bv_8_141_n351 )  ;
assign n976 =  ( rd_addr ) == ( bv_8_142_n353 )  ;
assign n977 =  ( rd_addr ) == ( bv_8_143_n355 )  ;
assign n978 =  ( rd_addr ) == ( bv_8_144_n357 )  ;
assign n979 =  ( rd_addr ) == ( bv_8_145_n359 )  ;
assign n980 =  ( rd_addr ) == ( bv_8_146_n361 )  ;
assign n981 =  ( rd_addr ) == ( bv_8_147_n363 )  ;
assign n982 =  ( rd_addr ) == ( bv_8_148_n365 )  ;
assign n983 =  ( rd_addr ) == ( bv_8_149_n367 )  ;
assign n984 =  ( rd_addr ) == ( bv_8_150_n369 )  ;
assign n985 =  ( rd_addr ) == ( bv_8_151_n371 )  ;
assign n986 =  ( rd_addr ) == ( bv_8_152_n373 )  ;
assign n987 =  ( rd_addr ) == ( bv_8_153_n375 )  ;
assign n988 =  ( rd_addr ) == ( bv_8_154_n377 )  ;
assign n989 =  ( rd_addr ) == ( bv_8_155_n379 )  ;
assign n990 =  ( rd_addr ) == ( bv_8_156_n381 )  ;
assign n991 =  ( rd_addr ) == ( bv_8_157_n383 )  ;
assign n992 =  ( rd_addr ) == ( bv_8_158_n385 )  ;
assign n993 =  ( rd_addr ) == ( bv_8_159_n387 )  ;
assign n994 =  ( rd_addr ) == ( bv_8_160_n389 )  ;
assign n995 =  ( rd_addr ) == ( bv_8_161_n391 )  ;
assign n996 =  ( rd_addr ) == ( bv_8_162_n393 )  ;
assign n997 =  ( rd_addr ) == ( bv_8_163_n395 )  ;
assign n998 =  ( rd_addr ) == ( bv_8_164_n397 )  ;
assign n999 =  ( rd_addr ) == ( bv_8_165_n399 )  ;
assign n1000 =  ( rd_addr ) == ( bv_8_166_n401 )  ;
assign n1001 =  ( rd_addr ) == ( bv_8_167_n403 )  ;
assign n1002 =  ( rd_addr ) == ( bv_8_168_n405 )  ;
assign n1003 =  ( rd_addr ) == ( bv_8_169_n407 )  ;
assign n1004 =  ( rd_addr ) == ( bv_8_170_n409 )  ;
assign n1005 =  ( rd_addr ) == ( bv_8_171_n411 )  ;
assign n1006 =  ( rd_addr ) == ( bv_8_172_n413 )  ;
assign n1007 =  ( rd_addr ) == ( bv_8_173_n415 )  ;
assign n1008 =  ( rd_addr ) == ( bv_8_174_n417 )  ;
assign n1009 =  ( rd_addr ) == ( bv_8_175_n419 )  ;
assign n1010 =  ( rd_addr ) == ( bv_8_176_n421 )  ;
assign n1011 =  ( rd_addr ) == ( bv_8_177_n423 )  ;
assign n1012 =  ( rd_addr ) == ( bv_8_178_n425 )  ;
assign n1013 =  ( rd_addr ) == ( bv_8_179_n427 )  ;
assign n1014 =  ( rd_addr ) == ( bv_8_180_n429 )  ;
assign n1015 =  ( rd_addr ) == ( bv_8_181_n431 )  ;
assign n1016 =  ( rd_addr ) == ( bv_8_182_n433 )  ;
assign n1017 =  ( rd_addr ) == ( bv_8_183_n435 )  ;
assign n1018 =  ( rd_addr ) == ( bv_8_184_n437 )  ;
assign n1019 =  ( rd_addr ) == ( bv_8_185_n439 )  ;
assign n1020 =  ( rd_addr ) == ( bv_8_186_n441 )  ;
assign n1021 =  ( rd_addr ) == ( bv_8_187_n443 )  ;
assign n1022 =  ( rd_addr ) == ( bv_8_188_n445 )  ;
assign n1023 =  ( rd_addr ) == ( bv_8_189_n447 )  ;
assign n1024 =  ( rd_addr ) == ( bv_8_190_n449 )  ;
assign n1025 =  ( rd_addr ) == ( bv_8_191_n451 )  ;
assign n1026 =  ( rd_addr ) == ( bv_8_192_n453 )  ;
assign n1027 =  ( rd_addr ) == ( bv_8_193_n455 )  ;
assign n1028 =  ( rd_addr ) == ( bv_8_194_n457 )  ;
assign n1029 =  ( rd_addr ) == ( bv_8_195_n459 )  ;
assign n1030 =  ( rd_addr ) == ( bv_8_196_n461 )  ;
assign n1031 =  ( rd_addr ) == ( bv_8_197_n463 )  ;
assign n1032 =  ( rd_addr ) == ( bv_8_198_n465 )  ;
assign n1033 =  ( rd_addr ) == ( bv_8_199_n467 )  ;
assign n1034 =  ( rd_addr ) == ( bv_8_200_n469 )  ;
assign n1035 =  ( rd_addr ) == ( bv_8_201_n471 )  ;
assign n1036 =  ( rd_addr ) == ( bv_8_202_n473 )  ;
assign n1037 =  ( rd_addr ) == ( bv_8_203_n475 )  ;
assign n1038 =  ( rd_addr ) == ( bv_8_204_n477 )  ;
assign n1039 =  ( rd_addr ) == ( bv_8_205_n479 )  ;
assign n1040 =  ( rd_addr ) == ( bv_8_206_n481 )  ;
assign n1041 =  ( rd_addr ) == ( bv_8_207_n483 )  ;
assign n1042 =  ( rd_addr ) == ( bv_8_208_n485 )  ;
assign n1043 =  ( rd_addr ) == ( bv_8_209_n487 )  ;
assign n1044 =  ( rd_addr ) == ( bv_8_210_n489 )  ;
assign n1045 =  ( rd_addr ) == ( bv_8_211_n491 )  ;
assign n1046 =  ( rd_addr ) == ( bv_8_212_n493 )  ;
assign n1047 =  ( rd_addr ) == ( bv_8_213_n495 )  ;
assign n1048 =  ( rd_addr ) == ( bv_8_214_n497 )  ;
assign n1049 =  ( rd_addr ) == ( bv_8_215_n499 )  ;
assign n1050 =  ( rd_addr ) == ( bv_8_216_n501 )  ;
assign n1051 =  ( rd_addr ) == ( bv_8_217_n503 )  ;
assign n1052 =  ( rd_addr ) == ( bv_8_218_n505 )  ;
assign n1053 =  ( rd_addr ) == ( bv_8_219_n507 )  ;
assign n1054 =  ( rd_addr ) == ( bv_8_220_n509 )  ;
assign n1055 =  ( rd_addr ) == ( bv_8_221_n511 )  ;
assign n1056 =  ( rd_addr ) == ( bv_8_222_n513 )  ;
assign n1057 =  ( rd_addr ) == ( bv_8_223_n515 )  ;
assign n1058 =  ( rd_addr ) == ( bv_8_224_n517 )  ;
assign n1059 =  ( rd_addr ) == ( bv_8_225_n519 )  ;
assign n1060 =  ( rd_addr ) == ( bv_8_226_n521 )  ;
assign n1061 =  ( rd_addr ) == ( bv_8_227_n523 )  ;
assign n1062 =  ( rd_addr ) == ( bv_8_228_n525 )  ;
assign n1063 =  ( rd_addr ) == ( bv_8_229_n527 )  ;
assign n1064 =  ( rd_addr ) == ( bv_8_230_n529 )  ;
assign n1065 =  ( rd_addr ) == ( bv_8_231_n531 )  ;
assign n1066 =  ( rd_addr ) == ( bv_8_232_n533 )  ;
assign n1067 =  ( rd_addr ) == ( bv_8_233_n535 )  ;
assign n1068 =  ( rd_addr ) == ( bv_8_234_n537 )  ;
assign n1069 =  ( rd_addr ) == ( bv_8_235_n539 )  ;
assign n1070 =  ( rd_addr ) == ( bv_8_236_n541 )  ;
assign n1071 =  ( rd_addr ) == ( bv_8_237_n543 )  ;
assign n1072 =  ( rd_addr ) == ( bv_8_238_n545 )  ;
assign n1073 =  ( rd_addr ) == ( bv_8_239_n547 )  ;
assign n1074 =  ( rd_addr ) == ( bv_8_240_n549 )  ;
assign n1075 =  ( rd_addr ) == ( bv_8_241_n551 )  ;
assign n1076 =  ( rd_addr ) == ( bv_8_242_n553 )  ;
assign n1077 =  ( rd_addr ) == ( bv_8_243_n555 )  ;
assign n1078 =  ( rd_addr ) == ( bv_8_244_n557 )  ;
assign n1079 =  ( rd_addr ) == ( bv_8_245_n559 )  ;
assign n1080 =  ( rd_addr ) == ( bv_8_246_n561 )  ;
assign n1081 =  ( rd_addr ) == ( bv_8_247_n563 )  ;
assign n1082 =  ( rd_addr ) == ( bv_8_248_n565 )  ;
assign n1083 =  ( rd_addr ) == ( bv_8_249_n567 )  ;
assign n1084 =  ( rd_addr ) == ( bv_8_250_n569 )  ;
assign n1085 =  ( rd_addr ) == ( bv_8_251_n571 )  ;
assign n1086 =  ( rd_addr ) == ( bv_8_252_n573 )  ;
assign n1087 =  ( rd_addr ) == ( bv_8_253_n575 )  ;
assign n1088 =  ( rd_addr ) == ( bv_8_254_n577 )  ;
assign n1089 =  ( n1088 ) ? ( iram_254 ) : ( iram_255 ) ;
assign n1090 =  ( n1087 ) ? ( iram_253 ) : ( n1089 ) ;
assign n1091 =  ( n1086 ) ? ( iram_252 ) : ( n1090 ) ;
assign n1092 =  ( n1085 ) ? ( iram_251 ) : ( n1091 ) ;
assign n1093 =  ( n1084 ) ? ( iram_250 ) : ( n1092 ) ;
assign n1094 =  ( n1083 ) ? ( iram_249 ) : ( n1093 ) ;
assign n1095 =  ( n1082 ) ? ( iram_248 ) : ( n1094 ) ;
assign n1096 =  ( n1081 ) ? ( iram_247 ) : ( n1095 ) ;
assign n1097 =  ( n1080 ) ? ( iram_246 ) : ( n1096 ) ;
assign n1098 =  ( n1079 ) ? ( iram_245 ) : ( n1097 ) ;
assign n1099 =  ( n1078 ) ? ( iram_244 ) : ( n1098 ) ;
assign n1100 =  ( n1077 ) ? ( iram_243 ) : ( n1099 ) ;
assign n1101 =  ( n1076 ) ? ( iram_242 ) : ( n1100 ) ;
assign n1102 =  ( n1075 ) ? ( iram_241 ) : ( n1101 ) ;
assign n1103 =  ( n1074 ) ? ( iram_240 ) : ( n1102 ) ;
assign n1104 =  ( n1073 ) ? ( iram_239 ) : ( n1103 ) ;
assign n1105 =  ( n1072 ) ? ( iram_238 ) : ( n1104 ) ;
assign n1106 =  ( n1071 ) ? ( iram_237 ) : ( n1105 ) ;
assign n1107 =  ( n1070 ) ? ( iram_236 ) : ( n1106 ) ;
assign n1108 =  ( n1069 ) ? ( iram_235 ) : ( n1107 ) ;
assign n1109 =  ( n1068 ) ? ( iram_234 ) : ( n1108 ) ;
assign n1110 =  ( n1067 ) ? ( iram_233 ) : ( n1109 ) ;
assign n1111 =  ( n1066 ) ? ( iram_232 ) : ( n1110 ) ;
assign n1112 =  ( n1065 ) ? ( iram_231 ) : ( n1111 ) ;
assign n1113 =  ( n1064 ) ? ( iram_230 ) : ( n1112 ) ;
assign n1114 =  ( n1063 ) ? ( iram_229 ) : ( n1113 ) ;
assign n1115 =  ( n1062 ) ? ( iram_228 ) : ( n1114 ) ;
assign n1116 =  ( n1061 ) ? ( iram_227 ) : ( n1115 ) ;
assign n1117 =  ( n1060 ) ? ( iram_226 ) : ( n1116 ) ;
assign n1118 =  ( n1059 ) ? ( iram_225 ) : ( n1117 ) ;
assign n1119 =  ( n1058 ) ? ( iram_224 ) : ( n1118 ) ;
assign n1120 =  ( n1057 ) ? ( iram_223 ) : ( n1119 ) ;
assign n1121 =  ( n1056 ) ? ( iram_222 ) : ( n1120 ) ;
assign n1122 =  ( n1055 ) ? ( iram_221 ) : ( n1121 ) ;
assign n1123 =  ( n1054 ) ? ( iram_220 ) : ( n1122 ) ;
assign n1124 =  ( n1053 ) ? ( iram_219 ) : ( n1123 ) ;
assign n1125 =  ( n1052 ) ? ( iram_218 ) : ( n1124 ) ;
assign n1126 =  ( n1051 ) ? ( iram_217 ) : ( n1125 ) ;
assign n1127 =  ( n1050 ) ? ( iram_216 ) : ( n1126 ) ;
assign n1128 =  ( n1049 ) ? ( iram_215 ) : ( n1127 ) ;
assign n1129 =  ( n1048 ) ? ( iram_214 ) : ( n1128 ) ;
assign n1130 =  ( n1047 ) ? ( iram_213 ) : ( n1129 ) ;
assign n1131 =  ( n1046 ) ? ( iram_212 ) : ( n1130 ) ;
assign n1132 =  ( n1045 ) ? ( iram_211 ) : ( n1131 ) ;
assign n1133 =  ( n1044 ) ? ( iram_210 ) : ( n1132 ) ;
assign n1134 =  ( n1043 ) ? ( iram_209 ) : ( n1133 ) ;
assign n1135 =  ( n1042 ) ? ( iram_208 ) : ( n1134 ) ;
assign n1136 =  ( n1041 ) ? ( iram_207 ) : ( n1135 ) ;
assign n1137 =  ( n1040 ) ? ( iram_206 ) : ( n1136 ) ;
assign n1138 =  ( n1039 ) ? ( iram_205 ) : ( n1137 ) ;
assign n1139 =  ( n1038 ) ? ( iram_204 ) : ( n1138 ) ;
assign n1140 =  ( n1037 ) ? ( iram_203 ) : ( n1139 ) ;
assign n1141 =  ( n1036 ) ? ( iram_202 ) : ( n1140 ) ;
assign n1142 =  ( n1035 ) ? ( iram_201 ) : ( n1141 ) ;
assign n1143 =  ( n1034 ) ? ( iram_200 ) : ( n1142 ) ;
assign n1144 =  ( n1033 ) ? ( iram_199 ) : ( n1143 ) ;
assign n1145 =  ( n1032 ) ? ( iram_198 ) : ( n1144 ) ;
assign n1146 =  ( n1031 ) ? ( iram_197 ) : ( n1145 ) ;
assign n1147 =  ( n1030 ) ? ( iram_196 ) : ( n1146 ) ;
assign n1148 =  ( n1029 ) ? ( iram_195 ) : ( n1147 ) ;
assign n1149 =  ( n1028 ) ? ( iram_194 ) : ( n1148 ) ;
assign n1150 =  ( n1027 ) ? ( iram_193 ) : ( n1149 ) ;
assign n1151 =  ( n1026 ) ? ( iram_192 ) : ( n1150 ) ;
assign n1152 =  ( n1025 ) ? ( iram_191 ) : ( n1151 ) ;
assign n1153 =  ( n1024 ) ? ( iram_190 ) : ( n1152 ) ;
assign n1154 =  ( n1023 ) ? ( iram_189 ) : ( n1153 ) ;
assign n1155 =  ( n1022 ) ? ( iram_188 ) : ( n1154 ) ;
assign n1156 =  ( n1021 ) ? ( iram_187 ) : ( n1155 ) ;
assign n1157 =  ( n1020 ) ? ( iram_186 ) : ( n1156 ) ;
assign n1158 =  ( n1019 ) ? ( iram_185 ) : ( n1157 ) ;
assign n1159 =  ( n1018 ) ? ( iram_184 ) : ( n1158 ) ;
assign n1160 =  ( n1017 ) ? ( iram_183 ) : ( n1159 ) ;
assign n1161 =  ( n1016 ) ? ( iram_182 ) : ( n1160 ) ;
assign n1162 =  ( n1015 ) ? ( iram_181 ) : ( n1161 ) ;
assign n1163 =  ( n1014 ) ? ( iram_180 ) : ( n1162 ) ;
assign n1164 =  ( n1013 ) ? ( iram_179 ) : ( n1163 ) ;
assign n1165 =  ( n1012 ) ? ( iram_178 ) : ( n1164 ) ;
assign n1166 =  ( n1011 ) ? ( iram_177 ) : ( n1165 ) ;
assign n1167 =  ( n1010 ) ? ( iram_176 ) : ( n1166 ) ;
assign n1168 =  ( n1009 ) ? ( iram_175 ) : ( n1167 ) ;
assign n1169 =  ( n1008 ) ? ( iram_174 ) : ( n1168 ) ;
assign n1170 =  ( n1007 ) ? ( iram_173 ) : ( n1169 ) ;
assign n1171 =  ( n1006 ) ? ( iram_172 ) : ( n1170 ) ;
assign n1172 =  ( n1005 ) ? ( iram_171 ) : ( n1171 ) ;
assign n1173 =  ( n1004 ) ? ( iram_170 ) : ( n1172 ) ;
assign n1174 =  ( n1003 ) ? ( iram_169 ) : ( n1173 ) ;
assign n1175 =  ( n1002 ) ? ( iram_168 ) : ( n1174 ) ;
assign n1176 =  ( n1001 ) ? ( iram_167 ) : ( n1175 ) ;
assign n1177 =  ( n1000 ) ? ( iram_166 ) : ( n1176 ) ;
assign n1178 =  ( n999 ) ? ( iram_165 ) : ( n1177 ) ;
assign n1179 =  ( n998 ) ? ( iram_164 ) : ( n1178 ) ;
assign n1180 =  ( n997 ) ? ( iram_163 ) : ( n1179 ) ;
assign n1181 =  ( n996 ) ? ( iram_162 ) : ( n1180 ) ;
assign n1182 =  ( n995 ) ? ( iram_161 ) : ( n1181 ) ;
assign n1183 =  ( n994 ) ? ( iram_160 ) : ( n1182 ) ;
assign n1184 =  ( n993 ) ? ( iram_159 ) : ( n1183 ) ;
assign n1185 =  ( n992 ) ? ( iram_158 ) : ( n1184 ) ;
assign n1186 =  ( n991 ) ? ( iram_157 ) : ( n1185 ) ;
assign n1187 =  ( n990 ) ? ( iram_156 ) : ( n1186 ) ;
assign n1188 =  ( n989 ) ? ( iram_155 ) : ( n1187 ) ;
assign n1189 =  ( n988 ) ? ( iram_154 ) : ( n1188 ) ;
assign n1190 =  ( n987 ) ? ( iram_153 ) : ( n1189 ) ;
assign n1191 =  ( n986 ) ? ( iram_152 ) : ( n1190 ) ;
assign n1192 =  ( n985 ) ? ( iram_151 ) : ( n1191 ) ;
assign n1193 =  ( n984 ) ? ( iram_150 ) : ( n1192 ) ;
assign n1194 =  ( n983 ) ? ( iram_149 ) : ( n1193 ) ;
assign n1195 =  ( n982 ) ? ( iram_148 ) : ( n1194 ) ;
assign n1196 =  ( n981 ) ? ( iram_147 ) : ( n1195 ) ;
assign n1197 =  ( n980 ) ? ( iram_146 ) : ( n1196 ) ;
assign n1198 =  ( n979 ) ? ( iram_145 ) : ( n1197 ) ;
assign n1199 =  ( n978 ) ? ( iram_144 ) : ( n1198 ) ;
assign n1200 =  ( n977 ) ? ( iram_143 ) : ( n1199 ) ;
assign n1201 =  ( n976 ) ? ( iram_142 ) : ( n1200 ) ;
assign n1202 =  ( n975 ) ? ( iram_141 ) : ( n1201 ) ;
assign n1203 =  ( n974 ) ? ( iram_140 ) : ( n1202 ) ;
assign n1204 =  ( n973 ) ? ( iram_139 ) : ( n1203 ) ;
assign n1205 =  ( n972 ) ? ( iram_138 ) : ( n1204 ) ;
assign n1206 =  ( n971 ) ? ( iram_137 ) : ( n1205 ) ;
assign n1207 =  ( n970 ) ? ( iram_136 ) : ( n1206 ) ;
assign n1208 =  ( n969 ) ? ( iram_135 ) : ( n1207 ) ;
assign n1209 =  ( n968 ) ? ( iram_134 ) : ( n1208 ) ;
assign n1210 =  ( n967 ) ? ( iram_133 ) : ( n1209 ) ;
assign n1211 =  ( n966 ) ? ( iram_132 ) : ( n1210 ) ;
assign n1212 =  ( n965 ) ? ( iram_131 ) : ( n1211 ) ;
assign n1213 =  ( n964 ) ? ( iram_130 ) : ( n1212 ) ;
assign n1214 =  ( n963 ) ? ( iram_129 ) : ( n1213 ) ;
assign n1215 =  ( n962 ) ? ( iram_128 ) : ( n1214 ) ;
assign n1216 =  ( n961 ) ? ( iram_127 ) : ( n1215 ) ;
assign n1217 =  ( n960 ) ? ( iram_126 ) : ( n1216 ) ;
assign n1218 =  ( n959 ) ? ( iram_125 ) : ( n1217 ) ;
assign n1219 =  ( n958 ) ? ( iram_124 ) : ( n1218 ) ;
assign n1220 =  ( n957 ) ? ( iram_123 ) : ( n1219 ) ;
assign n1221 =  ( n956 ) ? ( iram_122 ) : ( n1220 ) ;
assign n1222 =  ( n955 ) ? ( iram_121 ) : ( n1221 ) ;
assign n1223 =  ( n954 ) ? ( iram_120 ) : ( n1222 ) ;
assign n1224 =  ( n953 ) ? ( iram_119 ) : ( n1223 ) ;
assign n1225 =  ( n952 ) ? ( iram_118 ) : ( n1224 ) ;
assign n1226 =  ( n951 ) ? ( iram_117 ) : ( n1225 ) ;
assign n1227 =  ( n950 ) ? ( iram_116 ) : ( n1226 ) ;
assign n1228 =  ( n949 ) ? ( iram_115 ) : ( n1227 ) ;
assign n1229 =  ( n948 ) ? ( iram_114 ) : ( n1228 ) ;
assign n1230 =  ( n947 ) ? ( iram_113 ) : ( n1229 ) ;
assign n1231 =  ( n946 ) ? ( iram_112 ) : ( n1230 ) ;
assign n1232 =  ( n945 ) ? ( iram_111 ) : ( n1231 ) ;
assign n1233 =  ( n944 ) ? ( iram_110 ) : ( n1232 ) ;
assign n1234 =  ( n943 ) ? ( iram_109 ) : ( n1233 ) ;
assign n1235 =  ( n942 ) ? ( iram_108 ) : ( n1234 ) ;
assign n1236 =  ( n941 ) ? ( iram_107 ) : ( n1235 ) ;
assign n1237 =  ( n940 ) ? ( iram_106 ) : ( n1236 ) ;
assign n1238 =  ( n939 ) ? ( iram_105 ) : ( n1237 ) ;
assign n1239 =  ( n938 ) ? ( iram_104 ) : ( n1238 ) ;
assign n1240 =  ( n937 ) ? ( iram_103 ) : ( n1239 ) ;
assign n1241 =  ( n936 ) ? ( iram_102 ) : ( n1240 ) ;
assign n1242 =  ( n935 ) ? ( iram_101 ) : ( n1241 ) ;
assign n1243 =  ( n934 ) ? ( iram_100 ) : ( n1242 ) ;
assign n1244 =  ( n933 ) ? ( iram_99 ) : ( n1243 ) ;
assign n1245 =  ( n932 ) ? ( iram_98 ) : ( n1244 ) ;
assign n1246 =  ( n931 ) ? ( iram_97 ) : ( n1245 ) ;
assign n1247 =  ( n930 ) ? ( iram_96 ) : ( n1246 ) ;
assign n1248 =  ( n929 ) ? ( iram_95 ) : ( n1247 ) ;
assign n1249 =  ( n928 ) ? ( iram_94 ) : ( n1248 ) ;
assign n1250 =  ( n927 ) ? ( iram_93 ) : ( n1249 ) ;
assign n1251 =  ( n926 ) ? ( iram_92 ) : ( n1250 ) ;
assign n1252 =  ( n925 ) ? ( iram_91 ) : ( n1251 ) ;
assign n1253 =  ( n924 ) ? ( iram_90 ) : ( n1252 ) ;
assign n1254 =  ( n923 ) ? ( iram_89 ) : ( n1253 ) ;
assign n1255 =  ( n922 ) ? ( iram_88 ) : ( n1254 ) ;
assign n1256 =  ( n921 ) ? ( iram_87 ) : ( n1255 ) ;
assign n1257 =  ( n920 ) ? ( iram_86 ) : ( n1256 ) ;
assign n1258 =  ( n919 ) ? ( iram_85 ) : ( n1257 ) ;
assign n1259 =  ( n918 ) ? ( iram_84 ) : ( n1258 ) ;
assign n1260 =  ( n917 ) ? ( iram_83 ) : ( n1259 ) ;
assign n1261 =  ( n916 ) ? ( iram_82 ) : ( n1260 ) ;
assign n1262 =  ( n915 ) ? ( iram_81 ) : ( n1261 ) ;
assign n1263 =  ( n914 ) ? ( iram_80 ) : ( n1262 ) ;
assign n1264 =  ( n913 ) ? ( iram_79 ) : ( n1263 ) ;
assign n1265 =  ( n912 ) ? ( iram_78 ) : ( n1264 ) ;
assign n1266 =  ( n911 ) ? ( iram_77 ) : ( n1265 ) ;
assign n1267 =  ( n910 ) ? ( iram_76 ) : ( n1266 ) ;
assign n1268 =  ( n909 ) ? ( iram_75 ) : ( n1267 ) ;
assign n1269 =  ( n908 ) ? ( iram_74 ) : ( n1268 ) ;
assign n1270 =  ( n907 ) ? ( iram_73 ) : ( n1269 ) ;
assign n1271 =  ( n906 ) ? ( iram_72 ) : ( n1270 ) ;
assign n1272 =  ( n905 ) ? ( iram_71 ) : ( n1271 ) ;
assign n1273 =  ( n904 ) ? ( iram_70 ) : ( n1272 ) ;
assign n1274 =  ( n903 ) ? ( iram_69 ) : ( n1273 ) ;
assign n1275 =  ( n902 ) ? ( iram_68 ) : ( n1274 ) ;
assign n1276 =  ( n901 ) ? ( iram_67 ) : ( n1275 ) ;
assign n1277 =  ( n900 ) ? ( iram_66 ) : ( n1276 ) ;
assign n1278 =  ( n899 ) ? ( iram_65 ) : ( n1277 ) ;
assign n1279 =  ( n898 ) ? ( iram_64 ) : ( n1278 ) ;
assign n1280 =  ( n897 ) ? ( iram_63 ) : ( n1279 ) ;
assign n1281 =  ( n896 ) ? ( iram_62 ) : ( n1280 ) ;
assign n1282 =  ( n895 ) ? ( iram_61 ) : ( n1281 ) ;
assign n1283 =  ( n894 ) ? ( iram_60 ) : ( n1282 ) ;
assign n1284 =  ( n893 ) ? ( iram_59 ) : ( n1283 ) ;
assign n1285 =  ( n892 ) ? ( iram_58 ) : ( n1284 ) ;
assign n1286 =  ( n891 ) ? ( iram_57 ) : ( n1285 ) ;
assign n1287 =  ( n890 ) ? ( iram_56 ) : ( n1286 ) ;
assign n1288 =  ( n889 ) ? ( iram_55 ) : ( n1287 ) ;
assign n1289 =  ( n888 ) ? ( iram_54 ) : ( n1288 ) ;
assign n1290 =  ( n887 ) ? ( iram_53 ) : ( n1289 ) ;
assign n1291 =  ( n886 ) ? ( iram_52 ) : ( n1290 ) ;
assign n1292 =  ( n885 ) ? ( iram_51 ) : ( n1291 ) ;
assign n1293 =  ( n884 ) ? ( iram_50 ) : ( n1292 ) ;
assign n1294 =  ( n883 ) ? ( iram_49 ) : ( n1293 ) ;
assign n1295 =  ( n882 ) ? ( iram_48 ) : ( n1294 ) ;
assign n1296 =  ( n881 ) ? ( iram_47 ) : ( n1295 ) ;
assign n1297 =  ( n880 ) ? ( iram_46 ) : ( n1296 ) ;
assign n1298 =  ( n879 ) ? ( iram_45 ) : ( n1297 ) ;
assign n1299 =  ( n878 ) ? ( iram_44 ) : ( n1298 ) ;
assign n1300 =  ( n877 ) ? ( iram_43 ) : ( n1299 ) ;
assign n1301 =  ( n876 ) ? ( iram_42 ) : ( n1300 ) ;
assign n1302 =  ( n875 ) ? ( iram_41 ) : ( n1301 ) ;
assign n1303 =  ( n874 ) ? ( iram_40 ) : ( n1302 ) ;
assign n1304 =  ( n873 ) ? ( iram_39 ) : ( n1303 ) ;
assign n1305 =  ( n872 ) ? ( iram_38 ) : ( n1304 ) ;
assign n1306 =  ( n871 ) ? ( iram_37 ) : ( n1305 ) ;
assign n1307 =  ( n870 ) ? ( iram_36 ) : ( n1306 ) ;
assign n1308 =  ( n869 ) ? ( iram_35 ) : ( n1307 ) ;
assign n1309 =  ( n868 ) ? ( iram_34 ) : ( n1308 ) ;
assign n1310 =  ( n867 ) ? ( iram_33 ) : ( n1309 ) ;
assign n1311 =  ( n866 ) ? ( iram_32 ) : ( n1310 ) ;
assign n1312 =  ( n865 ) ? ( iram_31 ) : ( n1311 ) ;
assign n1313 =  ( n864 ) ? ( iram_30 ) : ( n1312 ) ;
assign n1314 =  ( n863 ) ? ( iram_29 ) : ( n1313 ) ;
assign n1315 =  ( n862 ) ? ( iram_28 ) : ( n1314 ) ;
assign n1316 =  ( n861 ) ? ( iram_27 ) : ( n1315 ) ;
assign n1317 =  ( n860 ) ? ( iram_26 ) : ( n1316 ) ;
assign n1318 =  ( n859 ) ? ( iram_25 ) : ( n1317 ) ;
assign n1319 =  ( n858 ) ? ( iram_24 ) : ( n1318 ) ;
assign n1320 =  ( n857 ) ? ( iram_23 ) : ( n1319 ) ;
assign n1321 =  ( n856 ) ? ( iram_22 ) : ( n1320 ) ;
assign n1322 =  ( n855 ) ? ( iram_21 ) : ( n1321 ) ;
assign n1323 =  ( n854 ) ? ( iram_20 ) : ( n1322 ) ;
assign n1324 =  ( n853 ) ? ( iram_19 ) : ( n1323 ) ;
assign n1325 =  ( n852 ) ? ( iram_18 ) : ( n1324 ) ;
assign n1326 =  ( n851 ) ? ( iram_17 ) : ( n1325 ) ;
assign n1327 =  ( n850 ) ? ( iram_16 ) : ( n1326 ) ;
assign n1328 =  ( n849 ) ? ( iram_15 ) : ( n1327 ) ;
assign n1329 =  ( n848 ) ? ( iram_14 ) : ( n1328 ) ;
assign n1330 =  ( n847 ) ? ( iram_13 ) : ( n1329 ) ;
assign n1331 =  ( n846 ) ? ( iram_12 ) : ( n1330 ) ;
assign n1332 =  ( n845 ) ? ( iram_11 ) : ( n1331 ) ;
assign n1333 =  ( n844 ) ? ( iram_10 ) : ( n1332 ) ;
assign n1334 =  ( n843 ) ? ( iram_9 ) : ( n1333 ) ;
assign n1335 =  ( n842 ) ? ( iram_8 ) : ( n1334 ) ;
assign n1336 =  ( n841 ) ? ( iram_7 ) : ( n1335 ) ;
assign n1337 =  ( n840 ) ? ( iram_6 ) : ( n1336 ) ;
assign n1338 =  ( n839 ) ? ( iram_5 ) : ( n1337 ) ;
assign n1339 =  ( n838 ) ? ( iram_4 ) : ( n1338 ) ;
assign n1340 =  ( n837 ) ? ( iram_3 ) : ( n1339 ) ;
assign n1341 =  ( n836 ) ? ( iram_2 ) : ( n1340 ) ;
assign n1342 =  ( n835 ) ? ( iram_1 ) : ( n1341 ) ;
assign n1343 =  ( n834 ) ? ( iram_0 ) : ( n1342 ) ;
assign n1344 =  ( bit_addr ) ? ( n833 ) : ( n1343 ) ;
assign n1345 = rd_addr[7:7] ;
assign n1346 =  ( n1345 ) == ( bv_1_1_n34 )  ;
assign n1347 = rd_addr[6:3] ;
assign n1348 =  { ( bv_1_1_n34 ) , ( n1347 ) }  ;
assign n1349 =  { ( n1348 ) , ( bv_3_0_n46 ) }  ;
assign n1350 = rd_addr[6:3] ;
assign n1351 =  { ( bv_4_2_n12 ) , ( n1350 ) }  ;
assign n1352 =  ( n1346 ) ? ( n1349 ) : ( n1351 ) ;
assign n1353 =  ( bit_addr ) ? ( n1352 ) : ( rd_addr ) ;
assign n1354 = n1353[7:0] ;
assign n1355 =  ( n1354 ) == ( bv_8_0_n69 )  ;
assign n1356 =  ( n1354 ) == ( bv_8_1_n71 )  ;
assign n1357 =  ( n1354 ) == ( bv_8_2_n73 )  ;
assign n1358 =  ( n1354 ) == ( bv_8_3_n75 )  ;
assign n1359 =  ( n1354 ) == ( bv_8_4_n77 )  ;
assign n1360 =  ( n1354 ) == ( bv_8_5_n79 )  ;
assign n1361 =  ( n1354 ) == ( bv_8_6_n81 )  ;
assign n1362 =  ( n1354 ) == ( bv_8_7_n83 )  ;
assign n1363 =  ( n1354 ) == ( bv_8_8_n85 )  ;
assign n1364 =  ( n1354 ) == ( bv_8_9_n87 )  ;
assign n1365 =  ( n1354 ) == ( bv_8_10_n89 )  ;
assign n1366 =  ( n1354 ) == ( bv_8_11_n91 )  ;
assign n1367 =  ( n1354 ) == ( bv_8_12_n93 )  ;
assign n1368 =  ( n1354 ) == ( bv_8_13_n95 )  ;
assign n1369 =  ( n1354 ) == ( bv_8_14_n97 )  ;
assign n1370 =  ( n1354 ) == ( bv_8_15_n99 )  ;
assign n1371 =  ( n1354 ) == ( bv_8_16_n101 )  ;
assign n1372 =  ( n1354 ) == ( bv_8_17_n103 )  ;
assign n1373 =  ( n1354 ) == ( bv_8_18_n105 )  ;
assign n1374 =  ( n1354 ) == ( bv_8_19_n107 )  ;
assign n1375 =  ( n1354 ) == ( bv_8_20_n109 )  ;
assign n1376 =  ( n1354 ) == ( bv_8_21_n111 )  ;
assign n1377 =  ( n1354 ) == ( bv_8_22_n113 )  ;
assign n1378 =  ( n1354 ) == ( bv_8_23_n115 )  ;
assign n1379 =  ( n1354 ) == ( bv_8_24_n117 )  ;
assign n1380 =  ( n1354 ) == ( bv_8_25_n119 )  ;
assign n1381 =  ( n1354 ) == ( bv_8_26_n121 )  ;
assign n1382 =  ( n1354 ) == ( bv_8_27_n123 )  ;
assign n1383 =  ( n1354 ) == ( bv_8_28_n125 )  ;
assign n1384 =  ( n1354 ) == ( bv_8_29_n127 )  ;
assign n1385 =  ( n1354 ) == ( bv_8_30_n129 )  ;
assign n1386 =  ( n1354 ) == ( bv_8_31_n131 )  ;
assign n1387 =  ( n1354 ) == ( bv_8_32_n133 )  ;
assign n1388 =  ( n1354 ) == ( bv_8_33_n135 )  ;
assign n1389 =  ( n1354 ) == ( bv_8_34_n137 )  ;
assign n1390 =  ( n1354 ) == ( bv_8_35_n139 )  ;
assign n1391 =  ( n1354 ) == ( bv_8_36_n141 )  ;
assign n1392 =  ( n1354 ) == ( bv_8_37_n143 )  ;
assign n1393 =  ( n1354 ) == ( bv_8_38_n145 )  ;
assign n1394 =  ( n1354 ) == ( bv_8_39_n147 )  ;
assign n1395 =  ( n1354 ) == ( bv_8_40_n149 )  ;
assign n1396 =  ( n1354 ) == ( bv_8_41_n151 )  ;
assign n1397 =  ( n1354 ) == ( bv_8_42_n153 )  ;
assign n1398 =  ( n1354 ) == ( bv_8_43_n155 )  ;
assign n1399 =  ( n1354 ) == ( bv_8_44_n157 )  ;
assign n1400 =  ( n1354 ) == ( bv_8_45_n159 )  ;
assign n1401 =  ( n1354 ) == ( bv_8_46_n161 )  ;
assign n1402 =  ( n1354 ) == ( bv_8_47_n163 )  ;
assign n1403 =  ( n1354 ) == ( bv_8_48_n165 )  ;
assign n1404 =  ( n1354 ) == ( bv_8_49_n167 )  ;
assign n1405 =  ( n1354 ) == ( bv_8_50_n169 )  ;
assign n1406 =  ( n1354 ) == ( bv_8_51_n171 )  ;
assign n1407 =  ( n1354 ) == ( bv_8_52_n173 )  ;
assign n1408 =  ( n1354 ) == ( bv_8_53_n175 )  ;
assign n1409 =  ( n1354 ) == ( bv_8_54_n177 )  ;
assign n1410 =  ( n1354 ) == ( bv_8_55_n179 )  ;
assign n1411 =  ( n1354 ) == ( bv_8_56_n181 )  ;
assign n1412 =  ( n1354 ) == ( bv_8_57_n183 )  ;
assign n1413 =  ( n1354 ) == ( bv_8_58_n185 )  ;
assign n1414 =  ( n1354 ) == ( bv_8_59_n187 )  ;
assign n1415 =  ( n1354 ) == ( bv_8_60_n189 )  ;
assign n1416 =  ( n1354 ) == ( bv_8_61_n191 )  ;
assign n1417 =  ( n1354 ) == ( bv_8_62_n193 )  ;
assign n1418 =  ( n1354 ) == ( bv_8_63_n195 )  ;
assign n1419 =  ( n1354 ) == ( bv_8_64_n197 )  ;
assign n1420 =  ( n1354 ) == ( bv_8_65_n199 )  ;
assign n1421 =  ( n1354 ) == ( bv_8_66_n201 )  ;
assign n1422 =  ( n1354 ) == ( bv_8_67_n203 )  ;
assign n1423 =  ( n1354 ) == ( bv_8_68_n205 )  ;
assign n1424 =  ( n1354 ) == ( bv_8_69_n207 )  ;
assign n1425 =  ( n1354 ) == ( bv_8_70_n209 )  ;
assign n1426 =  ( n1354 ) == ( bv_8_71_n211 )  ;
assign n1427 =  ( n1354 ) == ( bv_8_72_n213 )  ;
assign n1428 =  ( n1354 ) == ( bv_8_73_n215 )  ;
assign n1429 =  ( n1354 ) == ( bv_8_74_n217 )  ;
assign n1430 =  ( n1354 ) == ( bv_8_75_n219 )  ;
assign n1431 =  ( n1354 ) == ( bv_8_76_n221 )  ;
assign n1432 =  ( n1354 ) == ( bv_8_77_n223 )  ;
assign n1433 =  ( n1354 ) == ( bv_8_78_n225 )  ;
assign n1434 =  ( n1354 ) == ( bv_8_79_n227 )  ;
assign n1435 =  ( n1354 ) == ( bv_8_80_n229 )  ;
assign n1436 =  ( n1354 ) == ( bv_8_81_n231 )  ;
assign n1437 =  ( n1354 ) == ( bv_8_82_n233 )  ;
assign n1438 =  ( n1354 ) == ( bv_8_83_n235 )  ;
assign n1439 =  ( n1354 ) == ( bv_8_84_n237 )  ;
assign n1440 =  ( n1354 ) == ( bv_8_85_n239 )  ;
assign n1441 =  ( n1354 ) == ( bv_8_86_n241 )  ;
assign n1442 =  ( n1354 ) == ( bv_8_87_n243 )  ;
assign n1443 =  ( n1354 ) == ( bv_8_88_n245 )  ;
assign n1444 =  ( n1354 ) == ( bv_8_89_n247 )  ;
assign n1445 =  ( n1354 ) == ( bv_8_90_n249 )  ;
assign n1446 =  ( n1354 ) == ( bv_8_91_n251 )  ;
assign n1447 =  ( n1354 ) == ( bv_8_92_n253 )  ;
assign n1448 =  ( n1354 ) == ( bv_8_93_n255 )  ;
assign n1449 =  ( n1354 ) == ( bv_8_94_n257 )  ;
assign n1450 =  ( n1354 ) == ( bv_8_95_n259 )  ;
assign n1451 =  ( n1354 ) == ( bv_8_96_n261 )  ;
assign n1452 =  ( n1354 ) == ( bv_8_97_n263 )  ;
assign n1453 =  ( n1354 ) == ( bv_8_98_n265 )  ;
assign n1454 =  ( n1354 ) == ( bv_8_99_n267 )  ;
assign n1455 =  ( n1354 ) == ( bv_8_100_n269 )  ;
assign n1456 =  ( n1354 ) == ( bv_8_101_n271 )  ;
assign n1457 =  ( n1354 ) == ( bv_8_102_n273 )  ;
assign n1458 =  ( n1354 ) == ( bv_8_103_n275 )  ;
assign n1459 =  ( n1354 ) == ( bv_8_104_n277 )  ;
assign n1460 =  ( n1354 ) == ( bv_8_105_n279 )  ;
assign n1461 =  ( n1354 ) == ( bv_8_106_n281 )  ;
assign n1462 =  ( n1354 ) == ( bv_8_107_n283 )  ;
assign n1463 =  ( n1354 ) == ( bv_8_108_n285 )  ;
assign n1464 =  ( n1354 ) == ( bv_8_109_n287 )  ;
assign n1465 =  ( n1354 ) == ( bv_8_110_n289 )  ;
assign n1466 =  ( n1354 ) == ( bv_8_111_n291 )  ;
assign n1467 =  ( n1354 ) == ( bv_8_112_n293 )  ;
assign n1468 =  ( n1354 ) == ( bv_8_113_n295 )  ;
assign n1469 =  ( n1354 ) == ( bv_8_114_n297 )  ;
assign n1470 =  ( n1354 ) == ( bv_8_115_n299 )  ;
assign n1471 =  ( n1354 ) == ( bv_8_116_n301 )  ;
assign n1472 =  ( n1354 ) == ( bv_8_117_n303 )  ;
assign n1473 =  ( n1354 ) == ( bv_8_118_n305 )  ;
assign n1474 =  ( n1354 ) == ( bv_8_119_n307 )  ;
assign n1475 =  ( n1354 ) == ( bv_8_120_n309 )  ;
assign n1476 =  ( n1354 ) == ( bv_8_121_n311 )  ;
assign n1477 =  ( n1354 ) == ( bv_8_122_n313 )  ;
assign n1478 =  ( n1354 ) == ( bv_8_123_n315 )  ;
assign n1479 =  ( n1354 ) == ( bv_8_124_n317 )  ;
assign n1480 =  ( n1354 ) == ( bv_8_125_n319 )  ;
assign n1481 =  ( n1354 ) == ( bv_8_126_n321 )  ;
assign n1482 =  ( n1354 ) == ( bv_8_127_n323 )  ;
assign n1483 =  ( n1354 ) == ( bv_8_128_n325 )  ;
assign n1484 =  ( n1354 ) == ( bv_8_129_n327 )  ;
assign n1485 =  ( n1354 ) == ( bv_8_130_n329 )  ;
assign n1486 =  ( n1354 ) == ( bv_8_131_n331 )  ;
assign n1487 =  ( n1354 ) == ( bv_8_132_n333 )  ;
assign n1488 =  ( n1354 ) == ( bv_8_133_n335 )  ;
assign n1489 =  ( n1354 ) == ( bv_8_134_n337 )  ;
assign n1490 =  ( n1354 ) == ( bv_8_135_n339 )  ;
assign n1491 =  ( n1354 ) == ( bv_8_136_n341 )  ;
assign n1492 =  ( n1354 ) == ( bv_8_137_n343 )  ;
assign n1493 =  ( n1354 ) == ( bv_8_138_n345 )  ;
assign n1494 =  ( n1354 ) == ( bv_8_139_n347 )  ;
assign n1495 =  ( n1354 ) == ( bv_8_140_n349 )  ;
assign n1496 =  ( n1354 ) == ( bv_8_141_n351 )  ;
assign n1497 =  ( n1354 ) == ( bv_8_142_n353 )  ;
assign n1498 =  ( n1354 ) == ( bv_8_143_n355 )  ;
assign n1499 =  ( n1354 ) == ( bv_8_144_n357 )  ;
assign n1500 =  ( n1354 ) == ( bv_8_145_n359 )  ;
assign n1501 =  ( n1354 ) == ( bv_8_146_n361 )  ;
assign n1502 =  ( n1354 ) == ( bv_8_147_n363 )  ;
assign n1503 =  ( n1354 ) == ( bv_8_148_n365 )  ;
assign n1504 =  ( n1354 ) == ( bv_8_149_n367 )  ;
assign n1505 =  ( n1354 ) == ( bv_8_150_n369 )  ;
assign n1506 =  ( n1354 ) == ( bv_8_151_n371 )  ;
assign n1507 =  ( n1354 ) == ( bv_8_152_n373 )  ;
assign n1508 =  ( n1354 ) == ( bv_8_153_n375 )  ;
assign n1509 =  ( n1354 ) == ( bv_8_154_n377 )  ;
assign n1510 =  ( n1354 ) == ( bv_8_155_n379 )  ;
assign n1511 =  ( n1354 ) == ( bv_8_156_n381 )  ;
assign n1512 =  ( n1354 ) == ( bv_8_157_n383 )  ;
assign n1513 =  ( n1354 ) == ( bv_8_158_n385 )  ;
assign n1514 =  ( n1354 ) == ( bv_8_159_n387 )  ;
assign n1515 =  ( n1354 ) == ( bv_8_160_n389 )  ;
assign n1516 =  ( n1354 ) == ( bv_8_161_n391 )  ;
assign n1517 =  ( n1354 ) == ( bv_8_162_n393 )  ;
assign n1518 =  ( n1354 ) == ( bv_8_163_n395 )  ;
assign n1519 =  ( n1354 ) == ( bv_8_164_n397 )  ;
assign n1520 =  ( n1354 ) == ( bv_8_165_n399 )  ;
assign n1521 =  ( n1354 ) == ( bv_8_166_n401 )  ;
assign n1522 =  ( n1354 ) == ( bv_8_167_n403 )  ;
assign n1523 =  ( n1354 ) == ( bv_8_168_n405 )  ;
assign n1524 =  ( n1354 ) == ( bv_8_169_n407 )  ;
assign n1525 =  ( n1354 ) == ( bv_8_170_n409 )  ;
assign n1526 =  ( n1354 ) == ( bv_8_171_n411 )  ;
assign n1527 =  ( n1354 ) == ( bv_8_172_n413 )  ;
assign n1528 =  ( n1354 ) == ( bv_8_173_n415 )  ;
assign n1529 =  ( n1354 ) == ( bv_8_174_n417 )  ;
assign n1530 =  ( n1354 ) == ( bv_8_175_n419 )  ;
assign n1531 =  ( n1354 ) == ( bv_8_176_n421 )  ;
assign n1532 =  ( n1354 ) == ( bv_8_177_n423 )  ;
assign n1533 =  ( n1354 ) == ( bv_8_178_n425 )  ;
assign n1534 =  ( n1354 ) == ( bv_8_179_n427 )  ;
assign n1535 =  ( n1354 ) == ( bv_8_180_n429 )  ;
assign n1536 =  ( n1354 ) == ( bv_8_181_n431 )  ;
assign n1537 =  ( n1354 ) == ( bv_8_182_n433 )  ;
assign n1538 =  ( n1354 ) == ( bv_8_183_n435 )  ;
assign n1539 =  ( n1354 ) == ( bv_8_184_n437 )  ;
assign n1540 =  ( n1354 ) == ( bv_8_185_n439 )  ;
assign n1541 =  ( n1354 ) == ( bv_8_186_n441 )  ;
assign n1542 =  ( n1354 ) == ( bv_8_187_n443 )  ;
assign n1543 =  ( n1354 ) == ( bv_8_188_n445 )  ;
assign n1544 =  ( n1354 ) == ( bv_8_189_n447 )  ;
assign n1545 =  ( n1354 ) == ( bv_8_190_n449 )  ;
assign n1546 =  ( n1354 ) == ( bv_8_191_n451 )  ;
assign n1547 =  ( n1354 ) == ( bv_8_192_n453 )  ;
assign n1548 =  ( n1354 ) == ( bv_8_193_n455 )  ;
assign n1549 =  ( n1354 ) == ( bv_8_194_n457 )  ;
assign n1550 =  ( n1354 ) == ( bv_8_195_n459 )  ;
assign n1551 =  ( n1354 ) == ( bv_8_196_n461 )  ;
assign n1552 =  ( n1354 ) == ( bv_8_197_n463 )  ;
assign n1553 =  ( n1354 ) == ( bv_8_198_n465 )  ;
assign n1554 =  ( n1354 ) == ( bv_8_199_n467 )  ;
assign n1555 =  ( n1354 ) == ( bv_8_200_n469 )  ;
assign n1556 =  ( n1354 ) == ( bv_8_201_n471 )  ;
assign n1557 =  ( n1354 ) == ( bv_8_202_n473 )  ;
assign n1558 =  ( n1354 ) == ( bv_8_203_n475 )  ;
assign n1559 =  ( n1354 ) == ( bv_8_204_n477 )  ;
assign n1560 =  ( n1354 ) == ( bv_8_205_n479 )  ;
assign n1561 =  ( n1354 ) == ( bv_8_206_n481 )  ;
assign n1562 =  ( n1354 ) == ( bv_8_207_n483 )  ;
assign n1563 =  ( n1354 ) == ( bv_8_208_n485 )  ;
assign n1564 =  ( n1354 ) == ( bv_8_209_n487 )  ;
assign n1565 =  ( n1354 ) == ( bv_8_210_n489 )  ;
assign n1566 =  ( n1354 ) == ( bv_8_211_n491 )  ;
assign n1567 =  ( n1354 ) == ( bv_8_212_n493 )  ;
assign n1568 =  ( n1354 ) == ( bv_8_213_n495 )  ;
assign n1569 =  ( n1354 ) == ( bv_8_214_n497 )  ;
assign n1570 =  ( n1354 ) == ( bv_8_215_n499 )  ;
assign n1571 =  ( n1354 ) == ( bv_8_216_n501 )  ;
assign n1572 =  ( n1354 ) == ( bv_8_217_n503 )  ;
assign n1573 =  ( n1354 ) == ( bv_8_218_n505 )  ;
assign n1574 =  ( n1354 ) == ( bv_8_219_n507 )  ;
assign n1575 =  ( n1354 ) == ( bv_8_220_n509 )  ;
assign n1576 =  ( n1354 ) == ( bv_8_221_n511 )  ;
assign n1577 =  ( n1354 ) == ( bv_8_222_n513 )  ;
assign n1578 =  ( n1354 ) == ( bv_8_223_n515 )  ;
assign n1579 =  ( n1354 ) == ( bv_8_224_n517 )  ;
assign n1580 =  ( n1354 ) == ( bv_8_225_n519 )  ;
assign n1581 =  ( n1354 ) == ( bv_8_226_n521 )  ;
assign n1582 =  ( n1354 ) == ( bv_8_227_n523 )  ;
assign n1583 =  ( n1354 ) == ( bv_8_228_n525 )  ;
assign n1584 =  ( n1354 ) == ( bv_8_229_n527 )  ;
assign n1585 =  ( n1354 ) == ( bv_8_230_n529 )  ;
assign n1586 =  ( n1354 ) == ( bv_8_231_n531 )  ;
assign n1587 =  ( n1354 ) == ( bv_8_232_n533 )  ;
assign n1588 =  ( n1354 ) == ( bv_8_233_n535 )  ;
assign n1589 =  ( n1354 ) == ( bv_8_234_n537 )  ;
assign n1590 =  ( n1354 ) == ( bv_8_235_n539 )  ;
assign n1591 =  ( n1354 ) == ( bv_8_236_n541 )  ;
assign n1592 =  ( n1354 ) == ( bv_8_237_n543 )  ;
assign n1593 =  ( n1354 ) == ( bv_8_238_n545 )  ;
assign n1594 =  ( n1354 ) == ( bv_8_239_n547 )  ;
assign n1595 =  ( n1354 ) == ( bv_8_240_n549 )  ;
assign n1596 =  ( n1354 ) == ( bv_8_241_n551 )  ;
assign n1597 =  ( n1354 ) == ( bv_8_242_n553 )  ;
assign n1598 =  ( n1354 ) == ( bv_8_243_n555 )  ;
assign n1599 =  ( n1354 ) == ( bv_8_244_n557 )  ;
assign n1600 =  ( n1354 ) == ( bv_8_245_n559 )  ;
assign n1601 =  ( n1354 ) == ( bv_8_246_n561 )  ;
assign n1602 =  ( n1354 ) == ( bv_8_247_n563 )  ;
assign n1603 =  ( n1354 ) == ( bv_8_248_n565 )  ;
assign n1604 =  ( n1354 ) == ( bv_8_249_n567 )  ;
assign n1605 =  ( n1354 ) == ( bv_8_250_n569 )  ;
assign n1606 =  ( n1354 ) == ( bv_8_251_n571 )  ;
assign n1607 =  ( n1354 ) == ( bv_8_252_n573 )  ;
assign n1608 =  ( n1354 ) == ( bv_8_253_n575 )  ;
assign n1609 =  ( n1354 ) == ( bv_8_254_n577 )  ;
assign n1610 =  ( n1609 ) ? ( iram_254 ) : ( iram_255 ) ;
assign n1611 =  ( n1608 ) ? ( iram_253 ) : ( n1610 ) ;
assign n1612 =  ( n1607 ) ? ( iram_252 ) : ( n1611 ) ;
assign n1613 =  ( n1606 ) ? ( iram_251 ) : ( n1612 ) ;
assign n1614 =  ( n1605 ) ? ( iram_250 ) : ( n1613 ) ;
assign n1615 =  ( n1604 ) ? ( iram_249 ) : ( n1614 ) ;
assign n1616 =  ( n1603 ) ? ( iram_248 ) : ( n1615 ) ;
assign n1617 =  ( n1602 ) ? ( iram_247 ) : ( n1616 ) ;
assign n1618 =  ( n1601 ) ? ( iram_246 ) : ( n1617 ) ;
assign n1619 =  ( n1600 ) ? ( iram_245 ) : ( n1618 ) ;
assign n1620 =  ( n1599 ) ? ( iram_244 ) : ( n1619 ) ;
assign n1621 =  ( n1598 ) ? ( iram_243 ) : ( n1620 ) ;
assign n1622 =  ( n1597 ) ? ( iram_242 ) : ( n1621 ) ;
assign n1623 =  ( n1596 ) ? ( iram_241 ) : ( n1622 ) ;
assign n1624 =  ( n1595 ) ? ( iram_240 ) : ( n1623 ) ;
assign n1625 =  ( n1594 ) ? ( iram_239 ) : ( n1624 ) ;
assign n1626 =  ( n1593 ) ? ( iram_238 ) : ( n1625 ) ;
assign n1627 =  ( n1592 ) ? ( iram_237 ) : ( n1626 ) ;
assign n1628 =  ( n1591 ) ? ( iram_236 ) : ( n1627 ) ;
assign n1629 =  ( n1590 ) ? ( iram_235 ) : ( n1628 ) ;
assign n1630 =  ( n1589 ) ? ( iram_234 ) : ( n1629 ) ;
assign n1631 =  ( n1588 ) ? ( iram_233 ) : ( n1630 ) ;
assign n1632 =  ( n1587 ) ? ( iram_232 ) : ( n1631 ) ;
assign n1633 =  ( n1586 ) ? ( iram_231 ) : ( n1632 ) ;
assign n1634 =  ( n1585 ) ? ( iram_230 ) : ( n1633 ) ;
assign n1635 =  ( n1584 ) ? ( iram_229 ) : ( n1634 ) ;
assign n1636 =  ( n1583 ) ? ( iram_228 ) : ( n1635 ) ;
assign n1637 =  ( n1582 ) ? ( iram_227 ) : ( n1636 ) ;
assign n1638 =  ( n1581 ) ? ( iram_226 ) : ( n1637 ) ;
assign n1639 =  ( n1580 ) ? ( iram_225 ) : ( n1638 ) ;
assign n1640 =  ( n1579 ) ? ( iram_224 ) : ( n1639 ) ;
assign n1641 =  ( n1578 ) ? ( iram_223 ) : ( n1640 ) ;
assign n1642 =  ( n1577 ) ? ( iram_222 ) : ( n1641 ) ;
assign n1643 =  ( n1576 ) ? ( iram_221 ) : ( n1642 ) ;
assign n1644 =  ( n1575 ) ? ( iram_220 ) : ( n1643 ) ;
assign n1645 =  ( n1574 ) ? ( iram_219 ) : ( n1644 ) ;
assign n1646 =  ( n1573 ) ? ( iram_218 ) : ( n1645 ) ;
assign n1647 =  ( n1572 ) ? ( iram_217 ) : ( n1646 ) ;
assign n1648 =  ( n1571 ) ? ( iram_216 ) : ( n1647 ) ;
assign n1649 =  ( n1570 ) ? ( iram_215 ) : ( n1648 ) ;
assign n1650 =  ( n1569 ) ? ( iram_214 ) : ( n1649 ) ;
assign n1651 =  ( n1568 ) ? ( iram_213 ) : ( n1650 ) ;
assign n1652 =  ( n1567 ) ? ( iram_212 ) : ( n1651 ) ;
assign n1653 =  ( n1566 ) ? ( iram_211 ) : ( n1652 ) ;
assign n1654 =  ( n1565 ) ? ( iram_210 ) : ( n1653 ) ;
assign n1655 =  ( n1564 ) ? ( iram_209 ) : ( n1654 ) ;
assign n1656 =  ( n1563 ) ? ( iram_208 ) : ( n1655 ) ;
assign n1657 =  ( n1562 ) ? ( iram_207 ) : ( n1656 ) ;
assign n1658 =  ( n1561 ) ? ( iram_206 ) : ( n1657 ) ;
assign n1659 =  ( n1560 ) ? ( iram_205 ) : ( n1658 ) ;
assign n1660 =  ( n1559 ) ? ( iram_204 ) : ( n1659 ) ;
assign n1661 =  ( n1558 ) ? ( iram_203 ) : ( n1660 ) ;
assign n1662 =  ( n1557 ) ? ( iram_202 ) : ( n1661 ) ;
assign n1663 =  ( n1556 ) ? ( iram_201 ) : ( n1662 ) ;
assign n1664 =  ( n1555 ) ? ( iram_200 ) : ( n1663 ) ;
assign n1665 =  ( n1554 ) ? ( iram_199 ) : ( n1664 ) ;
assign n1666 =  ( n1553 ) ? ( iram_198 ) : ( n1665 ) ;
assign n1667 =  ( n1552 ) ? ( iram_197 ) : ( n1666 ) ;
assign n1668 =  ( n1551 ) ? ( iram_196 ) : ( n1667 ) ;
assign n1669 =  ( n1550 ) ? ( iram_195 ) : ( n1668 ) ;
assign n1670 =  ( n1549 ) ? ( iram_194 ) : ( n1669 ) ;
assign n1671 =  ( n1548 ) ? ( iram_193 ) : ( n1670 ) ;
assign n1672 =  ( n1547 ) ? ( iram_192 ) : ( n1671 ) ;
assign n1673 =  ( n1546 ) ? ( iram_191 ) : ( n1672 ) ;
assign n1674 =  ( n1545 ) ? ( iram_190 ) : ( n1673 ) ;
assign n1675 =  ( n1544 ) ? ( iram_189 ) : ( n1674 ) ;
assign n1676 =  ( n1543 ) ? ( iram_188 ) : ( n1675 ) ;
assign n1677 =  ( n1542 ) ? ( iram_187 ) : ( n1676 ) ;
assign n1678 =  ( n1541 ) ? ( iram_186 ) : ( n1677 ) ;
assign n1679 =  ( n1540 ) ? ( iram_185 ) : ( n1678 ) ;
assign n1680 =  ( n1539 ) ? ( iram_184 ) : ( n1679 ) ;
assign n1681 =  ( n1538 ) ? ( iram_183 ) : ( n1680 ) ;
assign n1682 =  ( n1537 ) ? ( iram_182 ) : ( n1681 ) ;
assign n1683 =  ( n1536 ) ? ( iram_181 ) : ( n1682 ) ;
assign n1684 =  ( n1535 ) ? ( iram_180 ) : ( n1683 ) ;
assign n1685 =  ( n1534 ) ? ( iram_179 ) : ( n1684 ) ;
assign n1686 =  ( n1533 ) ? ( iram_178 ) : ( n1685 ) ;
assign n1687 =  ( n1532 ) ? ( iram_177 ) : ( n1686 ) ;
assign n1688 =  ( n1531 ) ? ( iram_176 ) : ( n1687 ) ;
assign n1689 =  ( n1530 ) ? ( iram_175 ) : ( n1688 ) ;
assign n1690 =  ( n1529 ) ? ( iram_174 ) : ( n1689 ) ;
assign n1691 =  ( n1528 ) ? ( iram_173 ) : ( n1690 ) ;
assign n1692 =  ( n1527 ) ? ( iram_172 ) : ( n1691 ) ;
assign n1693 =  ( n1526 ) ? ( iram_171 ) : ( n1692 ) ;
assign n1694 =  ( n1525 ) ? ( iram_170 ) : ( n1693 ) ;
assign n1695 =  ( n1524 ) ? ( iram_169 ) : ( n1694 ) ;
assign n1696 =  ( n1523 ) ? ( iram_168 ) : ( n1695 ) ;
assign n1697 =  ( n1522 ) ? ( iram_167 ) : ( n1696 ) ;
assign n1698 =  ( n1521 ) ? ( iram_166 ) : ( n1697 ) ;
assign n1699 =  ( n1520 ) ? ( iram_165 ) : ( n1698 ) ;
assign n1700 =  ( n1519 ) ? ( iram_164 ) : ( n1699 ) ;
assign n1701 =  ( n1518 ) ? ( iram_163 ) : ( n1700 ) ;
assign n1702 =  ( n1517 ) ? ( iram_162 ) : ( n1701 ) ;
assign n1703 =  ( n1516 ) ? ( iram_161 ) : ( n1702 ) ;
assign n1704 =  ( n1515 ) ? ( iram_160 ) : ( n1703 ) ;
assign n1705 =  ( n1514 ) ? ( iram_159 ) : ( n1704 ) ;
assign n1706 =  ( n1513 ) ? ( iram_158 ) : ( n1705 ) ;
assign n1707 =  ( n1512 ) ? ( iram_157 ) : ( n1706 ) ;
assign n1708 =  ( n1511 ) ? ( iram_156 ) : ( n1707 ) ;
assign n1709 =  ( n1510 ) ? ( iram_155 ) : ( n1708 ) ;
assign n1710 =  ( n1509 ) ? ( iram_154 ) : ( n1709 ) ;
assign n1711 =  ( n1508 ) ? ( iram_153 ) : ( n1710 ) ;
assign n1712 =  ( n1507 ) ? ( iram_152 ) : ( n1711 ) ;
assign n1713 =  ( n1506 ) ? ( iram_151 ) : ( n1712 ) ;
assign n1714 =  ( n1505 ) ? ( iram_150 ) : ( n1713 ) ;
assign n1715 =  ( n1504 ) ? ( iram_149 ) : ( n1714 ) ;
assign n1716 =  ( n1503 ) ? ( iram_148 ) : ( n1715 ) ;
assign n1717 =  ( n1502 ) ? ( iram_147 ) : ( n1716 ) ;
assign n1718 =  ( n1501 ) ? ( iram_146 ) : ( n1717 ) ;
assign n1719 =  ( n1500 ) ? ( iram_145 ) : ( n1718 ) ;
assign n1720 =  ( n1499 ) ? ( iram_144 ) : ( n1719 ) ;
assign n1721 =  ( n1498 ) ? ( iram_143 ) : ( n1720 ) ;
assign n1722 =  ( n1497 ) ? ( iram_142 ) : ( n1721 ) ;
assign n1723 =  ( n1496 ) ? ( iram_141 ) : ( n1722 ) ;
assign n1724 =  ( n1495 ) ? ( iram_140 ) : ( n1723 ) ;
assign n1725 =  ( n1494 ) ? ( iram_139 ) : ( n1724 ) ;
assign n1726 =  ( n1493 ) ? ( iram_138 ) : ( n1725 ) ;
assign n1727 =  ( n1492 ) ? ( iram_137 ) : ( n1726 ) ;
assign n1728 =  ( n1491 ) ? ( iram_136 ) : ( n1727 ) ;
assign n1729 =  ( n1490 ) ? ( iram_135 ) : ( n1728 ) ;
assign n1730 =  ( n1489 ) ? ( iram_134 ) : ( n1729 ) ;
assign n1731 =  ( n1488 ) ? ( iram_133 ) : ( n1730 ) ;
assign n1732 =  ( n1487 ) ? ( iram_132 ) : ( n1731 ) ;
assign n1733 =  ( n1486 ) ? ( iram_131 ) : ( n1732 ) ;
assign n1734 =  ( n1485 ) ? ( iram_130 ) : ( n1733 ) ;
assign n1735 =  ( n1484 ) ? ( iram_129 ) : ( n1734 ) ;
assign n1736 =  ( n1483 ) ? ( iram_128 ) : ( n1735 ) ;
assign n1737 =  ( n1482 ) ? ( iram_127 ) : ( n1736 ) ;
assign n1738 =  ( n1481 ) ? ( iram_126 ) : ( n1737 ) ;
assign n1739 =  ( n1480 ) ? ( iram_125 ) : ( n1738 ) ;
assign n1740 =  ( n1479 ) ? ( iram_124 ) : ( n1739 ) ;
assign n1741 =  ( n1478 ) ? ( iram_123 ) : ( n1740 ) ;
assign n1742 =  ( n1477 ) ? ( iram_122 ) : ( n1741 ) ;
assign n1743 =  ( n1476 ) ? ( iram_121 ) : ( n1742 ) ;
assign n1744 =  ( n1475 ) ? ( iram_120 ) : ( n1743 ) ;
assign n1745 =  ( n1474 ) ? ( iram_119 ) : ( n1744 ) ;
assign n1746 =  ( n1473 ) ? ( iram_118 ) : ( n1745 ) ;
assign n1747 =  ( n1472 ) ? ( iram_117 ) : ( n1746 ) ;
assign n1748 =  ( n1471 ) ? ( iram_116 ) : ( n1747 ) ;
assign n1749 =  ( n1470 ) ? ( iram_115 ) : ( n1748 ) ;
assign n1750 =  ( n1469 ) ? ( iram_114 ) : ( n1749 ) ;
assign n1751 =  ( n1468 ) ? ( iram_113 ) : ( n1750 ) ;
assign n1752 =  ( n1467 ) ? ( iram_112 ) : ( n1751 ) ;
assign n1753 =  ( n1466 ) ? ( iram_111 ) : ( n1752 ) ;
assign n1754 =  ( n1465 ) ? ( iram_110 ) : ( n1753 ) ;
assign n1755 =  ( n1464 ) ? ( iram_109 ) : ( n1754 ) ;
assign n1756 =  ( n1463 ) ? ( iram_108 ) : ( n1755 ) ;
assign n1757 =  ( n1462 ) ? ( iram_107 ) : ( n1756 ) ;
assign n1758 =  ( n1461 ) ? ( iram_106 ) : ( n1757 ) ;
assign n1759 =  ( n1460 ) ? ( iram_105 ) : ( n1758 ) ;
assign n1760 =  ( n1459 ) ? ( iram_104 ) : ( n1759 ) ;
assign n1761 =  ( n1458 ) ? ( iram_103 ) : ( n1760 ) ;
assign n1762 =  ( n1457 ) ? ( iram_102 ) : ( n1761 ) ;
assign n1763 =  ( n1456 ) ? ( iram_101 ) : ( n1762 ) ;
assign n1764 =  ( n1455 ) ? ( iram_100 ) : ( n1763 ) ;
assign n1765 =  ( n1454 ) ? ( iram_99 ) : ( n1764 ) ;
assign n1766 =  ( n1453 ) ? ( iram_98 ) : ( n1765 ) ;
assign n1767 =  ( n1452 ) ? ( iram_97 ) : ( n1766 ) ;
assign n1768 =  ( n1451 ) ? ( iram_96 ) : ( n1767 ) ;
assign n1769 =  ( n1450 ) ? ( iram_95 ) : ( n1768 ) ;
assign n1770 =  ( n1449 ) ? ( iram_94 ) : ( n1769 ) ;
assign n1771 =  ( n1448 ) ? ( iram_93 ) : ( n1770 ) ;
assign n1772 =  ( n1447 ) ? ( iram_92 ) : ( n1771 ) ;
assign n1773 =  ( n1446 ) ? ( iram_91 ) : ( n1772 ) ;
assign n1774 =  ( n1445 ) ? ( iram_90 ) : ( n1773 ) ;
assign n1775 =  ( n1444 ) ? ( iram_89 ) : ( n1774 ) ;
assign n1776 =  ( n1443 ) ? ( iram_88 ) : ( n1775 ) ;
assign n1777 =  ( n1442 ) ? ( iram_87 ) : ( n1776 ) ;
assign n1778 =  ( n1441 ) ? ( iram_86 ) : ( n1777 ) ;
assign n1779 =  ( n1440 ) ? ( iram_85 ) : ( n1778 ) ;
assign n1780 =  ( n1439 ) ? ( iram_84 ) : ( n1779 ) ;
assign n1781 =  ( n1438 ) ? ( iram_83 ) : ( n1780 ) ;
assign n1782 =  ( n1437 ) ? ( iram_82 ) : ( n1781 ) ;
assign n1783 =  ( n1436 ) ? ( iram_81 ) : ( n1782 ) ;
assign n1784 =  ( n1435 ) ? ( iram_80 ) : ( n1783 ) ;
assign n1785 =  ( n1434 ) ? ( iram_79 ) : ( n1784 ) ;
assign n1786 =  ( n1433 ) ? ( iram_78 ) : ( n1785 ) ;
assign n1787 =  ( n1432 ) ? ( iram_77 ) : ( n1786 ) ;
assign n1788 =  ( n1431 ) ? ( iram_76 ) : ( n1787 ) ;
assign n1789 =  ( n1430 ) ? ( iram_75 ) : ( n1788 ) ;
assign n1790 =  ( n1429 ) ? ( iram_74 ) : ( n1789 ) ;
assign n1791 =  ( n1428 ) ? ( iram_73 ) : ( n1790 ) ;
assign n1792 =  ( n1427 ) ? ( iram_72 ) : ( n1791 ) ;
assign n1793 =  ( n1426 ) ? ( iram_71 ) : ( n1792 ) ;
assign n1794 =  ( n1425 ) ? ( iram_70 ) : ( n1793 ) ;
assign n1795 =  ( n1424 ) ? ( iram_69 ) : ( n1794 ) ;
assign n1796 =  ( n1423 ) ? ( iram_68 ) : ( n1795 ) ;
assign n1797 =  ( n1422 ) ? ( iram_67 ) : ( n1796 ) ;
assign n1798 =  ( n1421 ) ? ( iram_66 ) : ( n1797 ) ;
assign n1799 =  ( n1420 ) ? ( iram_65 ) : ( n1798 ) ;
assign n1800 =  ( n1419 ) ? ( iram_64 ) : ( n1799 ) ;
assign n1801 =  ( n1418 ) ? ( iram_63 ) : ( n1800 ) ;
assign n1802 =  ( n1417 ) ? ( iram_62 ) : ( n1801 ) ;
assign n1803 =  ( n1416 ) ? ( iram_61 ) : ( n1802 ) ;
assign n1804 =  ( n1415 ) ? ( iram_60 ) : ( n1803 ) ;
assign n1805 =  ( n1414 ) ? ( iram_59 ) : ( n1804 ) ;
assign n1806 =  ( n1413 ) ? ( iram_58 ) : ( n1805 ) ;
assign n1807 =  ( n1412 ) ? ( iram_57 ) : ( n1806 ) ;
assign n1808 =  ( n1411 ) ? ( iram_56 ) : ( n1807 ) ;
assign n1809 =  ( n1410 ) ? ( iram_55 ) : ( n1808 ) ;
assign n1810 =  ( n1409 ) ? ( iram_54 ) : ( n1809 ) ;
assign n1811 =  ( n1408 ) ? ( iram_53 ) : ( n1810 ) ;
assign n1812 =  ( n1407 ) ? ( iram_52 ) : ( n1811 ) ;
assign n1813 =  ( n1406 ) ? ( iram_51 ) : ( n1812 ) ;
assign n1814 =  ( n1405 ) ? ( iram_50 ) : ( n1813 ) ;
assign n1815 =  ( n1404 ) ? ( iram_49 ) : ( n1814 ) ;
assign n1816 =  ( n1403 ) ? ( iram_48 ) : ( n1815 ) ;
assign n1817 =  ( n1402 ) ? ( iram_47 ) : ( n1816 ) ;
assign n1818 =  ( n1401 ) ? ( iram_46 ) : ( n1817 ) ;
assign n1819 =  ( n1400 ) ? ( iram_45 ) : ( n1818 ) ;
assign n1820 =  ( n1399 ) ? ( iram_44 ) : ( n1819 ) ;
assign n1821 =  ( n1398 ) ? ( iram_43 ) : ( n1820 ) ;
assign n1822 =  ( n1397 ) ? ( iram_42 ) : ( n1821 ) ;
assign n1823 =  ( n1396 ) ? ( iram_41 ) : ( n1822 ) ;
assign n1824 =  ( n1395 ) ? ( iram_40 ) : ( n1823 ) ;
assign n1825 =  ( n1394 ) ? ( iram_39 ) : ( n1824 ) ;
assign n1826 =  ( n1393 ) ? ( iram_38 ) : ( n1825 ) ;
assign n1827 =  ( n1392 ) ? ( iram_37 ) : ( n1826 ) ;
assign n1828 =  ( n1391 ) ? ( iram_36 ) : ( n1827 ) ;
assign n1829 =  ( n1390 ) ? ( iram_35 ) : ( n1828 ) ;
assign n1830 =  ( n1389 ) ? ( iram_34 ) : ( n1829 ) ;
assign n1831 =  ( n1388 ) ? ( iram_33 ) : ( n1830 ) ;
assign n1832 =  ( n1387 ) ? ( iram_32 ) : ( n1831 ) ;
assign n1833 =  ( n1386 ) ? ( iram_31 ) : ( n1832 ) ;
assign n1834 =  ( n1385 ) ? ( iram_30 ) : ( n1833 ) ;
assign n1835 =  ( n1384 ) ? ( iram_29 ) : ( n1834 ) ;
assign n1836 =  ( n1383 ) ? ( iram_28 ) : ( n1835 ) ;
assign n1837 =  ( n1382 ) ? ( iram_27 ) : ( n1836 ) ;
assign n1838 =  ( n1381 ) ? ( iram_26 ) : ( n1837 ) ;
assign n1839 =  ( n1380 ) ? ( iram_25 ) : ( n1838 ) ;
assign n1840 =  ( n1379 ) ? ( iram_24 ) : ( n1839 ) ;
assign n1841 =  ( n1378 ) ? ( iram_23 ) : ( n1840 ) ;
assign n1842 =  ( n1377 ) ? ( iram_22 ) : ( n1841 ) ;
assign n1843 =  ( n1376 ) ? ( iram_21 ) : ( n1842 ) ;
assign n1844 =  ( n1375 ) ? ( iram_20 ) : ( n1843 ) ;
assign n1845 =  ( n1374 ) ? ( iram_19 ) : ( n1844 ) ;
assign n1846 =  ( n1373 ) ? ( iram_18 ) : ( n1845 ) ;
assign n1847 =  ( n1372 ) ? ( iram_17 ) : ( n1846 ) ;
assign n1848 =  ( n1371 ) ? ( iram_16 ) : ( n1847 ) ;
assign n1849 =  ( n1370 ) ? ( iram_15 ) : ( n1848 ) ;
assign n1850 =  ( n1369 ) ? ( iram_14 ) : ( n1849 ) ;
assign n1851 =  ( n1368 ) ? ( iram_13 ) : ( n1850 ) ;
assign n1852 =  ( n1367 ) ? ( iram_12 ) : ( n1851 ) ;
assign n1853 =  ( n1366 ) ? ( iram_11 ) : ( n1852 ) ;
assign n1854 =  ( n1365 ) ? ( iram_10 ) : ( n1853 ) ;
assign n1855 =  ( n1364 ) ? ( iram_9 ) : ( n1854 ) ;
assign n1856 =  ( n1363 ) ? ( iram_8 ) : ( n1855 ) ;
assign n1857 =  ( n1362 ) ? ( iram_7 ) : ( n1856 ) ;
assign n1858 =  ( n1361 ) ? ( iram_6 ) : ( n1857 ) ;
assign n1859 =  ( n1360 ) ? ( iram_5 ) : ( n1858 ) ;
assign n1860 =  ( n1359 ) ? ( iram_4 ) : ( n1859 ) ;
assign n1861 =  ( n1358 ) ? ( iram_3 ) : ( n1860 ) ;
assign n1862 =  ( n1357 ) ? ( iram_2 ) : ( n1861 ) ;
assign n1863 =  ( n1356 ) ? ( iram_1 ) : ( n1862 ) ;
assign n1864 =  ( n1355 ) ? ( iram_0 ) : ( n1863 ) ;
assign n1865 = rd_addr[7:7] ;
assign n1866 =  ( n1865 ) == ( bv_1_1_n34 )  ;
assign n1867 = rd_addr[6:3] ;
assign n1868 =  { ( bv_1_1_n34 ) , ( n1867 ) }  ;
assign n1869 =  { ( n1868 ) , ( bv_3_0_n46 ) }  ;
assign n1870 = rd_addr[6:3] ;
assign n1871 =  { ( bv_4_2_n12 ) , ( n1870 ) }  ;
assign n1872 =  ( n1866 ) ? ( n1869 ) : ( n1871 ) ;
assign n1873 =  ( bit_addr ) ? ( n1872 ) : ( rd_addr ) ;
assign n1874 = n1873[7:0] ;
assign n1875 =  ( n1874 ) == ( bv_8_0_n69 )  ;
assign n1876 =  ( n1874 ) == ( bv_8_1_n71 )  ;
assign n1877 =  ( n1874 ) == ( bv_8_2_n73 )  ;
assign n1878 =  ( n1874 ) == ( bv_8_3_n75 )  ;
assign n1879 =  ( n1874 ) == ( bv_8_4_n77 )  ;
assign n1880 =  ( n1874 ) == ( bv_8_5_n79 )  ;
assign n1881 =  ( n1874 ) == ( bv_8_6_n81 )  ;
assign n1882 =  ( n1874 ) == ( bv_8_7_n83 )  ;
assign n1883 =  ( n1874 ) == ( bv_8_8_n85 )  ;
assign n1884 =  ( n1874 ) == ( bv_8_9_n87 )  ;
assign n1885 =  ( n1874 ) == ( bv_8_10_n89 )  ;
assign n1886 =  ( n1874 ) == ( bv_8_11_n91 )  ;
assign n1887 =  ( n1874 ) == ( bv_8_12_n93 )  ;
assign n1888 =  ( n1874 ) == ( bv_8_13_n95 )  ;
assign n1889 =  ( n1874 ) == ( bv_8_14_n97 )  ;
assign n1890 =  ( n1874 ) == ( bv_8_15_n99 )  ;
assign n1891 =  ( n1874 ) == ( bv_8_16_n101 )  ;
assign n1892 =  ( n1874 ) == ( bv_8_17_n103 )  ;
assign n1893 =  ( n1874 ) == ( bv_8_18_n105 )  ;
assign n1894 =  ( n1874 ) == ( bv_8_19_n107 )  ;
assign n1895 =  ( n1874 ) == ( bv_8_20_n109 )  ;
assign n1896 =  ( n1874 ) == ( bv_8_21_n111 )  ;
assign n1897 =  ( n1874 ) == ( bv_8_22_n113 )  ;
assign n1898 =  ( n1874 ) == ( bv_8_23_n115 )  ;
assign n1899 =  ( n1874 ) == ( bv_8_24_n117 )  ;
assign n1900 =  ( n1874 ) == ( bv_8_25_n119 )  ;
assign n1901 =  ( n1874 ) == ( bv_8_26_n121 )  ;
assign n1902 =  ( n1874 ) == ( bv_8_27_n123 )  ;
assign n1903 =  ( n1874 ) == ( bv_8_28_n125 )  ;
assign n1904 =  ( n1874 ) == ( bv_8_29_n127 )  ;
assign n1905 =  ( n1874 ) == ( bv_8_30_n129 )  ;
assign n1906 =  ( n1874 ) == ( bv_8_31_n131 )  ;
assign n1907 =  ( n1874 ) == ( bv_8_32_n133 )  ;
assign n1908 =  ( n1874 ) == ( bv_8_33_n135 )  ;
assign n1909 =  ( n1874 ) == ( bv_8_34_n137 )  ;
assign n1910 =  ( n1874 ) == ( bv_8_35_n139 )  ;
assign n1911 =  ( n1874 ) == ( bv_8_36_n141 )  ;
assign n1912 =  ( n1874 ) == ( bv_8_37_n143 )  ;
assign n1913 =  ( n1874 ) == ( bv_8_38_n145 )  ;
assign n1914 =  ( n1874 ) == ( bv_8_39_n147 )  ;
assign n1915 =  ( n1874 ) == ( bv_8_40_n149 )  ;
assign n1916 =  ( n1874 ) == ( bv_8_41_n151 )  ;
assign n1917 =  ( n1874 ) == ( bv_8_42_n153 )  ;
assign n1918 =  ( n1874 ) == ( bv_8_43_n155 )  ;
assign n1919 =  ( n1874 ) == ( bv_8_44_n157 )  ;
assign n1920 =  ( n1874 ) == ( bv_8_45_n159 )  ;
assign n1921 =  ( n1874 ) == ( bv_8_46_n161 )  ;
assign n1922 =  ( n1874 ) == ( bv_8_47_n163 )  ;
assign n1923 =  ( n1874 ) == ( bv_8_48_n165 )  ;
assign n1924 =  ( n1874 ) == ( bv_8_49_n167 )  ;
assign n1925 =  ( n1874 ) == ( bv_8_50_n169 )  ;
assign n1926 =  ( n1874 ) == ( bv_8_51_n171 )  ;
assign n1927 =  ( n1874 ) == ( bv_8_52_n173 )  ;
assign n1928 =  ( n1874 ) == ( bv_8_53_n175 )  ;
assign n1929 =  ( n1874 ) == ( bv_8_54_n177 )  ;
assign n1930 =  ( n1874 ) == ( bv_8_55_n179 )  ;
assign n1931 =  ( n1874 ) == ( bv_8_56_n181 )  ;
assign n1932 =  ( n1874 ) == ( bv_8_57_n183 )  ;
assign n1933 =  ( n1874 ) == ( bv_8_58_n185 )  ;
assign n1934 =  ( n1874 ) == ( bv_8_59_n187 )  ;
assign n1935 =  ( n1874 ) == ( bv_8_60_n189 )  ;
assign n1936 =  ( n1874 ) == ( bv_8_61_n191 )  ;
assign n1937 =  ( n1874 ) == ( bv_8_62_n193 )  ;
assign n1938 =  ( n1874 ) == ( bv_8_63_n195 )  ;
assign n1939 =  ( n1874 ) == ( bv_8_64_n197 )  ;
assign n1940 =  ( n1874 ) == ( bv_8_65_n199 )  ;
assign n1941 =  ( n1874 ) == ( bv_8_66_n201 )  ;
assign n1942 =  ( n1874 ) == ( bv_8_67_n203 )  ;
assign n1943 =  ( n1874 ) == ( bv_8_68_n205 )  ;
assign n1944 =  ( n1874 ) == ( bv_8_69_n207 )  ;
assign n1945 =  ( n1874 ) == ( bv_8_70_n209 )  ;
assign n1946 =  ( n1874 ) == ( bv_8_71_n211 )  ;
assign n1947 =  ( n1874 ) == ( bv_8_72_n213 )  ;
assign n1948 =  ( n1874 ) == ( bv_8_73_n215 )  ;
assign n1949 =  ( n1874 ) == ( bv_8_74_n217 )  ;
assign n1950 =  ( n1874 ) == ( bv_8_75_n219 )  ;
assign n1951 =  ( n1874 ) == ( bv_8_76_n221 )  ;
assign n1952 =  ( n1874 ) == ( bv_8_77_n223 )  ;
assign n1953 =  ( n1874 ) == ( bv_8_78_n225 )  ;
assign n1954 =  ( n1874 ) == ( bv_8_79_n227 )  ;
assign n1955 =  ( n1874 ) == ( bv_8_80_n229 )  ;
assign n1956 =  ( n1874 ) == ( bv_8_81_n231 )  ;
assign n1957 =  ( n1874 ) == ( bv_8_82_n233 )  ;
assign n1958 =  ( n1874 ) == ( bv_8_83_n235 )  ;
assign n1959 =  ( n1874 ) == ( bv_8_84_n237 )  ;
assign n1960 =  ( n1874 ) == ( bv_8_85_n239 )  ;
assign n1961 =  ( n1874 ) == ( bv_8_86_n241 )  ;
assign n1962 =  ( n1874 ) == ( bv_8_87_n243 )  ;
assign n1963 =  ( n1874 ) == ( bv_8_88_n245 )  ;
assign n1964 =  ( n1874 ) == ( bv_8_89_n247 )  ;
assign n1965 =  ( n1874 ) == ( bv_8_90_n249 )  ;
assign n1966 =  ( n1874 ) == ( bv_8_91_n251 )  ;
assign n1967 =  ( n1874 ) == ( bv_8_92_n253 )  ;
assign n1968 =  ( n1874 ) == ( bv_8_93_n255 )  ;
assign n1969 =  ( n1874 ) == ( bv_8_94_n257 )  ;
assign n1970 =  ( n1874 ) == ( bv_8_95_n259 )  ;
assign n1971 =  ( n1874 ) == ( bv_8_96_n261 )  ;
assign n1972 =  ( n1874 ) == ( bv_8_97_n263 )  ;
assign n1973 =  ( n1874 ) == ( bv_8_98_n265 )  ;
assign n1974 =  ( n1874 ) == ( bv_8_99_n267 )  ;
assign n1975 =  ( n1874 ) == ( bv_8_100_n269 )  ;
assign n1976 =  ( n1874 ) == ( bv_8_101_n271 )  ;
assign n1977 =  ( n1874 ) == ( bv_8_102_n273 )  ;
assign n1978 =  ( n1874 ) == ( bv_8_103_n275 )  ;
assign n1979 =  ( n1874 ) == ( bv_8_104_n277 )  ;
assign n1980 =  ( n1874 ) == ( bv_8_105_n279 )  ;
assign n1981 =  ( n1874 ) == ( bv_8_106_n281 )  ;
assign n1982 =  ( n1874 ) == ( bv_8_107_n283 )  ;
assign n1983 =  ( n1874 ) == ( bv_8_108_n285 )  ;
assign n1984 =  ( n1874 ) == ( bv_8_109_n287 )  ;
assign n1985 =  ( n1874 ) == ( bv_8_110_n289 )  ;
assign n1986 =  ( n1874 ) == ( bv_8_111_n291 )  ;
assign n1987 =  ( n1874 ) == ( bv_8_112_n293 )  ;
assign n1988 =  ( n1874 ) == ( bv_8_113_n295 )  ;
assign n1989 =  ( n1874 ) == ( bv_8_114_n297 )  ;
assign n1990 =  ( n1874 ) == ( bv_8_115_n299 )  ;
assign n1991 =  ( n1874 ) == ( bv_8_116_n301 )  ;
assign n1992 =  ( n1874 ) == ( bv_8_117_n303 )  ;
assign n1993 =  ( n1874 ) == ( bv_8_118_n305 )  ;
assign n1994 =  ( n1874 ) == ( bv_8_119_n307 )  ;
assign n1995 =  ( n1874 ) == ( bv_8_120_n309 )  ;
assign n1996 =  ( n1874 ) == ( bv_8_121_n311 )  ;
assign n1997 =  ( n1874 ) == ( bv_8_122_n313 )  ;
assign n1998 =  ( n1874 ) == ( bv_8_123_n315 )  ;
assign n1999 =  ( n1874 ) == ( bv_8_124_n317 )  ;
assign n2000 =  ( n1874 ) == ( bv_8_125_n319 )  ;
assign n2001 =  ( n1874 ) == ( bv_8_126_n321 )  ;
assign n2002 =  ( n1874 ) == ( bv_8_127_n323 )  ;
assign n2003 =  ( n1874 ) == ( bv_8_128_n325 )  ;
assign n2004 =  ( n1874 ) == ( bv_8_129_n327 )  ;
assign n2005 =  ( n1874 ) == ( bv_8_130_n329 )  ;
assign n2006 =  ( n1874 ) == ( bv_8_131_n331 )  ;
assign n2007 =  ( n1874 ) == ( bv_8_132_n333 )  ;
assign n2008 =  ( n1874 ) == ( bv_8_133_n335 )  ;
assign n2009 =  ( n1874 ) == ( bv_8_134_n337 )  ;
assign n2010 =  ( n1874 ) == ( bv_8_135_n339 )  ;
assign n2011 =  ( n1874 ) == ( bv_8_136_n341 )  ;
assign n2012 =  ( n1874 ) == ( bv_8_137_n343 )  ;
assign n2013 =  ( n1874 ) == ( bv_8_138_n345 )  ;
assign n2014 =  ( n1874 ) == ( bv_8_139_n347 )  ;
assign n2015 =  ( n1874 ) == ( bv_8_140_n349 )  ;
assign n2016 =  ( n1874 ) == ( bv_8_141_n351 )  ;
assign n2017 =  ( n1874 ) == ( bv_8_142_n353 )  ;
assign n2018 =  ( n1874 ) == ( bv_8_143_n355 )  ;
assign n2019 =  ( n1874 ) == ( bv_8_144_n357 )  ;
assign n2020 =  ( n1874 ) == ( bv_8_145_n359 )  ;
assign n2021 =  ( n1874 ) == ( bv_8_146_n361 )  ;
assign n2022 =  ( n1874 ) == ( bv_8_147_n363 )  ;
assign n2023 =  ( n1874 ) == ( bv_8_148_n365 )  ;
assign n2024 =  ( n1874 ) == ( bv_8_149_n367 )  ;
assign n2025 =  ( n1874 ) == ( bv_8_150_n369 )  ;
assign n2026 =  ( n1874 ) == ( bv_8_151_n371 )  ;
assign n2027 =  ( n1874 ) == ( bv_8_152_n373 )  ;
assign n2028 =  ( n1874 ) == ( bv_8_153_n375 )  ;
assign n2029 =  ( n1874 ) == ( bv_8_154_n377 )  ;
assign n2030 =  ( n1874 ) == ( bv_8_155_n379 )  ;
assign n2031 =  ( n1874 ) == ( bv_8_156_n381 )  ;
assign n2032 =  ( n1874 ) == ( bv_8_157_n383 )  ;
assign n2033 =  ( n1874 ) == ( bv_8_158_n385 )  ;
assign n2034 =  ( n1874 ) == ( bv_8_159_n387 )  ;
assign n2035 =  ( n1874 ) == ( bv_8_160_n389 )  ;
assign n2036 =  ( n1874 ) == ( bv_8_161_n391 )  ;
assign n2037 =  ( n1874 ) == ( bv_8_162_n393 )  ;
assign n2038 =  ( n1874 ) == ( bv_8_163_n395 )  ;
assign n2039 =  ( n1874 ) == ( bv_8_164_n397 )  ;
assign n2040 =  ( n1874 ) == ( bv_8_165_n399 )  ;
assign n2041 =  ( n1874 ) == ( bv_8_166_n401 )  ;
assign n2042 =  ( n1874 ) == ( bv_8_167_n403 )  ;
assign n2043 =  ( n1874 ) == ( bv_8_168_n405 )  ;
assign n2044 =  ( n1874 ) == ( bv_8_169_n407 )  ;
assign n2045 =  ( n1874 ) == ( bv_8_170_n409 )  ;
assign n2046 =  ( n1874 ) == ( bv_8_171_n411 )  ;
assign n2047 =  ( n1874 ) == ( bv_8_172_n413 )  ;
assign n2048 =  ( n1874 ) == ( bv_8_173_n415 )  ;
assign n2049 =  ( n1874 ) == ( bv_8_174_n417 )  ;
assign n2050 =  ( n1874 ) == ( bv_8_175_n419 )  ;
assign n2051 =  ( n1874 ) == ( bv_8_176_n421 )  ;
assign n2052 =  ( n1874 ) == ( bv_8_177_n423 )  ;
assign n2053 =  ( n1874 ) == ( bv_8_178_n425 )  ;
assign n2054 =  ( n1874 ) == ( bv_8_179_n427 )  ;
assign n2055 =  ( n1874 ) == ( bv_8_180_n429 )  ;
assign n2056 =  ( n1874 ) == ( bv_8_181_n431 )  ;
assign n2057 =  ( n1874 ) == ( bv_8_182_n433 )  ;
assign n2058 =  ( n1874 ) == ( bv_8_183_n435 )  ;
assign n2059 =  ( n1874 ) == ( bv_8_184_n437 )  ;
assign n2060 =  ( n1874 ) == ( bv_8_185_n439 )  ;
assign n2061 =  ( n1874 ) == ( bv_8_186_n441 )  ;
assign n2062 =  ( n1874 ) == ( bv_8_187_n443 )  ;
assign n2063 =  ( n1874 ) == ( bv_8_188_n445 )  ;
assign n2064 =  ( n1874 ) == ( bv_8_189_n447 )  ;
assign n2065 =  ( n1874 ) == ( bv_8_190_n449 )  ;
assign n2066 =  ( n1874 ) == ( bv_8_191_n451 )  ;
assign n2067 =  ( n1874 ) == ( bv_8_192_n453 )  ;
assign n2068 =  ( n1874 ) == ( bv_8_193_n455 )  ;
assign n2069 =  ( n1874 ) == ( bv_8_194_n457 )  ;
assign n2070 =  ( n1874 ) == ( bv_8_195_n459 )  ;
assign n2071 =  ( n1874 ) == ( bv_8_196_n461 )  ;
assign n2072 =  ( n1874 ) == ( bv_8_197_n463 )  ;
assign n2073 =  ( n1874 ) == ( bv_8_198_n465 )  ;
assign n2074 =  ( n1874 ) == ( bv_8_199_n467 )  ;
assign n2075 =  ( n1874 ) == ( bv_8_200_n469 )  ;
assign n2076 =  ( n1874 ) == ( bv_8_201_n471 )  ;
assign n2077 =  ( n1874 ) == ( bv_8_202_n473 )  ;
assign n2078 =  ( n1874 ) == ( bv_8_203_n475 )  ;
assign n2079 =  ( n1874 ) == ( bv_8_204_n477 )  ;
assign n2080 =  ( n1874 ) == ( bv_8_205_n479 )  ;
assign n2081 =  ( n1874 ) == ( bv_8_206_n481 )  ;
assign n2082 =  ( n1874 ) == ( bv_8_207_n483 )  ;
assign n2083 =  ( n1874 ) == ( bv_8_208_n485 )  ;
assign n2084 =  ( n1874 ) == ( bv_8_209_n487 )  ;
assign n2085 =  ( n1874 ) == ( bv_8_210_n489 )  ;
assign n2086 =  ( n1874 ) == ( bv_8_211_n491 )  ;
assign n2087 =  ( n1874 ) == ( bv_8_212_n493 )  ;
assign n2088 =  ( n1874 ) == ( bv_8_213_n495 )  ;
assign n2089 =  ( n1874 ) == ( bv_8_214_n497 )  ;
assign n2090 =  ( n1874 ) == ( bv_8_215_n499 )  ;
assign n2091 =  ( n1874 ) == ( bv_8_216_n501 )  ;
assign n2092 =  ( n1874 ) == ( bv_8_217_n503 )  ;
assign n2093 =  ( n1874 ) == ( bv_8_218_n505 )  ;
assign n2094 =  ( n1874 ) == ( bv_8_219_n507 )  ;
assign n2095 =  ( n1874 ) == ( bv_8_220_n509 )  ;
assign n2096 =  ( n1874 ) == ( bv_8_221_n511 )  ;
assign n2097 =  ( n1874 ) == ( bv_8_222_n513 )  ;
assign n2098 =  ( n1874 ) == ( bv_8_223_n515 )  ;
assign n2099 =  ( n1874 ) == ( bv_8_224_n517 )  ;
assign n2100 =  ( n1874 ) == ( bv_8_225_n519 )  ;
assign n2101 =  ( n1874 ) == ( bv_8_226_n521 )  ;
assign n2102 =  ( n1874 ) == ( bv_8_227_n523 )  ;
assign n2103 =  ( n1874 ) == ( bv_8_228_n525 )  ;
assign n2104 =  ( n1874 ) == ( bv_8_229_n527 )  ;
assign n2105 =  ( n1874 ) == ( bv_8_230_n529 )  ;
assign n2106 =  ( n1874 ) == ( bv_8_231_n531 )  ;
assign n2107 =  ( n1874 ) == ( bv_8_232_n533 )  ;
assign n2108 =  ( n1874 ) == ( bv_8_233_n535 )  ;
assign n2109 =  ( n1874 ) == ( bv_8_234_n537 )  ;
assign n2110 =  ( n1874 ) == ( bv_8_235_n539 )  ;
assign n2111 =  ( n1874 ) == ( bv_8_236_n541 )  ;
assign n2112 =  ( n1874 ) == ( bv_8_237_n543 )  ;
assign n2113 =  ( n1874 ) == ( bv_8_238_n545 )  ;
assign n2114 =  ( n1874 ) == ( bv_8_239_n547 )  ;
assign n2115 =  ( n1874 ) == ( bv_8_240_n549 )  ;
assign n2116 =  ( n1874 ) == ( bv_8_241_n551 )  ;
assign n2117 =  ( n1874 ) == ( bv_8_242_n553 )  ;
assign n2118 =  ( n1874 ) == ( bv_8_243_n555 )  ;
assign n2119 =  ( n1874 ) == ( bv_8_244_n557 )  ;
assign n2120 =  ( n1874 ) == ( bv_8_245_n559 )  ;
assign n2121 =  ( n1874 ) == ( bv_8_246_n561 )  ;
assign n2122 =  ( n1874 ) == ( bv_8_247_n563 )  ;
assign n2123 =  ( n1874 ) == ( bv_8_248_n565 )  ;
assign n2124 =  ( n1874 ) == ( bv_8_249_n567 )  ;
assign n2125 =  ( n1874 ) == ( bv_8_250_n569 )  ;
assign n2126 =  ( n1874 ) == ( bv_8_251_n571 )  ;
assign n2127 =  ( n1874 ) == ( bv_8_252_n573 )  ;
assign n2128 =  ( n1874 ) == ( bv_8_253_n575 )  ;
assign n2129 =  ( n1874 ) == ( bv_8_254_n577 )  ;
assign n2130 =  ( n2129 ) ? ( iram_254 ) : ( iram_255 ) ;
assign n2131 =  ( n2128 ) ? ( iram_253 ) : ( n2130 ) ;
assign n2132 =  ( n2127 ) ? ( iram_252 ) : ( n2131 ) ;
assign n2133 =  ( n2126 ) ? ( iram_251 ) : ( n2132 ) ;
assign n2134 =  ( n2125 ) ? ( iram_250 ) : ( n2133 ) ;
assign n2135 =  ( n2124 ) ? ( iram_249 ) : ( n2134 ) ;
assign n2136 =  ( n2123 ) ? ( iram_248 ) : ( n2135 ) ;
assign n2137 =  ( n2122 ) ? ( iram_247 ) : ( n2136 ) ;
assign n2138 =  ( n2121 ) ? ( iram_246 ) : ( n2137 ) ;
assign n2139 =  ( n2120 ) ? ( iram_245 ) : ( n2138 ) ;
assign n2140 =  ( n2119 ) ? ( iram_244 ) : ( n2139 ) ;
assign n2141 =  ( n2118 ) ? ( iram_243 ) : ( n2140 ) ;
assign n2142 =  ( n2117 ) ? ( iram_242 ) : ( n2141 ) ;
assign n2143 =  ( n2116 ) ? ( iram_241 ) : ( n2142 ) ;
assign n2144 =  ( n2115 ) ? ( iram_240 ) : ( n2143 ) ;
assign n2145 =  ( n2114 ) ? ( iram_239 ) : ( n2144 ) ;
assign n2146 =  ( n2113 ) ? ( iram_238 ) : ( n2145 ) ;
assign n2147 =  ( n2112 ) ? ( iram_237 ) : ( n2146 ) ;
assign n2148 =  ( n2111 ) ? ( iram_236 ) : ( n2147 ) ;
assign n2149 =  ( n2110 ) ? ( iram_235 ) : ( n2148 ) ;
assign n2150 =  ( n2109 ) ? ( iram_234 ) : ( n2149 ) ;
assign n2151 =  ( n2108 ) ? ( iram_233 ) : ( n2150 ) ;
assign n2152 =  ( n2107 ) ? ( iram_232 ) : ( n2151 ) ;
assign n2153 =  ( n2106 ) ? ( iram_231 ) : ( n2152 ) ;
assign n2154 =  ( n2105 ) ? ( iram_230 ) : ( n2153 ) ;
assign n2155 =  ( n2104 ) ? ( iram_229 ) : ( n2154 ) ;
assign n2156 =  ( n2103 ) ? ( iram_228 ) : ( n2155 ) ;
assign n2157 =  ( n2102 ) ? ( iram_227 ) : ( n2156 ) ;
assign n2158 =  ( n2101 ) ? ( iram_226 ) : ( n2157 ) ;
assign n2159 =  ( n2100 ) ? ( iram_225 ) : ( n2158 ) ;
assign n2160 =  ( n2099 ) ? ( iram_224 ) : ( n2159 ) ;
assign n2161 =  ( n2098 ) ? ( iram_223 ) : ( n2160 ) ;
assign n2162 =  ( n2097 ) ? ( iram_222 ) : ( n2161 ) ;
assign n2163 =  ( n2096 ) ? ( iram_221 ) : ( n2162 ) ;
assign n2164 =  ( n2095 ) ? ( iram_220 ) : ( n2163 ) ;
assign n2165 =  ( n2094 ) ? ( iram_219 ) : ( n2164 ) ;
assign n2166 =  ( n2093 ) ? ( iram_218 ) : ( n2165 ) ;
assign n2167 =  ( n2092 ) ? ( iram_217 ) : ( n2166 ) ;
assign n2168 =  ( n2091 ) ? ( iram_216 ) : ( n2167 ) ;
assign n2169 =  ( n2090 ) ? ( iram_215 ) : ( n2168 ) ;
assign n2170 =  ( n2089 ) ? ( iram_214 ) : ( n2169 ) ;
assign n2171 =  ( n2088 ) ? ( iram_213 ) : ( n2170 ) ;
assign n2172 =  ( n2087 ) ? ( iram_212 ) : ( n2171 ) ;
assign n2173 =  ( n2086 ) ? ( iram_211 ) : ( n2172 ) ;
assign n2174 =  ( n2085 ) ? ( iram_210 ) : ( n2173 ) ;
assign n2175 =  ( n2084 ) ? ( iram_209 ) : ( n2174 ) ;
assign n2176 =  ( n2083 ) ? ( iram_208 ) : ( n2175 ) ;
assign n2177 =  ( n2082 ) ? ( iram_207 ) : ( n2176 ) ;
assign n2178 =  ( n2081 ) ? ( iram_206 ) : ( n2177 ) ;
assign n2179 =  ( n2080 ) ? ( iram_205 ) : ( n2178 ) ;
assign n2180 =  ( n2079 ) ? ( iram_204 ) : ( n2179 ) ;
assign n2181 =  ( n2078 ) ? ( iram_203 ) : ( n2180 ) ;
assign n2182 =  ( n2077 ) ? ( iram_202 ) : ( n2181 ) ;
assign n2183 =  ( n2076 ) ? ( iram_201 ) : ( n2182 ) ;
assign n2184 =  ( n2075 ) ? ( iram_200 ) : ( n2183 ) ;
assign n2185 =  ( n2074 ) ? ( iram_199 ) : ( n2184 ) ;
assign n2186 =  ( n2073 ) ? ( iram_198 ) : ( n2185 ) ;
assign n2187 =  ( n2072 ) ? ( iram_197 ) : ( n2186 ) ;
assign n2188 =  ( n2071 ) ? ( iram_196 ) : ( n2187 ) ;
assign n2189 =  ( n2070 ) ? ( iram_195 ) : ( n2188 ) ;
assign n2190 =  ( n2069 ) ? ( iram_194 ) : ( n2189 ) ;
assign n2191 =  ( n2068 ) ? ( iram_193 ) : ( n2190 ) ;
assign n2192 =  ( n2067 ) ? ( iram_192 ) : ( n2191 ) ;
assign n2193 =  ( n2066 ) ? ( iram_191 ) : ( n2192 ) ;
assign n2194 =  ( n2065 ) ? ( iram_190 ) : ( n2193 ) ;
assign n2195 =  ( n2064 ) ? ( iram_189 ) : ( n2194 ) ;
assign n2196 =  ( n2063 ) ? ( iram_188 ) : ( n2195 ) ;
assign n2197 =  ( n2062 ) ? ( iram_187 ) : ( n2196 ) ;
assign n2198 =  ( n2061 ) ? ( iram_186 ) : ( n2197 ) ;
assign n2199 =  ( n2060 ) ? ( iram_185 ) : ( n2198 ) ;
assign n2200 =  ( n2059 ) ? ( iram_184 ) : ( n2199 ) ;
assign n2201 =  ( n2058 ) ? ( iram_183 ) : ( n2200 ) ;
assign n2202 =  ( n2057 ) ? ( iram_182 ) : ( n2201 ) ;
assign n2203 =  ( n2056 ) ? ( iram_181 ) : ( n2202 ) ;
assign n2204 =  ( n2055 ) ? ( iram_180 ) : ( n2203 ) ;
assign n2205 =  ( n2054 ) ? ( iram_179 ) : ( n2204 ) ;
assign n2206 =  ( n2053 ) ? ( iram_178 ) : ( n2205 ) ;
assign n2207 =  ( n2052 ) ? ( iram_177 ) : ( n2206 ) ;
assign n2208 =  ( n2051 ) ? ( iram_176 ) : ( n2207 ) ;
assign n2209 =  ( n2050 ) ? ( iram_175 ) : ( n2208 ) ;
assign n2210 =  ( n2049 ) ? ( iram_174 ) : ( n2209 ) ;
assign n2211 =  ( n2048 ) ? ( iram_173 ) : ( n2210 ) ;
assign n2212 =  ( n2047 ) ? ( iram_172 ) : ( n2211 ) ;
assign n2213 =  ( n2046 ) ? ( iram_171 ) : ( n2212 ) ;
assign n2214 =  ( n2045 ) ? ( iram_170 ) : ( n2213 ) ;
assign n2215 =  ( n2044 ) ? ( iram_169 ) : ( n2214 ) ;
assign n2216 =  ( n2043 ) ? ( iram_168 ) : ( n2215 ) ;
assign n2217 =  ( n2042 ) ? ( iram_167 ) : ( n2216 ) ;
assign n2218 =  ( n2041 ) ? ( iram_166 ) : ( n2217 ) ;
assign n2219 =  ( n2040 ) ? ( iram_165 ) : ( n2218 ) ;
assign n2220 =  ( n2039 ) ? ( iram_164 ) : ( n2219 ) ;
assign n2221 =  ( n2038 ) ? ( iram_163 ) : ( n2220 ) ;
assign n2222 =  ( n2037 ) ? ( iram_162 ) : ( n2221 ) ;
assign n2223 =  ( n2036 ) ? ( iram_161 ) : ( n2222 ) ;
assign n2224 =  ( n2035 ) ? ( iram_160 ) : ( n2223 ) ;
assign n2225 =  ( n2034 ) ? ( iram_159 ) : ( n2224 ) ;
assign n2226 =  ( n2033 ) ? ( iram_158 ) : ( n2225 ) ;
assign n2227 =  ( n2032 ) ? ( iram_157 ) : ( n2226 ) ;
assign n2228 =  ( n2031 ) ? ( iram_156 ) : ( n2227 ) ;
assign n2229 =  ( n2030 ) ? ( iram_155 ) : ( n2228 ) ;
assign n2230 =  ( n2029 ) ? ( iram_154 ) : ( n2229 ) ;
assign n2231 =  ( n2028 ) ? ( iram_153 ) : ( n2230 ) ;
assign n2232 =  ( n2027 ) ? ( iram_152 ) : ( n2231 ) ;
assign n2233 =  ( n2026 ) ? ( iram_151 ) : ( n2232 ) ;
assign n2234 =  ( n2025 ) ? ( iram_150 ) : ( n2233 ) ;
assign n2235 =  ( n2024 ) ? ( iram_149 ) : ( n2234 ) ;
assign n2236 =  ( n2023 ) ? ( iram_148 ) : ( n2235 ) ;
assign n2237 =  ( n2022 ) ? ( iram_147 ) : ( n2236 ) ;
assign n2238 =  ( n2021 ) ? ( iram_146 ) : ( n2237 ) ;
assign n2239 =  ( n2020 ) ? ( iram_145 ) : ( n2238 ) ;
assign n2240 =  ( n2019 ) ? ( iram_144 ) : ( n2239 ) ;
assign n2241 =  ( n2018 ) ? ( iram_143 ) : ( n2240 ) ;
assign n2242 =  ( n2017 ) ? ( iram_142 ) : ( n2241 ) ;
assign n2243 =  ( n2016 ) ? ( iram_141 ) : ( n2242 ) ;
assign n2244 =  ( n2015 ) ? ( iram_140 ) : ( n2243 ) ;
assign n2245 =  ( n2014 ) ? ( iram_139 ) : ( n2244 ) ;
assign n2246 =  ( n2013 ) ? ( iram_138 ) : ( n2245 ) ;
assign n2247 =  ( n2012 ) ? ( iram_137 ) : ( n2246 ) ;
assign n2248 =  ( n2011 ) ? ( iram_136 ) : ( n2247 ) ;
assign n2249 =  ( n2010 ) ? ( iram_135 ) : ( n2248 ) ;
assign n2250 =  ( n2009 ) ? ( iram_134 ) : ( n2249 ) ;
assign n2251 =  ( n2008 ) ? ( iram_133 ) : ( n2250 ) ;
assign n2252 =  ( n2007 ) ? ( iram_132 ) : ( n2251 ) ;
assign n2253 =  ( n2006 ) ? ( iram_131 ) : ( n2252 ) ;
assign n2254 =  ( n2005 ) ? ( iram_130 ) : ( n2253 ) ;
assign n2255 =  ( n2004 ) ? ( iram_129 ) : ( n2254 ) ;
assign n2256 =  ( n2003 ) ? ( iram_128 ) : ( n2255 ) ;
assign n2257 =  ( n2002 ) ? ( iram_127 ) : ( n2256 ) ;
assign n2258 =  ( n2001 ) ? ( iram_126 ) : ( n2257 ) ;
assign n2259 =  ( n2000 ) ? ( iram_125 ) : ( n2258 ) ;
assign n2260 =  ( n1999 ) ? ( iram_124 ) : ( n2259 ) ;
assign n2261 =  ( n1998 ) ? ( iram_123 ) : ( n2260 ) ;
assign n2262 =  ( n1997 ) ? ( iram_122 ) : ( n2261 ) ;
assign n2263 =  ( n1996 ) ? ( iram_121 ) : ( n2262 ) ;
assign n2264 =  ( n1995 ) ? ( iram_120 ) : ( n2263 ) ;
assign n2265 =  ( n1994 ) ? ( iram_119 ) : ( n2264 ) ;
assign n2266 =  ( n1993 ) ? ( iram_118 ) : ( n2265 ) ;
assign n2267 =  ( n1992 ) ? ( iram_117 ) : ( n2266 ) ;
assign n2268 =  ( n1991 ) ? ( iram_116 ) : ( n2267 ) ;
assign n2269 =  ( n1990 ) ? ( iram_115 ) : ( n2268 ) ;
assign n2270 =  ( n1989 ) ? ( iram_114 ) : ( n2269 ) ;
assign n2271 =  ( n1988 ) ? ( iram_113 ) : ( n2270 ) ;
assign n2272 =  ( n1987 ) ? ( iram_112 ) : ( n2271 ) ;
assign n2273 =  ( n1986 ) ? ( iram_111 ) : ( n2272 ) ;
assign n2274 =  ( n1985 ) ? ( iram_110 ) : ( n2273 ) ;
assign n2275 =  ( n1984 ) ? ( iram_109 ) : ( n2274 ) ;
assign n2276 =  ( n1983 ) ? ( iram_108 ) : ( n2275 ) ;
assign n2277 =  ( n1982 ) ? ( iram_107 ) : ( n2276 ) ;
assign n2278 =  ( n1981 ) ? ( iram_106 ) : ( n2277 ) ;
assign n2279 =  ( n1980 ) ? ( iram_105 ) : ( n2278 ) ;
assign n2280 =  ( n1979 ) ? ( iram_104 ) : ( n2279 ) ;
assign n2281 =  ( n1978 ) ? ( iram_103 ) : ( n2280 ) ;
assign n2282 =  ( n1977 ) ? ( iram_102 ) : ( n2281 ) ;
assign n2283 =  ( n1976 ) ? ( iram_101 ) : ( n2282 ) ;
assign n2284 =  ( n1975 ) ? ( iram_100 ) : ( n2283 ) ;
assign n2285 =  ( n1974 ) ? ( iram_99 ) : ( n2284 ) ;
assign n2286 =  ( n1973 ) ? ( iram_98 ) : ( n2285 ) ;
assign n2287 =  ( n1972 ) ? ( iram_97 ) : ( n2286 ) ;
assign n2288 =  ( n1971 ) ? ( iram_96 ) : ( n2287 ) ;
assign n2289 =  ( n1970 ) ? ( iram_95 ) : ( n2288 ) ;
assign n2290 =  ( n1969 ) ? ( iram_94 ) : ( n2289 ) ;
assign n2291 =  ( n1968 ) ? ( iram_93 ) : ( n2290 ) ;
assign n2292 =  ( n1967 ) ? ( iram_92 ) : ( n2291 ) ;
assign n2293 =  ( n1966 ) ? ( iram_91 ) : ( n2292 ) ;
assign n2294 =  ( n1965 ) ? ( iram_90 ) : ( n2293 ) ;
assign n2295 =  ( n1964 ) ? ( iram_89 ) : ( n2294 ) ;
assign n2296 =  ( n1963 ) ? ( iram_88 ) : ( n2295 ) ;
assign n2297 =  ( n1962 ) ? ( iram_87 ) : ( n2296 ) ;
assign n2298 =  ( n1961 ) ? ( iram_86 ) : ( n2297 ) ;
assign n2299 =  ( n1960 ) ? ( iram_85 ) : ( n2298 ) ;
assign n2300 =  ( n1959 ) ? ( iram_84 ) : ( n2299 ) ;
assign n2301 =  ( n1958 ) ? ( iram_83 ) : ( n2300 ) ;
assign n2302 =  ( n1957 ) ? ( iram_82 ) : ( n2301 ) ;
assign n2303 =  ( n1956 ) ? ( iram_81 ) : ( n2302 ) ;
assign n2304 =  ( n1955 ) ? ( iram_80 ) : ( n2303 ) ;
assign n2305 =  ( n1954 ) ? ( iram_79 ) : ( n2304 ) ;
assign n2306 =  ( n1953 ) ? ( iram_78 ) : ( n2305 ) ;
assign n2307 =  ( n1952 ) ? ( iram_77 ) : ( n2306 ) ;
assign n2308 =  ( n1951 ) ? ( iram_76 ) : ( n2307 ) ;
assign n2309 =  ( n1950 ) ? ( iram_75 ) : ( n2308 ) ;
assign n2310 =  ( n1949 ) ? ( iram_74 ) : ( n2309 ) ;
assign n2311 =  ( n1948 ) ? ( iram_73 ) : ( n2310 ) ;
assign n2312 =  ( n1947 ) ? ( iram_72 ) : ( n2311 ) ;
assign n2313 =  ( n1946 ) ? ( iram_71 ) : ( n2312 ) ;
assign n2314 =  ( n1945 ) ? ( iram_70 ) : ( n2313 ) ;
assign n2315 =  ( n1944 ) ? ( iram_69 ) : ( n2314 ) ;
assign n2316 =  ( n1943 ) ? ( iram_68 ) : ( n2315 ) ;
assign n2317 =  ( n1942 ) ? ( iram_67 ) : ( n2316 ) ;
assign n2318 =  ( n1941 ) ? ( iram_66 ) : ( n2317 ) ;
assign n2319 =  ( n1940 ) ? ( iram_65 ) : ( n2318 ) ;
assign n2320 =  ( n1939 ) ? ( iram_64 ) : ( n2319 ) ;
assign n2321 =  ( n1938 ) ? ( iram_63 ) : ( n2320 ) ;
assign n2322 =  ( n1937 ) ? ( iram_62 ) : ( n2321 ) ;
assign n2323 =  ( n1936 ) ? ( iram_61 ) : ( n2322 ) ;
assign n2324 =  ( n1935 ) ? ( iram_60 ) : ( n2323 ) ;
assign n2325 =  ( n1934 ) ? ( iram_59 ) : ( n2324 ) ;
assign n2326 =  ( n1933 ) ? ( iram_58 ) : ( n2325 ) ;
assign n2327 =  ( n1932 ) ? ( iram_57 ) : ( n2326 ) ;
assign n2328 =  ( n1931 ) ? ( iram_56 ) : ( n2327 ) ;
assign n2329 =  ( n1930 ) ? ( iram_55 ) : ( n2328 ) ;
assign n2330 =  ( n1929 ) ? ( iram_54 ) : ( n2329 ) ;
assign n2331 =  ( n1928 ) ? ( iram_53 ) : ( n2330 ) ;
assign n2332 =  ( n1927 ) ? ( iram_52 ) : ( n2331 ) ;
assign n2333 =  ( n1926 ) ? ( iram_51 ) : ( n2332 ) ;
assign n2334 =  ( n1925 ) ? ( iram_50 ) : ( n2333 ) ;
assign n2335 =  ( n1924 ) ? ( iram_49 ) : ( n2334 ) ;
assign n2336 =  ( n1923 ) ? ( iram_48 ) : ( n2335 ) ;
assign n2337 =  ( n1922 ) ? ( iram_47 ) : ( n2336 ) ;
assign n2338 =  ( n1921 ) ? ( iram_46 ) : ( n2337 ) ;
assign n2339 =  ( n1920 ) ? ( iram_45 ) : ( n2338 ) ;
assign n2340 =  ( n1919 ) ? ( iram_44 ) : ( n2339 ) ;
assign n2341 =  ( n1918 ) ? ( iram_43 ) : ( n2340 ) ;
assign n2342 =  ( n1917 ) ? ( iram_42 ) : ( n2341 ) ;
assign n2343 =  ( n1916 ) ? ( iram_41 ) : ( n2342 ) ;
assign n2344 =  ( n1915 ) ? ( iram_40 ) : ( n2343 ) ;
assign n2345 =  ( n1914 ) ? ( iram_39 ) : ( n2344 ) ;
assign n2346 =  ( n1913 ) ? ( iram_38 ) : ( n2345 ) ;
assign n2347 =  ( n1912 ) ? ( iram_37 ) : ( n2346 ) ;
assign n2348 =  ( n1911 ) ? ( iram_36 ) : ( n2347 ) ;
assign n2349 =  ( n1910 ) ? ( iram_35 ) : ( n2348 ) ;
assign n2350 =  ( n1909 ) ? ( iram_34 ) : ( n2349 ) ;
assign n2351 =  ( n1908 ) ? ( iram_33 ) : ( n2350 ) ;
assign n2352 =  ( n1907 ) ? ( iram_32 ) : ( n2351 ) ;
assign n2353 =  ( n1906 ) ? ( iram_31 ) : ( n2352 ) ;
assign n2354 =  ( n1905 ) ? ( iram_30 ) : ( n2353 ) ;
assign n2355 =  ( n1904 ) ? ( iram_29 ) : ( n2354 ) ;
assign n2356 =  ( n1903 ) ? ( iram_28 ) : ( n2355 ) ;
assign n2357 =  ( n1902 ) ? ( iram_27 ) : ( n2356 ) ;
assign n2358 =  ( n1901 ) ? ( iram_26 ) : ( n2357 ) ;
assign n2359 =  ( n1900 ) ? ( iram_25 ) : ( n2358 ) ;
assign n2360 =  ( n1899 ) ? ( iram_24 ) : ( n2359 ) ;
assign n2361 =  ( n1898 ) ? ( iram_23 ) : ( n2360 ) ;
assign n2362 =  ( n1897 ) ? ( iram_22 ) : ( n2361 ) ;
assign n2363 =  ( n1896 ) ? ( iram_21 ) : ( n2362 ) ;
assign n2364 =  ( n1895 ) ? ( iram_20 ) : ( n2363 ) ;
assign n2365 =  ( n1894 ) ? ( iram_19 ) : ( n2364 ) ;
assign n2366 =  ( n1893 ) ? ( iram_18 ) : ( n2365 ) ;
assign n2367 =  ( n1892 ) ? ( iram_17 ) : ( n2366 ) ;
assign n2368 =  ( n1891 ) ? ( iram_16 ) : ( n2367 ) ;
assign n2369 =  ( n1890 ) ? ( iram_15 ) : ( n2368 ) ;
assign n2370 =  ( n1889 ) ? ( iram_14 ) : ( n2369 ) ;
assign n2371 =  ( n1888 ) ? ( iram_13 ) : ( n2370 ) ;
assign n2372 =  ( n1887 ) ? ( iram_12 ) : ( n2371 ) ;
assign n2373 =  ( n1886 ) ? ( iram_11 ) : ( n2372 ) ;
assign n2374 =  ( n1885 ) ? ( iram_10 ) : ( n2373 ) ;
assign n2375 =  ( n1884 ) ? ( iram_9 ) : ( n2374 ) ;
assign n2376 =  ( n1883 ) ? ( iram_8 ) : ( n2375 ) ;
assign n2377 =  ( n1882 ) ? ( iram_7 ) : ( n2376 ) ;
assign n2378 =  ( n1881 ) ? ( iram_6 ) : ( n2377 ) ;
assign n2379 =  ( n1880 ) ? ( iram_5 ) : ( n2378 ) ;
assign n2380 =  ( n1879 ) ? ( iram_4 ) : ( n2379 ) ;
assign n2381 =  ( n1878 ) ? ( iram_3 ) : ( n2380 ) ;
assign n2382 =  ( n1877 ) ? ( iram_2 ) : ( n2381 ) ;
assign n2383 =  ( n1876 ) ? ( iram_1 ) : ( n2382 ) ;
assign n2384 =  ( n1875 ) ? ( iram_0 ) : ( n2383 ) ;
assign n2385 = rd_addr[7:7] ;
assign n2386 =  ( n2385 ) == ( bv_1_1_n34 )  ;
assign n2387 = rd_addr[6:3] ;
assign n2388 =  { ( bv_1_1_n34 ) , ( n2387 ) }  ;
assign n2389 =  { ( n2388 ) , ( bv_3_0_n46 ) }  ;
assign n2390 = rd_addr[6:3] ;
assign n2391 =  { ( bv_4_2_n12 ) , ( n2390 ) }  ;
assign n2392 =  ( n2386 ) ? ( n2389 ) : ( n2391 ) ;
assign n2393 =  ( bit_addr ) ? ( n2392 ) : ( rd_addr ) ;
assign n2394 = wr_addr[7:7] ;
assign n2395 =  ( n2394 ) == ( bv_1_1_n34 )  ;
assign n2396 = wr_addr[6:3] ;
assign n2397 =  { ( bv_1_1_n34 ) , ( n2396 ) }  ;
assign n2398 =  { ( n2397 ) , ( bv_3_0_n46 ) }  ;
assign n2399 = wr_addr[6:3] ;
assign n2400 =  { ( bv_4_2_n12 ) , ( n2399 ) }  ;
assign n2401 =  ( n2395 ) ? ( n2398 ) : ( n2400 ) ;
assign n2402 =  ( bit_addr_r ) ? ( n2401 ) : ( wr_addr ) ;
assign n2403 =  ( n2393 ) == ( n2402 )  ;
assign n2404 = n2393[7:0] ;
assign n2405 =  ( n2404 ) == ( bv_8_0_n69 )  ;
assign n2406 =  ( n2404 ) == ( bv_8_1_n71 )  ;
assign n2407 =  ( n2404 ) == ( bv_8_2_n73 )  ;
assign n2408 =  ( n2404 ) == ( bv_8_3_n75 )  ;
assign n2409 =  ( n2404 ) == ( bv_8_4_n77 )  ;
assign n2410 =  ( n2404 ) == ( bv_8_5_n79 )  ;
assign n2411 =  ( n2404 ) == ( bv_8_6_n81 )  ;
assign n2412 =  ( n2404 ) == ( bv_8_7_n83 )  ;
assign n2413 =  ( n2404 ) == ( bv_8_8_n85 )  ;
assign n2414 =  ( n2404 ) == ( bv_8_9_n87 )  ;
assign n2415 =  ( n2404 ) == ( bv_8_10_n89 )  ;
assign n2416 =  ( n2404 ) == ( bv_8_11_n91 )  ;
assign n2417 =  ( n2404 ) == ( bv_8_12_n93 )  ;
assign n2418 =  ( n2404 ) == ( bv_8_13_n95 )  ;
assign n2419 =  ( n2404 ) == ( bv_8_14_n97 )  ;
assign n2420 =  ( n2404 ) == ( bv_8_15_n99 )  ;
assign n2421 =  ( n2404 ) == ( bv_8_16_n101 )  ;
assign n2422 =  ( n2404 ) == ( bv_8_17_n103 )  ;
assign n2423 =  ( n2404 ) == ( bv_8_18_n105 )  ;
assign n2424 =  ( n2404 ) == ( bv_8_19_n107 )  ;
assign n2425 =  ( n2404 ) == ( bv_8_20_n109 )  ;
assign n2426 =  ( n2404 ) == ( bv_8_21_n111 )  ;
assign n2427 =  ( n2404 ) == ( bv_8_22_n113 )  ;
assign n2428 =  ( n2404 ) == ( bv_8_23_n115 )  ;
assign n2429 =  ( n2404 ) == ( bv_8_24_n117 )  ;
assign n2430 =  ( n2404 ) == ( bv_8_25_n119 )  ;
assign n2431 =  ( n2404 ) == ( bv_8_26_n121 )  ;
assign n2432 =  ( n2404 ) == ( bv_8_27_n123 )  ;
assign n2433 =  ( n2404 ) == ( bv_8_28_n125 )  ;
assign n2434 =  ( n2404 ) == ( bv_8_29_n127 )  ;
assign n2435 =  ( n2404 ) == ( bv_8_30_n129 )  ;
assign n2436 =  ( n2404 ) == ( bv_8_31_n131 )  ;
assign n2437 =  ( n2404 ) == ( bv_8_32_n133 )  ;
assign n2438 =  ( n2404 ) == ( bv_8_33_n135 )  ;
assign n2439 =  ( n2404 ) == ( bv_8_34_n137 )  ;
assign n2440 =  ( n2404 ) == ( bv_8_35_n139 )  ;
assign n2441 =  ( n2404 ) == ( bv_8_36_n141 )  ;
assign n2442 =  ( n2404 ) == ( bv_8_37_n143 )  ;
assign n2443 =  ( n2404 ) == ( bv_8_38_n145 )  ;
assign n2444 =  ( n2404 ) == ( bv_8_39_n147 )  ;
assign n2445 =  ( n2404 ) == ( bv_8_40_n149 )  ;
assign n2446 =  ( n2404 ) == ( bv_8_41_n151 )  ;
assign n2447 =  ( n2404 ) == ( bv_8_42_n153 )  ;
assign n2448 =  ( n2404 ) == ( bv_8_43_n155 )  ;
assign n2449 =  ( n2404 ) == ( bv_8_44_n157 )  ;
assign n2450 =  ( n2404 ) == ( bv_8_45_n159 )  ;
assign n2451 =  ( n2404 ) == ( bv_8_46_n161 )  ;
assign n2452 =  ( n2404 ) == ( bv_8_47_n163 )  ;
assign n2453 =  ( n2404 ) == ( bv_8_48_n165 )  ;
assign n2454 =  ( n2404 ) == ( bv_8_49_n167 )  ;
assign n2455 =  ( n2404 ) == ( bv_8_50_n169 )  ;
assign n2456 =  ( n2404 ) == ( bv_8_51_n171 )  ;
assign n2457 =  ( n2404 ) == ( bv_8_52_n173 )  ;
assign n2458 =  ( n2404 ) == ( bv_8_53_n175 )  ;
assign n2459 =  ( n2404 ) == ( bv_8_54_n177 )  ;
assign n2460 =  ( n2404 ) == ( bv_8_55_n179 )  ;
assign n2461 =  ( n2404 ) == ( bv_8_56_n181 )  ;
assign n2462 =  ( n2404 ) == ( bv_8_57_n183 )  ;
assign n2463 =  ( n2404 ) == ( bv_8_58_n185 )  ;
assign n2464 =  ( n2404 ) == ( bv_8_59_n187 )  ;
assign n2465 =  ( n2404 ) == ( bv_8_60_n189 )  ;
assign n2466 =  ( n2404 ) == ( bv_8_61_n191 )  ;
assign n2467 =  ( n2404 ) == ( bv_8_62_n193 )  ;
assign n2468 =  ( n2404 ) == ( bv_8_63_n195 )  ;
assign n2469 =  ( n2404 ) == ( bv_8_64_n197 )  ;
assign n2470 =  ( n2404 ) == ( bv_8_65_n199 )  ;
assign n2471 =  ( n2404 ) == ( bv_8_66_n201 )  ;
assign n2472 =  ( n2404 ) == ( bv_8_67_n203 )  ;
assign n2473 =  ( n2404 ) == ( bv_8_68_n205 )  ;
assign n2474 =  ( n2404 ) == ( bv_8_69_n207 )  ;
assign n2475 =  ( n2404 ) == ( bv_8_70_n209 )  ;
assign n2476 =  ( n2404 ) == ( bv_8_71_n211 )  ;
assign n2477 =  ( n2404 ) == ( bv_8_72_n213 )  ;
assign n2478 =  ( n2404 ) == ( bv_8_73_n215 )  ;
assign n2479 =  ( n2404 ) == ( bv_8_74_n217 )  ;
assign n2480 =  ( n2404 ) == ( bv_8_75_n219 )  ;
assign n2481 =  ( n2404 ) == ( bv_8_76_n221 )  ;
assign n2482 =  ( n2404 ) == ( bv_8_77_n223 )  ;
assign n2483 =  ( n2404 ) == ( bv_8_78_n225 )  ;
assign n2484 =  ( n2404 ) == ( bv_8_79_n227 )  ;
assign n2485 =  ( n2404 ) == ( bv_8_80_n229 )  ;
assign n2486 =  ( n2404 ) == ( bv_8_81_n231 )  ;
assign n2487 =  ( n2404 ) == ( bv_8_82_n233 )  ;
assign n2488 =  ( n2404 ) == ( bv_8_83_n235 )  ;
assign n2489 =  ( n2404 ) == ( bv_8_84_n237 )  ;
assign n2490 =  ( n2404 ) == ( bv_8_85_n239 )  ;
assign n2491 =  ( n2404 ) == ( bv_8_86_n241 )  ;
assign n2492 =  ( n2404 ) == ( bv_8_87_n243 )  ;
assign n2493 =  ( n2404 ) == ( bv_8_88_n245 )  ;
assign n2494 =  ( n2404 ) == ( bv_8_89_n247 )  ;
assign n2495 =  ( n2404 ) == ( bv_8_90_n249 )  ;
assign n2496 =  ( n2404 ) == ( bv_8_91_n251 )  ;
assign n2497 =  ( n2404 ) == ( bv_8_92_n253 )  ;
assign n2498 =  ( n2404 ) == ( bv_8_93_n255 )  ;
assign n2499 =  ( n2404 ) == ( bv_8_94_n257 )  ;
assign n2500 =  ( n2404 ) == ( bv_8_95_n259 )  ;
assign n2501 =  ( n2404 ) == ( bv_8_96_n261 )  ;
assign n2502 =  ( n2404 ) == ( bv_8_97_n263 )  ;
assign n2503 =  ( n2404 ) == ( bv_8_98_n265 )  ;
assign n2504 =  ( n2404 ) == ( bv_8_99_n267 )  ;
assign n2505 =  ( n2404 ) == ( bv_8_100_n269 )  ;
assign n2506 =  ( n2404 ) == ( bv_8_101_n271 )  ;
assign n2507 =  ( n2404 ) == ( bv_8_102_n273 )  ;
assign n2508 =  ( n2404 ) == ( bv_8_103_n275 )  ;
assign n2509 =  ( n2404 ) == ( bv_8_104_n277 )  ;
assign n2510 =  ( n2404 ) == ( bv_8_105_n279 )  ;
assign n2511 =  ( n2404 ) == ( bv_8_106_n281 )  ;
assign n2512 =  ( n2404 ) == ( bv_8_107_n283 )  ;
assign n2513 =  ( n2404 ) == ( bv_8_108_n285 )  ;
assign n2514 =  ( n2404 ) == ( bv_8_109_n287 )  ;
assign n2515 =  ( n2404 ) == ( bv_8_110_n289 )  ;
assign n2516 =  ( n2404 ) == ( bv_8_111_n291 )  ;
assign n2517 =  ( n2404 ) == ( bv_8_112_n293 )  ;
assign n2518 =  ( n2404 ) == ( bv_8_113_n295 )  ;
assign n2519 =  ( n2404 ) == ( bv_8_114_n297 )  ;
assign n2520 =  ( n2404 ) == ( bv_8_115_n299 )  ;
assign n2521 =  ( n2404 ) == ( bv_8_116_n301 )  ;
assign n2522 =  ( n2404 ) == ( bv_8_117_n303 )  ;
assign n2523 =  ( n2404 ) == ( bv_8_118_n305 )  ;
assign n2524 =  ( n2404 ) == ( bv_8_119_n307 )  ;
assign n2525 =  ( n2404 ) == ( bv_8_120_n309 )  ;
assign n2526 =  ( n2404 ) == ( bv_8_121_n311 )  ;
assign n2527 =  ( n2404 ) == ( bv_8_122_n313 )  ;
assign n2528 =  ( n2404 ) == ( bv_8_123_n315 )  ;
assign n2529 =  ( n2404 ) == ( bv_8_124_n317 )  ;
assign n2530 =  ( n2404 ) == ( bv_8_125_n319 )  ;
assign n2531 =  ( n2404 ) == ( bv_8_126_n321 )  ;
assign n2532 =  ( n2404 ) == ( bv_8_127_n323 )  ;
assign n2533 =  ( n2404 ) == ( bv_8_128_n325 )  ;
assign n2534 =  ( n2404 ) == ( bv_8_129_n327 )  ;
assign n2535 =  ( n2404 ) == ( bv_8_130_n329 )  ;
assign n2536 =  ( n2404 ) == ( bv_8_131_n331 )  ;
assign n2537 =  ( n2404 ) == ( bv_8_132_n333 )  ;
assign n2538 =  ( n2404 ) == ( bv_8_133_n335 )  ;
assign n2539 =  ( n2404 ) == ( bv_8_134_n337 )  ;
assign n2540 =  ( n2404 ) == ( bv_8_135_n339 )  ;
assign n2541 =  ( n2404 ) == ( bv_8_136_n341 )  ;
assign n2542 =  ( n2404 ) == ( bv_8_137_n343 )  ;
assign n2543 =  ( n2404 ) == ( bv_8_138_n345 )  ;
assign n2544 =  ( n2404 ) == ( bv_8_139_n347 )  ;
assign n2545 =  ( n2404 ) == ( bv_8_140_n349 )  ;
assign n2546 =  ( n2404 ) == ( bv_8_141_n351 )  ;
assign n2547 =  ( n2404 ) == ( bv_8_142_n353 )  ;
assign n2548 =  ( n2404 ) == ( bv_8_143_n355 )  ;
assign n2549 =  ( n2404 ) == ( bv_8_144_n357 )  ;
assign n2550 =  ( n2404 ) == ( bv_8_145_n359 )  ;
assign n2551 =  ( n2404 ) == ( bv_8_146_n361 )  ;
assign n2552 =  ( n2404 ) == ( bv_8_147_n363 )  ;
assign n2553 =  ( n2404 ) == ( bv_8_148_n365 )  ;
assign n2554 =  ( n2404 ) == ( bv_8_149_n367 )  ;
assign n2555 =  ( n2404 ) == ( bv_8_150_n369 )  ;
assign n2556 =  ( n2404 ) == ( bv_8_151_n371 )  ;
assign n2557 =  ( n2404 ) == ( bv_8_152_n373 )  ;
assign n2558 =  ( n2404 ) == ( bv_8_153_n375 )  ;
assign n2559 =  ( n2404 ) == ( bv_8_154_n377 )  ;
assign n2560 =  ( n2404 ) == ( bv_8_155_n379 )  ;
assign n2561 =  ( n2404 ) == ( bv_8_156_n381 )  ;
assign n2562 =  ( n2404 ) == ( bv_8_157_n383 )  ;
assign n2563 =  ( n2404 ) == ( bv_8_158_n385 )  ;
assign n2564 =  ( n2404 ) == ( bv_8_159_n387 )  ;
assign n2565 =  ( n2404 ) == ( bv_8_160_n389 )  ;
assign n2566 =  ( n2404 ) == ( bv_8_161_n391 )  ;
assign n2567 =  ( n2404 ) == ( bv_8_162_n393 )  ;
assign n2568 =  ( n2404 ) == ( bv_8_163_n395 )  ;
assign n2569 =  ( n2404 ) == ( bv_8_164_n397 )  ;
assign n2570 =  ( n2404 ) == ( bv_8_165_n399 )  ;
assign n2571 =  ( n2404 ) == ( bv_8_166_n401 )  ;
assign n2572 =  ( n2404 ) == ( bv_8_167_n403 )  ;
assign n2573 =  ( n2404 ) == ( bv_8_168_n405 )  ;
assign n2574 =  ( n2404 ) == ( bv_8_169_n407 )  ;
assign n2575 =  ( n2404 ) == ( bv_8_170_n409 )  ;
assign n2576 =  ( n2404 ) == ( bv_8_171_n411 )  ;
assign n2577 =  ( n2404 ) == ( bv_8_172_n413 )  ;
assign n2578 =  ( n2404 ) == ( bv_8_173_n415 )  ;
assign n2579 =  ( n2404 ) == ( bv_8_174_n417 )  ;
assign n2580 =  ( n2404 ) == ( bv_8_175_n419 )  ;
assign n2581 =  ( n2404 ) == ( bv_8_176_n421 )  ;
assign n2582 =  ( n2404 ) == ( bv_8_177_n423 )  ;
assign n2583 =  ( n2404 ) == ( bv_8_178_n425 )  ;
assign n2584 =  ( n2404 ) == ( bv_8_179_n427 )  ;
assign n2585 =  ( n2404 ) == ( bv_8_180_n429 )  ;
assign n2586 =  ( n2404 ) == ( bv_8_181_n431 )  ;
assign n2587 =  ( n2404 ) == ( bv_8_182_n433 )  ;
assign n2588 =  ( n2404 ) == ( bv_8_183_n435 )  ;
assign n2589 =  ( n2404 ) == ( bv_8_184_n437 )  ;
assign n2590 =  ( n2404 ) == ( bv_8_185_n439 )  ;
assign n2591 =  ( n2404 ) == ( bv_8_186_n441 )  ;
assign n2592 =  ( n2404 ) == ( bv_8_187_n443 )  ;
assign n2593 =  ( n2404 ) == ( bv_8_188_n445 )  ;
assign n2594 =  ( n2404 ) == ( bv_8_189_n447 )  ;
assign n2595 =  ( n2404 ) == ( bv_8_190_n449 )  ;
assign n2596 =  ( n2404 ) == ( bv_8_191_n451 )  ;
assign n2597 =  ( n2404 ) == ( bv_8_192_n453 )  ;
assign n2598 =  ( n2404 ) == ( bv_8_193_n455 )  ;
assign n2599 =  ( n2404 ) == ( bv_8_194_n457 )  ;
assign n2600 =  ( n2404 ) == ( bv_8_195_n459 )  ;
assign n2601 =  ( n2404 ) == ( bv_8_196_n461 )  ;
assign n2602 =  ( n2404 ) == ( bv_8_197_n463 )  ;
assign n2603 =  ( n2404 ) == ( bv_8_198_n465 )  ;
assign n2604 =  ( n2404 ) == ( bv_8_199_n467 )  ;
assign n2605 =  ( n2404 ) == ( bv_8_200_n469 )  ;
assign n2606 =  ( n2404 ) == ( bv_8_201_n471 )  ;
assign n2607 =  ( n2404 ) == ( bv_8_202_n473 )  ;
assign n2608 =  ( n2404 ) == ( bv_8_203_n475 )  ;
assign n2609 =  ( n2404 ) == ( bv_8_204_n477 )  ;
assign n2610 =  ( n2404 ) == ( bv_8_205_n479 )  ;
assign n2611 =  ( n2404 ) == ( bv_8_206_n481 )  ;
assign n2612 =  ( n2404 ) == ( bv_8_207_n483 )  ;
assign n2613 =  ( n2404 ) == ( bv_8_208_n485 )  ;
assign n2614 =  ( n2404 ) == ( bv_8_209_n487 )  ;
assign n2615 =  ( n2404 ) == ( bv_8_210_n489 )  ;
assign n2616 =  ( n2404 ) == ( bv_8_211_n491 )  ;
assign n2617 =  ( n2404 ) == ( bv_8_212_n493 )  ;
assign n2618 =  ( n2404 ) == ( bv_8_213_n495 )  ;
assign n2619 =  ( n2404 ) == ( bv_8_214_n497 )  ;
assign n2620 =  ( n2404 ) == ( bv_8_215_n499 )  ;
assign n2621 =  ( n2404 ) == ( bv_8_216_n501 )  ;
assign n2622 =  ( n2404 ) == ( bv_8_217_n503 )  ;
assign n2623 =  ( n2404 ) == ( bv_8_218_n505 )  ;
assign n2624 =  ( n2404 ) == ( bv_8_219_n507 )  ;
assign n2625 =  ( n2404 ) == ( bv_8_220_n509 )  ;
assign n2626 =  ( n2404 ) == ( bv_8_221_n511 )  ;
assign n2627 =  ( n2404 ) == ( bv_8_222_n513 )  ;
assign n2628 =  ( n2404 ) == ( bv_8_223_n515 )  ;
assign n2629 =  ( n2404 ) == ( bv_8_224_n517 )  ;
assign n2630 =  ( n2404 ) == ( bv_8_225_n519 )  ;
assign n2631 =  ( n2404 ) == ( bv_8_226_n521 )  ;
assign n2632 =  ( n2404 ) == ( bv_8_227_n523 )  ;
assign n2633 =  ( n2404 ) == ( bv_8_228_n525 )  ;
assign n2634 =  ( n2404 ) == ( bv_8_229_n527 )  ;
assign n2635 =  ( n2404 ) == ( bv_8_230_n529 )  ;
assign n2636 =  ( n2404 ) == ( bv_8_231_n531 )  ;
assign n2637 =  ( n2404 ) == ( bv_8_232_n533 )  ;
assign n2638 =  ( n2404 ) == ( bv_8_233_n535 )  ;
assign n2639 =  ( n2404 ) == ( bv_8_234_n537 )  ;
assign n2640 =  ( n2404 ) == ( bv_8_235_n539 )  ;
assign n2641 =  ( n2404 ) == ( bv_8_236_n541 )  ;
assign n2642 =  ( n2404 ) == ( bv_8_237_n543 )  ;
assign n2643 =  ( n2404 ) == ( bv_8_238_n545 )  ;
assign n2644 =  ( n2404 ) == ( bv_8_239_n547 )  ;
assign n2645 =  ( n2404 ) == ( bv_8_240_n549 )  ;
assign n2646 =  ( n2404 ) == ( bv_8_241_n551 )  ;
assign n2647 =  ( n2404 ) == ( bv_8_242_n553 )  ;
assign n2648 =  ( n2404 ) == ( bv_8_243_n555 )  ;
assign n2649 =  ( n2404 ) == ( bv_8_244_n557 )  ;
assign n2650 =  ( n2404 ) == ( bv_8_245_n559 )  ;
assign n2651 =  ( n2404 ) == ( bv_8_246_n561 )  ;
assign n2652 =  ( n2404 ) == ( bv_8_247_n563 )  ;
assign n2653 =  ( n2404 ) == ( bv_8_248_n565 )  ;
assign n2654 =  ( n2404 ) == ( bv_8_249_n567 )  ;
assign n2655 =  ( n2404 ) == ( bv_8_250_n569 )  ;
assign n2656 =  ( n2404 ) == ( bv_8_251_n571 )  ;
assign n2657 =  ( n2404 ) == ( bv_8_252_n573 )  ;
assign n2658 =  ( n2404 ) == ( bv_8_253_n575 )  ;
assign n2659 =  ( n2404 ) == ( bv_8_254_n577 )  ;
assign n2660 =  ( n2659 ) ? ( iram_254 ) : ( iram_255 ) ;
assign n2661 =  ( n2658 ) ? ( iram_253 ) : ( n2660 ) ;
assign n2662 =  ( n2657 ) ? ( iram_252 ) : ( n2661 ) ;
assign n2663 =  ( n2656 ) ? ( iram_251 ) : ( n2662 ) ;
assign n2664 =  ( n2655 ) ? ( iram_250 ) : ( n2663 ) ;
assign n2665 =  ( n2654 ) ? ( iram_249 ) : ( n2664 ) ;
assign n2666 =  ( n2653 ) ? ( iram_248 ) : ( n2665 ) ;
assign n2667 =  ( n2652 ) ? ( iram_247 ) : ( n2666 ) ;
assign n2668 =  ( n2651 ) ? ( iram_246 ) : ( n2667 ) ;
assign n2669 =  ( n2650 ) ? ( iram_245 ) : ( n2668 ) ;
assign n2670 =  ( n2649 ) ? ( iram_244 ) : ( n2669 ) ;
assign n2671 =  ( n2648 ) ? ( iram_243 ) : ( n2670 ) ;
assign n2672 =  ( n2647 ) ? ( iram_242 ) : ( n2671 ) ;
assign n2673 =  ( n2646 ) ? ( iram_241 ) : ( n2672 ) ;
assign n2674 =  ( n2645 ) ? ( iram_240 ) : ( n2673 ) ;
assign n2675 =  ( n2644 ) ? ( iram_239 ) : ( n2674 ) ;
assign n2676 =  ( n2643 ) ? ( iram_238 ) : ( n2675 ) ;
assign n2677 =  ( n2642 ) ? ( iram_237 ) : ( n2676 ) ;
assign n2678 =  ( n2641 ) ? ( iram_236 ) : ( n2677 ) ;
assign n2679 =  ( n2640 ) ? ( iram_235 ) : ( n2678 ) ;
assign n2680 =  ( n2639 ) ? ( iram_234 ) : ( n2679 ) ;
assign n2681 =  ( n2638 ) ? ( iram_233 ) : ( n2680 ) ;
assign n2682 =  ( n2637 ) ? ( iram_232 ) : ( n2681 ) ;
assign n2683 =  ( n2636 ) ? ( iram_231 ) : ( n2682 ) ;
assign n2684 =  ( n2635 ) ? ( iram_230 ) : ( n2683 ) ;
assign n2685 =  ( n2634 ) ? ( iram_229 ) : ( n2684 ) ;
assign n2686 =  ( n2633 ) ? ( iram_228 ) : ( n2685 ) ;
assign n2687 =  ( n2632 ) ? ( iram_227 ) : ( n2686 ) ;
assign n2688 =  ( n2631 ) ? ( iram_226 ) : ( n2687 ) ;
assign n2689 =  ( n2630 ) ? ( iram_225 ) : ( n2688 ) ;
assign n2690 =  ( n2629 ) ? ( iram_224 ) : ( n2689 ) ;
assign n2691 =  ( n2628 ) ? ( iram_223 ) : ( n2690 ) ;
assign n2692 =  ( n2627 ) ? ( iram_222 ) : ( n2691 ) ;
assign n2693 =  ( n2626 ) ? ( iram_221 ) : ( n2692 ) ;
assign n2694 =  ( n2625 ) ? ( iram_220 ) : ( n2693 ) ;
assign n2695 =  ( n2624 ) ? ( iram_219 ) : ( n2694 ) ;
assign n2696 =  ( n2623 ) ? ( iram_218 ) : ( n2695 ) ;
assign n2697 =  ( n2622 ) ? ( iram_217 ) : ( n2696 ) ;
assign n2698 =  ( n2621 ) ? ( iram_216 ) : ( n2697 ) ;
assign n2699 =  ( n2620 ) ? ( iram_215 ) : ( n2698 ) ;
assign n2700 =  ( n2619 ) ? ( iram_214 ) : ( n2699 ) ;
assign n2701 =  ( n2618 ) ? ( iram_213 ) : ( n2700 ) ;
assign n2702 =  ( n2617 ) ? ( iram_212 ) : ( n2701 ) ;
assign n2703 =  ( n2616 ) ? ( iram_211 ) : ( n2702 ) ;
assign n2704 =  ( n2615 ) ? ( iram_210 ) : ( n2703 ) ;
assign n2705 =  ( n2614 ) ? ( iram_209 ) : ( n2704 ) ;
assign n2706 =  ( n2613 ) ? ( iram_208 ) : ( n2705 ) ;
assign n2707 =  ( n2612 ) ? ( iram_207 ) : ( n2706 ) ;
assign n2708 =  ( n2611 ) ? ( iram_206 ) : ( n2707 ) ;
assign n2709 =  ( n2610 ) ? ( iram_205 ) : ( n2708 ) ;
assign n2710 =  ( n2609 ) ? ( iram_204 ) : ( n2709 ) ;
assign n2711 =  ( n2608 ) ? ( iram_203 ) : ( n2710 ) ;
assign n2712 =  ( n2607 ) ? ( iram_202 ) : ( n2711 ) ;
assign n2713 =  ( n2606 ) ? ( iram_201 ) : ( n2712 ) ;
assign n2714 =  ( n2605 ) ? ( iram_200 ) : ( n2713 ) ;
assign n2715 =  ( n2604 ) ? ( iram_199 ) : ( n2714 ) ;
assign n2716 =  ( n2603 ) ? ( iram_198 ) : ( n2715 ) ;
assign n2717 =  ( n2602 ) ? ( iram_197 ) : ( n2716 ) ;
assign n2718 =  ( n2601 ) ? ( iram_196 ) : ( n2717 ) ;
assign n2719 =  ( n2600 ) ? ( iram_195 ) : ( n2718 ) ;
assign n2720 =  ( n2599 ) ? ( iram_194 ) : ( n2719 ) ;
assign n2721 =  ( n2598 ) ? ( iram_193 ) : ( n2720 ) ;
assign n2722 =  ( n2597 ) ? ( iram_192 ) : ( n2721 ) ;
assign n2723 =  ( n2596 ) ? ( iram_191 ) : ( n2722 ) ;
assign n2724 =  ( n2595 ) ? ( iram_190 ) : ( n2723 ) ;
assign n2725 =  ( n2594 ) ? ( iram_189 ) : ( n2724 ) ;
assign n2726 =  ( n2593 ) ? ( iram_188 ) : ( n2725 ) ;
assign n2727 =  ( n2592 ) ? ( iram_187 ) : ( n2726 ) ;
assign n2728 =  ( n2591 ) ? ( iram_186 ) : ( n2727 ) ;
assign n2729 =  ( n2590 ) ? ( iram_185 ) : ( n2728 ) ;
assign n2730 =  ( n2589 ) ? ( iram_184 ) : ( n2729 ) ;
assign n2731 =  ( n2588 ) ? ( iram_183 ) : ( n2730 ) ;
assign n2732 =  ( n2587 ) ? ( iram_182 ) : ( n2731 ) ;
assign n2733 =  ( n2586 ) ? ( iram_181 ) : ( n2732 ) ;
assign n2734 =  ( n2585 ) ? ( iram_180 ) : ( n2733 ) ;
assign n2735 =  ( n2584 ) ? ( iram_179 ) : ( n2734 ) ;
assign n2736 =  ( n2583 ) ? ( iram_178 ) : ( n2735 ) ;
assign n2737 =  ( n2582 ) ? ( iram_177 ) : ( n2736 ) ;
assign n2738 =  ( n2581 ) ? ( iram_176 ) : ( n2737 ) ;
assign n2739 =  ( n2580 ) ? ( iram_175 ) : ( n2738 ) ;
assign n2740 =  ( n2579 ) ? ( iram_174 ) : ( n2739 ) ;
assign n2741 =  ( n2578 ) ? ( iram_173 ) : ( n2740 ) ;
assign n2742 =  ( n2577 ) ? ( iram_172 ) : ( n2741 ) ;
assign n2743 =  ( n2576 ) ? ( iram_171 ) : ( n2742 ) ;
assign n2744 =  ( n2575 ) ? ( iram_170 ) : ( n2743 ) ;
assign n2745 =  ( n2574 ) ? ( iram_169 ) : ( n2744 ) ;
assign n2746 =  ( n2573 ) ? ( iram_168 ) : ( n2745 ) ;
assign n2747 =  ( n2572 ) ? ( iram_167 ) : ( n2746 ) ;
assign n2748 =  ( n2571 ) ? ( iram_166 ) : ( n2747 ) ;
assign n2749 =  ( n2570 ) ? ( iram_165 ) : ( n2748 ) ;
assign n2750 =  ( n2569 ) ? ( iram_164 ) : ( n2749 ) ;
assign n2751 =  ( n2568 ) ? ( iram_163 ) : ( n2750 ) ;
assign n2752 =  ( n2567 ) ? ( iram_162 ) : ( n2751 ) ;
assign n2753 =  ( n2566 ) ? ( iram_161 ) : ( n2752 ) ;
assign n2754 =  ( n2565 ) ? ( iram_160 ) : ( n2753 ) ;
assign n2755 =  ( n2564 ) ? ( iram_159 ) : ( n2754 ) ;
assign n2756 =  ( n2563 ) ? ( iram_158 ) : ( n2755 ) ;
assign n2757 =  ( n2562 ) ? ( iram_157 ) : ( n2756 ) ;
assign n2758 =  ( n2561 ) ? ( iram_156 ) : ( n2757 ) ;
assign n2759 =  ( n2560 ) ? ( iram_155 ) : ( n2758 ) ;
assign n2760 =  ( n2559 ) ? ( iram_154 ) : ( n2759 ) ;
assign n2761 =  ( n2558 ) ? ( iram_153 ) : ( n2760 ) ;
assign n2762 =  ( n2557 ) ? ( iram_152 ) : ( n2761 ) ;
assign n2763 =  ( n2556 ) ? ( iram_151 ) : ( n2762 ) ;
assign n2764 =  ( n2555 ) ? ( iram_150 ) : ( n2763 ) ;
assign n2765 =  ( n2554 ) ? ( iram_149 ) : ( n2764 ) ;
assign n2766 =  ( n2553 ) ? ( iram_148 ) : ( n2765 ) ;
assign n2767 =  ( n2552 ) ? ( iram_147 ) : ( n2766 ) ;
assign n2768 =  ( n2551 ) ? ( iram_146 ) : ( n2767 ) ;
assign n2769 =  ( n2550 ) ? ( iram_145 ) : ( n2768 ) ;
assign n2770 =  ( n2549 ) ? ( iram_144 ) : ( n2769 ) ;
assign n2771 =  ( n2548 ) ? ( iram_143 ) : ( n2770 ) ;
assign n2772 =  ( n2547 ) ? ( iram_142 ) : ( n2771 ) ;
assign n2773 =  ( n2546 ) ? ( iram_141 ) : ( n2772 ) ;
assign n2774 =  ( n2545 ) ? ( iram_140 ) : ( n2773 ) ;
assign n2775 =  ( n2544 ) ? ( iram_139 ) : ( n2774 ) ;
assign n2776 =  ( n2543 ) ? ( iram_138 ) : ( n2775 ) ;
assign n2777 =  ( n2542 ) ? ( iram_137 ) : ( n2776 ) ;
assign n2778 =  ( n2541 ) ? ( iram_136 ) : ( n2777 ) ;
assign n2779 =  ( n2540 ) ? ( iram_135 ) : ( n2778 ) ;
assign n2780 =  ( n2539 ) ? ( iram_134 ) : ( n2779 ) ;
assign n2781 =  ( n2538 ) ? ( iram_133 ) : ( n2780 ) ;
assign n2782 =  ( n2537 ) ? ( iram_132 ) : ( n2781 ) ;
assign n2783 =  ( n2536 ) ? ( iram_131 ) : ( n2782 ) ;
assign n2784 =  ( n2535 ) ? ( iram_130 ) : ( n2783 ) ;
assign n2785 =  ( n2534 ) ? ( iram_129 ) : ( n2784 ) ;
assign n2786 =  ( n2533 ) ? ( iram_128 ) : ( n2785 ) ;
assign n2787 =  ( n2532 ) ? ( iram_127 ) : ( n2786 ) ;
assign n2788 =  ( n2531 ) ? ( iram_126 ) : ( n2787 ) ;
assign n2789 =  ( n2530 ) ? ( iram_125 ) : ( n2788 ) ;
assign n2790 =  ( n2529 ) ? ( iram_124 ) : ( n2789 ) ;
assign n2791 =  ( n2528 ) ? ( iram_123 ) : ( n2790 ) ;
assign n2792 =  ( n2527 ) ? ( iram_122 ) : ( n2791 ) ;
assign n2793 =  ( n2526 ) ? ( iram_121 ) : ( n2792 ) ;
assign n2794 =  ( n2525 ) ? ( iram_120 ) : ( n2793 ) ;
assign n2795 =  ( n2524 ) ? ( iram_119 ) : ( n2794 ) ;
assign n2796 =  ( n2523 ) ? ( iram_118 ) : ( n2795 ) ;
assign n2797 =  ( n2522 ) ? ( iram_117 ) : ( n2796 ) ;
assign n2798 =  ( n2521 ) ? ( iram_116 ) : ( n2797 ) ;
assign n2799 =  ( n2520 ) ? ( iram_115 ) : ( n2798 ) ;
assign n2800 =  ( n2519 ) ? ( iram_114 ) : ( n2799 ) ;
assign n2801 =  ( n2518 ) ? ( iram_113 ) : ( n2800 ) ;
assign n2802 =  ( n2517 ) ? ( iram_112 ) : ( n2801 ) ;
assign n2803 =  ( n2516 ) ? ( iram_111 ) : ( n2802 ) ;
assign n2804 =  ( n2515 ) ? ( iram_110 ) : ( n2803 ) ;
assign n2805 =  ( n2514 ) ? ( iram_109 ) : ( n2804 ) ;
assign n2806 =  ( n2513 ) ? ( iram_108 ) : ( n2805 ) ;
assign n2807 =  ( n2512 ) ? ( iram_107 ) : ( n2806 ) ;
assign n2808 =  ( n2511 ) ? ( iram_106 ) : ( n2807 ) ;
assign n2809 =  ( n2510 ) ? ( iram_105 ) : ( n2808 ) ;
assign n2810 =  ( n2509 ) ? ( iram_104 ) : ( n2809 ) ;
assign n2811 =  ( n2508 ) ? ( iram_103 ) : ( n2810 ) ;
assign n2812 =  ( n2507 ) ? ( iram_102 ) : ( n2811 ) ;
assign n2813 =  ( n2506 ) ? ( iram_101 ) : ( n2812 ) ;
assign n2814 =  ( n2505 ) ? ( iram_100 ) : ( n2813 ) ;
assign n2815 =  ( n2504 ) ? ( iram_99 ) : ( n2814 ) ;
assign n2816 =  ( n2503 ) ? ( iram_98 ) : ( n2815 ) ;
assign n2817 =  ( n2502 ) ? ( iram_97 ) : ( n2816 ) ;
assign n2818 =  ( n2501 ) ? ( iram_96 ) : ( n2817 ) ;
assign n2819 =  ( n2500 ) ? ( iram_95 ) : ( n2818 ) ;
assign n2820 =  ( n2499 ) ? ( iram_94 ) : ( n2819 ) ;
assign n2821 =  ( n2498 ) ? ( iram_93 ) : ( n2820 ) ;
assign n2822 =  ( n2497 ) ? ( iram_92 ) : ( n2821 ) ;
assign n2823 =  ( n2496 ) ? ( iram_91 ) : ( n2822 ) ;
assign n2824 =  ( n2495 ) ? ( iram_90 ) : ( n2823 ) ;
assign n2825 =  ( n2494 ) ? ( iram_89 ) : ( n2824 ) ;
assign n2826 =  ( n2493 ) ? ( iram_88 ) : ( n2825 ) ;
assign n2827 =  ( n2492 ) ? ( iram_87 ) : ( n2826 ) ;
assign n2828 =  ( n2491 ) ? ( iram_86 ) : ( n2827 ) ;
assign n2829 =  ( n2490 ) ? ( iram_85 ) : ( n2828 ) ;
assign n2830 =  ( n2489 ) ? ( iram_84 ) : ( n2829 ) ;
assign n2831 =  ( n2488 ) ? ( iram_83 ) : ( n2830 ) ;
assign n2832 =  ( n2487 ) ? ( iram_82 ) : ( n2831 ) ;
assign n2833 =  ( n2486 ) ? ( iram_81 ) : ( n2832 ) ;
assign n2834 =  ( n2485 ) ? ( iram_80 ) : ( n2833 ) ;
assign n2835 =  ( n2484 ) ? ( iram_79 ) : ( n2834 ) ;
assign n2836 =  ( n2483 ) ? ( iram_78 ) : ( n2835 ) ;
assign n2837 =  ( n2482 ) ? ( iram_77 ) : ( n2836 ) ;
assign n2838 =  ( n2481 ) ? ( iram_76 ) : ( n2837 ) ;
assign n2839 =  ( n2480 ) ? ( iram_75 ) : ( n2838 ) ;
assign n2840 =  ( n2479 ) ? ( iram_74 ) : ( n2839 ) ;
assign n2841 =  ( n2478 ) ? ( iram_73 ) : ( n2840 ) ;
assign n2842 =  ( n2477 ) ? ( iram_72 ) : ( n2841 ) ;
assign n2843 =  ( n2476 ) ? ( iram_71 ) : ( n2842 ) ;
assign n2844 =  ( n2475 ) ? ( iram_70 ) : ( n2843 ) ;
assign n2845 =  ( n2474 ) ? ( iram_69 ) : ( n2844 ) ;
assign n2846 =  ( n2473 ) ? ( iram_68 ) : ( n2845 ) ;
assign n2847 =  ( n2472 ) ? ( iram_67 ) : ( n2846 ) ;
assign n2848 =  ( n2471 ) ? ( iram_66 ) : ( n2847 ) ;
assign n2849 =  ( n2470 ) ? ( iram_65 ) : ( n2848 ) ;
assign n2850 =  ( n2469 ) ? ( iram_64 ) : ( n2849 ) ;
assign n2851 =  ( n2468 ) ? ( iram_63 ) : ( n2850 ) ;
assign n2852 =  ( n2467 ) ? ( iram_62 ) : ( n2851 ) ;
assign n2853 =  ( n2466 ) ? ( iram_61 ) : ( n2852 ) ;
assign n2854 =  ( n2465 ) ? ( iram_60 ) : ( n2853 ) ;
assign n2855 =  ( n2464 ) ? ( iram_59 ) : ( n2854 ) ;
assign n2856 =  ( n2463 ) ? ( iram_58 ) : ( n2855 ) ;
assign n2857 =  ( n2462 ) ? ( iram_57 ) : ( n2856 ) ;
assign n2858 =  ( n2461 ) ? ( iram_56 ) : ( n2857 ) ;
assign n2859 =  ( n2460 ) ? ( iram_55 ) : ( n2858 ) ;
assign n2860 =  ( n2459 ) ? ( iram_54 ) : ( n2859 ) ;
assign n2861 =  ( n2458 ) ? ( iram_53 ) : ( n2860 ) ;
assign n2862 =  ( n2457 ) ? ( iram_52 ) : ( n2861 ) ;
assign n2863 =  ( n2456 ) ? ( iram_51 ) : ( n2862 ) ;
assign n2864 =  ( n2455 ) ? ( iram_50 ) : ( n2863 ) ;
assign n2865 =  ( n2454 ) ? ( iram_49 ) : ( n2864 ) ;
assign n2866 =  ( n2453 ) ? ( iram_48 ) : ( n2865 ) ;
assign n2867 =  ( n2452 ) ? ( iram_47 ) : ( n2866 ) ;
assign n2868 =  ( n2451 ) ? ( iram_46 ) : ( n2867 ) ;
assign n2869 =  ( n2450 ) ? ( iram_45 ) : ( n2868 ) ;
assign n2870 =  ( n2449 ) ? ( iram_44 ) : ( n2869 ) ;
assign n2871 =  ( n2448 ) ? ( iram_43 ) : ( n2870 ) ;
assign n2872 =  ( n2447 ) ? ( iram_42 ) : ( n2871 ) ;
assign n2873 =  ( n2446 ) ? ( iram_41 ) : ( n2872 ) ;
assign n2874 =  ( n2445 ) ? ( iram_40 ) : ( n2873 ) ;
assign n2875 =  ( n2444 ) ? ( iram_39 ) : ( n2874 ) ;
assign n2876 =  ( n2443 ) ? ( iram_38 ) : ( n2875 ) ;
assign n2877 =  ( n2442 ) ? ( iram_37 ) : ( n2876 ) ;
assign n2878 =  ( n2441 ) ? ( iram_36 ) : ( n2877 ) ;
assign n2879 =  ( n2440 ) ? ( iram_35 ) : ( n2878 ) ;
assign n2880 =  ( n2439 ) ? ( iram_34 ) : ( n2879 ) ;
assign n2881 =  ( n2438 ) ? ( iram_33 ) : ( n2880 ) ;
assign n2882 =  ( n2437 ) ? ( iram_32 ) : ( n2881 ) ;
assign n2883 =  ( n2436 ) ? ( iram_31 ) : ( n2882 ) ;
assign n2884 =  ( n2435 ) ? ( iram_30 ) : ( n2883 ) ;
assign n2885 =  ( n2434 ) ? ( iram_29 ) : ( n2884 ) ;
assign n2886 =  ( n2433 ) ? ( iram_28 ) : ( n2885 ) ;
assign n2887 =  ( n2432 ) ? ( iram_27 ) : ( n2886 ) ;
assign n2888 =  ( n2431 ) ? ( iram_26 ) : ( n2887 ) ;
assign n2889 =  ( n2430 ) ? ( iram_25 ) : ( n2888 ) ;
assign n2890 =  ( n2429 ) ? ( iram_24 ) : ( n2889 ) ;
assign n2891 =  ( n2428 ) ? ( iram_23 ) : ( n2890 ) ;
assign n2892 =  ( n2427 ) ? ( iram_22 ) : ( n2891 ) ;
assign n2893 =  ( n2426 ) ? ( iram_21 ) : ( n2892 ) ;
assign n2894 =  ( n2425 ) ? ( iram_20 ) : ( n2893 ) ;
assign n2895 =  ( n2424 ) ? ( iram_19 ) : ( n2894 ) ;
assign n2896 =  ( n2423 ) ? ( iram_18 ) : ( n2895 ) ;
assign n2897 =  ( n2422 ) ? ( iram_17 ) : ( n2896 ) ;
assign n2898 =  ( n2421 ) ? ( iram_16 ) : ( n2897 ) ;
assign n2899 =  ( n2420 ) ? ( iram_15 ) : ( n2898 ) ;
assign n2900 =  ( n2419 ) ? ( iram_14 ) : ( n2899 ) ;
assign n2901 =  ( n2418 ) ? ( iram_13 ) : ( n2900 ) ;
assign n2902 =  ( n2417 ) ? ( iram_12 ) : ( n2901 ) ;
assign n2903 =  ( n2416 ) ? ( iram_11 ) : ( n2902 ) ;
assign n2904 =  ( n2415 ) ? ( iram_10 ) : ( n2903 ) ;
assign n2905 =  ( n2414 ) ? ( iram_9 ) : ( n2904 ) ;
assign n2906 =  ( n2413 ) ? ( iram_8 ) : ( n2905 ) ;
assign n2907 =  ( n2412 ) ? ( iram_7 ) : ( n2906 ) ;
assign n2908 =  ( n2411 ) ? ( iram_6 ) : ( n2907 ) ;
assign n2909 =  ( n2410 ) ? ( iram_5 ) : ( n2908 ) ;
assign n2910 =  ( n2409 ) ? ( iram_4 ) : ( n2909 ) ;
assign n2911 =  ( n2408 ) ? ( iram_3 ) : ( n2910 ) ;
assign n2912 =  ( n2407 ) ? ( iram_2 ) : ( n2911 ) ;
assign n2913 =  ( n2406 ) ? ( iram_1 ) : ( n2912 ) ;
assign n2914 =  ( n2405 ) ? ( iram_0 ) : ( n2913 ) ;
assign n2915 =  ( n2403 ) ? ( ram_rd_data ) : ( n2914 ) ;
assign n2916 = rd_addr[7:7] ;
assign n2917 =  ( n2916 ) == ( bv_1_1_n34 )  ;
assign n2918 = rd_addr[6:3] ;
assign n2919 =  { ( bv_1_1_n34 ) , ( n2918 ) }  ;
assign n2920 =  { ( n2919 ) , ( bv_3_0_n46 ) }  ;
assign n2921 = rd_addr[6:3] ;
assign n2922 =  { ( bv_4_2_n12 ) , ( n2921 ) }  ;
assign n2923 =  ( n2917 ) ? ( n2920 ) : ( n2922 ) ;
assign n2924 =  ( bit_addr ) ? ( n2923 ) : ( rd_addr ) ;
assign n2925 =  ( n2924 ) == ( n51 )  ;
assign n2926 = n2924[7:0] ;
assign n2927 =  ( n2926 ) == ( bv_8_0_n69 )  ;
assign n2928 =  ( n2926 ) == ( bv_8_1_n71 )  ;
assign n2929 =  ( n2926 ) == ( bv_8_2_n73 )  ;
assign n2930 =  ( n2926 ) == ( bv_8_3_n75 )  ;
assign n2931 =  ( n2926 ) == ( bv_8_4_n77 )  ;
assign n2932 =  ( n2926 ) == ( bv_8_5_n79 )  ;
assign n2933 =  ( n2926 ) == ( bv_8_6_n81 )  ;
assign n2934 =  ( n2926 ) == ( bv_8_7_n83 )  ;
assign n2935 =  ( n2926 ) == ( bv_8_8_n85 )  ;
assign n2936 =  ( n2926 ) == ( bv_8_9_n87 )  ;
assign n2937 =  ( n2926 ) == ( bv_8_10_n89 )  ;
assign n2938 =  ( n2926 ) == ( bv_8_11_n91 )  ;
assign n2939 =  ( n2926 ) == ( bv_8_12_n93 )  ;
assign n2940 =  ( n2926 ) == ( bv_8_13_n95 )  ;
assign n2941 =  ( n2926 ) == ( bv_8_14_n97 )  ;
assign n2942 =  ( n2926 ) == ( bv_8_15_n99 )  ;
assign n2943 =  ( n2926 ) == ( bv_8_16_n101 )  ;
assign n2944 =  ( n2926 ) == ( bv_8_17_n103 )  ;
assign n2945 =  ( n2926 ) == ( bv_8_18_n105 )  ;
assign n2946 =  ( n2926 ) == ( bv_8_19_n107 )  ;
assign n2947 =  ( n2926 ) == ( bv_8_20_n109 )  ;
assign n2948 =  ( n2926 ) == ( bv_8_21_n111 )  ;
assign n2949 =  ( n2926 ) == ( bv_8_22_n113 )  ;
assign n2950 =  ( n2926 ) == ( bv_8_23_n115 )  ;
assign n2951 =  ( n2926 ) == ( bv_8_24_n117 )  ;
assign n2952 =  ( n2926 ) == ( bv_8_25_n119 )  ;
assign n2953 =  ( n2926 ) == ( bv_8_26_n121 )  ;
assign n2954 =  ( n2926 ) == ( bv_8_27_n123 )  ;
assign n2955 =  ( n2926 ) == ( bv_8_28_n125 )  ;
assign n2956 =  ( n2926 ) == ( bv_8_29_n127 )  ;
assign n2957 =  ( n2926 ) == ( bv_8_30_n129 )  ;
assign n2958 =  ( n2926 ) == ( bv_8_31_n131 )  ;
assign n2959 =  ( n2926 ) == ( bv_8_32_n133 )  ;
assign n2960 =  ( n2926 ) == ( bv_8_33_n135 )  ;
assign n2961 =  ( n2926 ) == ( bv_8_34_n137 )  ;
assign n2962 =  ( n2926 ) == ( bv_8_35_n139 )  ;
assign n2963 =  ( n2926 ) == ( bv_8_36_n141 )  ;
assign n2964 =  ( n2926 ) == ( bv_8_37_n143 )  ;
assign n2965 =  ( n2926 ) == ( bv_8_38_n145 )  ;
assign n2966 =  ( n2926 ) == ( bv_8_39_n147 )  ;
assign n2967 =  ( n2926 ) == ( bv_8_40_n149 )  ;
assign n2968 =  ( n2926 ) == ( bv_8_41_n151 )  ;
assign n2969 =  ( n2926 ) == ( bv_8_42_n153 )  ;
assign n2970 =  ( n2926 ) == ( bv_8_43_n155 )  ;
assign n2971 =  ( n2926 ) == ( bv_8_44_n157 )  ;
assign n2972 =  ( n2926 ) == ( bv_8_45_n159 )  ;
assign n2973 =  ( n2926 ) == ( bv_8_46_n161 )  ;
assign n2974 =  ( n2926 ) == ( bv_8_47_n163 )  ;
assign n2975 =  ( n2926 ) == ( bv_8_48_n165 )  ;
assign n2976 =  ( n2926 ) == ( bv_8_49_n167 )  ;
assign n2977 =  ( n2926 ) == ( bv_8_50_n169 )  ;
assign n2978 =  ( n2926 ) == ( bv_8_51_n171 )  ;
assign n2979 =  ( n2926 ) == ( bv_8_52_n173 )  ;
assign n2980 =  ( n2926 ) == ( bv_8_53_n175 )  ;
assign n2981 =  ( n2926 ) == ( bv_8_54_n177 )  ;
assign n2982 =  ( n2926 ) == ( bv_8_55_n179 )  ;
assign n2983 =  ( n2926 ) == ( bv_8_56_n181 )  ;
assign n2984 =  ( n2926 ) == ( bv_8_57_n183 )  ;
assign n2985 =  ( n2926 ) == ( bv_8_58_n185 )  ;
assign n2986 =  ( n2926 ) == ( bv_8_59_n187 )  ;
assign n2987 =  ( n2926 ) == ( bv_8_60_n189 )  ;
assign n2988 =  ( n2926 ) == ( bv_8_61_n191 )  ;
assign n2989 =  ( n2926 ) == ( bv_8_62_n193 )  ;
assign n2990 =  ( n2926 ) == ( bv_8_63_n195 )  ;
assign n2991 =  ( n2926 ) == ( bv_8_64_n197 )  ;
assign n2992 =  ( n2926 ) == ( bv_8_65_n199 )  ;
assign n2993 =  ( n2926 ) == ( bv_8_66_n201 )  ;
assign n2994 =  ( n2926 ) == ( bv_8_67_n203 )  ;
assign n2995 =  ( n2926 ) == ( bv_8_68_n205 )  ;
assign n2996 =  ( n2926 ) == ( bv_8_69_n207 )  ;
assign n2997 =  ( n2926 ) == ( bv_8_70_n209 )  ;
assign n2998 =  ( n2926 ) == ( bv_8_71_n211 )  ;
assign n2999 =  ( n2926 ) == ( bv_8_72_n213 )  ;
assign n3000 =  ( n2926 ) == ( bv_8_73_n215 )  ;
assign n3001 =  ( n2926 ) == ( bv_8_74_n217 )  ;
assign n3002 =  ( n2926 ) == ( bv_8_75_n219 )  ;
assign n3003 =  ( n2926 ) == ( bv_8_76_n221 )  ;
assign n3004 =  ( n2926 ) == ( bv_8_77_n223 )  ;
assign n3005 =  ( n2926 ) == ( bv_8_78_n225 )  ;
assign n3006 =  ( n2926 ) == ( bv_8_79_n227 )  ;
assign n3007 =  ( n2926 ) == ( bv_8_80_n229 )  ;
assign n3008 =  ( n2926 ) == ( bv_8_81_n231 )  ;
assign n3009 =  ( n2926 ) == ( bv_8_82_n233 )  ;
assign n3010 =  ( n2926 ) == ( bv_8_83_n235 )  ;
assign n3011 =  ( n2926 ) == ( bv_8_84_n237 )  ;
assign n3012 =  ( n2926 ) == ( bv_8_85_n239 )  ;
assign n3013 =  ( n2926 ) == ( bv_8_86_n241 )  ;
assign n3014 =  ( n2926 ) == ( bv_8_87_n243 )  ;
assign n3015 =  ( n2926 ) == ( bv_8_88_n245 )  ;
assign n3016 =  ( n2926 ) == ( bv_8_89_n247 )  ;
assign n3017 =  ( n2926 ) == ( bv_8_90_n249 )  ;
assign n3018 =  ( n2926 ) == ( bv_8_91_n251 )  ;
assign n3019 =  ( n2926 ) == ( bv_8_92_n253 )  ;
assign n3020 =  ( n2926 ) == ( bv_8_93_n255 )  ;
assign n3021 =  ( n2926 ) == ( bv_8_94_n257 )  ;
assign n3022 =  ( n2926 ) == ( bv_8_95_n259 )  ;
assign n3023 =  ( n2926 ) == ( bv_8_96_n261 )  ;
assign n3024 =  ( n2926 ) == ( bv_8_97_n263 )  ;
assign n3025 =  ( n2926 ) == ( bv_8_98_n265 )  ;
assign n3026 =  ( n2926 ) == ( bv_8_99_n267 )  ;
assign n3027 =  ( n2926 ) == ( bv_8_100_n269 )  ;
assign n3028 =  ( n2926 ) == ( bv_8_101_n271 )  ;
assign n3029 =  ( n2926 ) == ( bv_8_102_n273 )  ;
assign n3030 =  ( n2926 ) == ( bv_8_103_n275 )  ;
assign n3031 =  ( n2926 ) == ( bv_8_104_n277 )  ;
assign n3032 =  ( n2926 ) == ( bv_8_105_n279 )  ;
assign n3033 =  ( n2926 ) == ( bv_8_106_n281 )  ;
assign n3034 =  ( n2926 ) == ( bv_8_107_n283 )  ;
assign n3035 =  ( n2926 ) == ( bv_8_108_n285 )  ;
assign n3036 =  ( n2926 ) == ( bv_8_109_n287 )  ;
assign n3037 =  ( n2926 ) == ( bv_8_110_n289 )  ;
assign n3038 =  ( n2926 ) == ( bv_8_111_n291 )  ;
assign n3039 =  ( n2926 ) == ( bv_8_112_n293 )  ;
assign n3040 =  ( n2926 ) == ( bv_8_113_n295 )  ;
assign n3041 =  ( n2926 ) == ( bv_8_114_n297 )  ;
assign n3042 =  ( n2926 ) == ( bv_8_115_n299 )  ;
assign n3043 =  ( n2926 ) == ( bv_8_116_n301 )  ;
assign n3044 =  ( n2926 ) == ( bv_8_117_n303 )  ;
assign n3045 =  ( n2926 ) == ( bv_8_118_n305 )  ;
assign n3046 =  ( n2926 ) == ( bv_8_119_n307 )  ;
assign n3047 =  ( n2926 ) == ( bv_8_120_n309 )  ;
assign n3048 =  ( n2926 ) == ( bv_8_121_n311 )  ;
assign n3049 =  ( n2926 ) == ( bv_8_122_n313 )  ;
assign n3050 =  ( n2926 ) == ( bv_8_123_n315 )  ;
assign n3051 =  ( n2926 ) == ( bv_8_124_n317 )  ;
assign n3052 =  ( n2926 ) == ( bv_8_125_n319 )  ;
assign n3053 =  ( n2926 ) == ( bv_8_126_n321 )  ;
assign n3054 =  ( n2926 ) == ( bv_8_127_n323 )  ;
assign n3055 =  ( n2926 ) == ( bv_8_128_n325 )  ;
assign n3056 =  ( n2926 ) == ( bv_8_129_n327 )  ;
assign n3057 =  ( n2926 ) == ( bv_8_130_n329 )  ;
assign n3058 =  ( n2926 ) == ( bv_8_131_n331 )  ;
assign n3059 =  ( n2926 ) == ( bv_8_132_n333 )  ;
assign n3060 =  ( n2926 ) == ( bv_8_133_n335 )  ;
assign n3061 =  ( n2926 ) == ( bv_8_134_n337 )  ;
assign n3062 =  ( n2926 ) == ( bv_8_135_n339 )  ;
assign n3063 =  ( n2926 ) == ( bv_8_136_n341 )  ;
assign n3064 =  ( n2926 ) == ( bv_8_137_n343 )  ;
assign n3065 =  ( n2926 ) == ( bv_8_138_n345 )  ;
assign n3066 =  ( n2926 ) == ( bv_8_139_n347 )  ;
assign n3067 =  ( n2926 ) == ( bv_8_140_n349 )  ;
assign n3068 =  ( n2926 ) == ( bv_8_141_n351 )  ;
assign n3069 =  ( n2926 ) == ( bv_8_142_n353 )  ;
assign n3070 =  ( n2926 ) == ( bv_8_143_n355 )  ;
assign n3071 =  ( n2926 ) == ( bv_8_144_n357 )  ;
assign n3072 =  ( n2926 ) == ( bv_8_145_n359 )  ;
assign n3073 =  ( n2926 ) == ( bv_8_146_n361 )  ;
assign n3074 =  ( n2926 ) == ( bv_8_147_n363 )  ;
assign n3075 =  ( n2926 ) == ( bv_8_148_n365 )  ;
assign n3076 =  ( n2926 ) == ( bv_8_149_n367 )  ;
assign n3077 =  ( n2926 ) == ( bv_8_150_n369 )  ;
assign n3078 =  ( n2926 ) == ( bv_8_151_n371 )  ;
assign n3079 =  ( n2926 ) == ( bv_8_152_n373 )  ;
assign n3080 =  ( n2926 ) == ( bv_8_153_n375 )  ;
assign n3081 =  ( n2926 ) == ( bv_8_154_n377 )  ;
assign n3082 =  ( n2926 ) == ( bv_8_155_n379 )  ;
assign n3083 =  ( n2926 ) == ( bv_8_156_n381 )  ;
assign n3084 =  ( n2926 ) == ( bv_8_157_n383 )  ;
assign n3085 =  ( n2926 ) == ( bv_8_158_n385 )  ;
assign n3086 =  ( n2926 ) == ( bv_8_159_n387 )  ;
assign n3087 =  ( n2926 ) == ( bv_8_160_n389 )  ;
assign n3088 =  ( n2926 ) == ( bv_8_161_n391 )  ;
assign n3089 =  ( n2926 ) == ( bv_8_162_n393 )  ;
assign n3090 =  ( n2926 ) == ( bv_8_163_n395 )  ;
assign n3091 =  ( n2926 ) == ( bv_8_164_n397 )  ;
assign n3092 =  ( n2926 ) == ( bv_8_165_n399 )  ;
assign n3093 =  ( n2926 ) == ( bv_8_166_n401 )  ;
assign n3094 =  ( n2926 ) == ( bv_8_167_n403 )  ;
assign n3095 =  ( n2926 ) == ( bv_8_168_n405 )  ;
assign n3096 =  ( n2926 ) == ( bv_8_169_n407 )  ;
assign n3097 =  ( n2926 ) == ( bv_8_170_n409 )  ;
assign n3098 =  ( n2926 ) == ( bv_8_171_n411 )  ;
assign n3099 =  ( n2926 ) == ( bv_8_172_n413 )  ;
assign n3100 =  ( n2926 ) == ( bv_8_173_n415 )  ;
assign n3101 =  ( n2926 ) == ( bv_8_174_n417 )  ;
assign n3102 =  ( n2926 ) == ( bv_8_175_n419 )  ;
assign n3103 =  ( n2926 ) == ( bv_8_176_n421 )  ;
assign n3104 =  ( n2926 ) == ( bv_8_177_n423 )  ;
assign n3105 =  ( n2926 ) == ( bv_8_178_n425 )  ;
assign n3106 =  ( n2926 ) == ( bv_8_179_n427 )  ;
assign n3107 =  ( n2926 ) == ( bv_8_180_n429 )  ;
assign n3108 =  ( n2926 ) == ( bv_8_181_n431 )  ;
assign n3109 =  ( n2926 ) == ( bv_8_182_n433 )  ;
assign n3110 =  ( n2926 ) == ( bv_8_183_n435 )  ;
assign n3111 =  ( n2926 ) == ( bv_8_184_n437 )  ;
assign n3112 =  ( n2926 ) == ( bv_8_185_n439 )  ;
assign n3113 =  ( n2926 ) == ( bv_8_186_n441 )  ;
assign n3114 =  ( n2926 ) == ( bv_8_187_n443 )  ;
assign n3115 =  ( n2926 ) == ( bv_8_188_n445 )  ;
assign n3116 =  ( n2926 ) == ( bv_8_189_n447 )  ;
assign n3117 =  ( n2926 ) == ( bv_8_190_n449 )  ;
assign n3118 =  ( n2926 ) == ( bv_8_191_n451 )  ;
assign n3119 =  ( n2926 ) == ( bv_8_192_n453 )  ;
assign n3120 =  ( n2926 ) == ( bv_8_193_n455 )  ;
assign n3121 =  ( n2926 ) == ( bv_8_194_n457 )  ;
assign n3122 =  ( n2926 ) == ( bv_8_195_n459 )  ;
assign n3123 =  ( n2926 ) == ( bv_8_196_n461 )  ;
assign n3124 =  ( n2926 ) == ( bv_8_197_n463 )  ;
assign n3125 =  ( n2926 ) == ( bv_8_198_n465 )  ;
assign n3126 =  ( n2926 ) == ( bv_8_199_n467 )  ;
assign n3127 =  ( n2926 ) == ( bv_8_200_n469 )  ;
assign n3128 =  ( n2926 ) == ( bv_8_201_n471 )  ;
assign n3129 =  ( n2926 ) == ( bv_8_202_n473 )  ;
assign n3130 =  ( n2926 ) == ( bv_8_203_n475 )  ;
assign n3131 =  ( n2926 ) == ( bv_8_204_n477 )  ;
assign n3132 =  ( n2926 ) == ( bv_8_205_n479 )  ;
assign n3133 =  ( n2926 ) == ( bv_8_206_n481 )  ;
assign n3134 =  ( n2926 ) == ( bv_8_207_n483 )  ;
assign n3135 =  ( n2926 ) == ( bv_8_208_n485 )  ;
assign n3136 =  ( n2926 ) == ( bv_8_209_n487 )  ;
assign n3137 =  ( n2926 ) == ( bv_8_210_n489 )  ;
assign n3138 =  ( n2926 ) == ( bv_8_211_n491 )  ;
assign n3139 =  ( n2926 ) == ( bv_8_212_n493 )  ;
assign n3140 =  ( n2926 ) == ( bv_8_213_n495 )  ;
assign n3141 =  ( n2926 ) == ( bv_8_214_n497 )  ;
assign n3142 =  ( n2926 ) == ( bv_8_215_n499 )  ;
assign n3143 =  ( n2926 ) == ( bv_8_216_n501 )  ;
assign n3144 =  ( n2926 ) == ( bv_8_217_n503 )  ;
assign n3145 =  ( n2926 ) == ( bv_8_218_n505 )  ;
assign n3146 =  ( n2926 ) == ( bv_8_219_n507 )  ;
assign n3147 =  ( n2926 ) == ( bv_8_220_n509 )  ;
assign n3148 =  ( n2926 ) == ( bv_8_221_n511 )  ;
assign n3149 =  ( n2926 ) == ( bv_8_222_n513 )  ;
assign n3150 =  ( n2926 ) == ( bv_8_223_n515 )  ;
assign n3151 =  ( n2926 ) == ( bv_8_224_n517 )  ;
assign n3152 =  ( n2926 ) == ( bv_8_225_n519 )  ;
assign n3153 =  ( n2926 ) == ( bv_8_226_n521 )  ;
assign n3154 =  ( n2926 ) == ( bv_8_227_n523 )  ;
assign n3155 =  ( n2926 ) == ( bv_8_228_n525 )  ;
assign n3156 =  ( n2926 ) == ( bv_8_229_n527 )  ;
assign n3157 =  ( n2926 ) == ( bv_8_230_n529 )  ;
assign n3158 =  ( n2926 ) == ( bv_8_231_n531 )  ;
assign n3159 =  ( n2926 ) == ( bv_8_232_n533 )  ;
assign n3160 =  ( n2926 ) == ( bv_8_233_n535 )  ;
assign n3161 =  ( n2926 ) == ( bv_8_234_n537 )  ;
assign n3162 =  ( n2926 ) == ( bv_8_235_n539 )  ;
assign n3163 =  ( n2926 ) == ( bv_8_236_n541 )  ;
assign n3164 =  ( n2926 ) == ( bv_8_237_n543 )  ;
assign n3165 =  ( n2926 ) == ( bv_8_238_n545 )  ;
assign n3166 =  ( n2926 ) == ( bv_8_239_n547 )  ;
assign n3167 =  ( n2926 ) == ( bv_8_240_n549 )  ;
assign n3168 =  ( n2926 ) == ( bv_8_241_n551 )  ;
assign n3169 =  ( n2926 ) == ( bv_8_242_n553 )  ;
assign n3170 =  ( n2926 ) == ( bv_8_243_n555 )  ;
assign n3171 =  ( n2926 ) == ( bv_8_244_n557 )  ;
assign n3172 =  ( n2926 ) == ( bv_8_245_n559 )  ;
assign n3173 =  ( n2926 ) == ( bv_8_246_n561 )  ;
assign n3174 =  ( n2926 ) == ( bv_8_247_n563 )  ;
assign n3175 =  ( n2926 ) == ( bv_8_248_n565 )  ;
assign n3176 =  ( n2926 ) == ( bv_8_249_n567 )  ;
assign n3177 =  ( n2926 ) == ( bv_8_250_n569 )  ;
assign n3178 =  ( n2926 ) == ( bv_8_251_n571 )  ;
assign n3179 =  ( n2926 ) == ( bv_8_252_n573 )  ;
assign n3180 =  ( n2926 ) == ( bv_8_253_n575 )  ;
assign n3181 =  ( n2926 ) == ( bv_8_254_n577 )  ;
assign n3182 =  ( n3181 ) ? ( iram_254 ) : ( iram_255 ) ;
assign n3183 =  ( n3180 ) ? ( iram_253 ) : ( n3182 ) ;
assign n3184 =  ( n3179 ) ? ( iram_252 ) : ( n3183 ) ;
assign n3185 =  ( n3178 ) ? ( iram_251 ) : ( n3184 ) ;
assign n3186 =  ( n3177 ) ? ( iram_250 ) : ( n3185 ) ;
assign n3187 =  ( n3176 ) ? ( iram_249 ) : ( n3186 ) ;
assign n3188 =  ( n3175 ) ? ( iram_248 ) : ( n3187 ) ;
assign n3189 =  ( n3174 ) ? ( iram_247 ) : ( n3188 ) ;
assign n3190 =  ( n3173 ) ? ( iram_246 ) : ( n3189 ) ;
assign n3191 =  ( n3172 ) ? ( iram_245 ) : ( n3190 ) ;
assign n3192 =  ( n3171 ) ? ( iram_244 ) : ( n3191 ) ;
assign n3193 =  ( n3170 ) ? ( iram_243 ) : ( n3192 ) ;
assign n3194 =  ( n3169 ) ? ( iram_242 ) : ( n3193 ) ;
assign n3195 =  ( n3168 ) ? ( iram_241 ) : ( n3194 ) ;
assign n3196 =  ( n3167 ) ? ( iram_240 ) : ( n3195 ) ;
assign n3197 =  ( n3166 ) ? ( iram_239 ) : ( n3196 ) ;
assign n3198 =  ( n3165 ) ? ( iram_238 ) : ( n3197 ) ;
assign n3199 =  ( n3164 ) ? ( iram_237 ) : ( n3198 ) ;
assign n3200 =  ( n3163 ) ? ( iram_236 ) : ( n3199 ) ;
assign n3201 =  ( n3162 ) ? ( iram_235 ) : ( n3200 ) ;
assign n3202 =  ( n3161 ) ? ( iram_234 ) : ( n3201 ) ;
assign n3203 =  ( n3160 ) ? ( iram_233 ) : ( n3202 ) ;
assign n3204 =  ( n3159 ) ? ( iram_232 ) : ( n3203 ) ;
assign n3205 =  ( n3158 ) ? ( iram_231 ) : ( n3204 ) ;
assign n3206 =  ( n3157 ) ? ( iram_230 ) : ( n3205 ) ;
assign n3207 =  ( n3156 ) ? ( iram_229 ) : ( n3206 ) ;
assign n3208 =  ( n3155 ) ? ( iram_228 ) : ( n3207 ) ;
assign n3209 =  ( n3154 ) ? ( iram_227 ) : ( n3208 ) ;
assign n3210 =  ( n3153 ) ? ( iram_226 ) : ( n3209 ) ;
assign n3211 =  ( n3152 ) ? ( iram_225 ) : ( n3210 ) ;
assign n3212 =  ( n3151 ) ? ( iram_224 ) : ( n3211 ) ;
assign n3213 =  ( n3150 ) ? ( iram_223 ) : ( n3212 ) ;
assign n3214 =  ( n3149 ) ? ( iram_222 ) : ( n3213 ) ;
assign n3215 =  ( n3148 ) ? ( iram_221 ) : ( n3214 ) ;
assign n3216 =  ( n3147 ) ? ( iram_220 ) : ( n3215 ) ;
assign n3217 =  ( n3146 ) ? ( iram_219 ) : ( n3216 ) ;
assign n3218 =  ( n3145 ) ? ( iram_218 ) : ( n3217 ) ;
assign n3219 =  ( n3144 ) ? ( iram_217 ) : ( n3218 ) ;
assign n3220 =  ( n3143 ) ? ( iram_216 ) : ( n3219 ) ;
assign n3221 =  ( n3142 ) ? ( iram_215 ) : ( n3220 ) ;
assign n3222 =  ( n3141 ) ? ( iram_214 ) : ( n3221 ) ;
assign n3223 =  ( n3140 ) ? ( iram_213 ) : ( n3222 ) ;
assign n3224 =  ( n3139 ) ? ( iram_212 ) : ( n3223 ) ;
assign n3225 =  ( n3138 ) ? ( iram_211 ) : ( n3224 ) ;
assign n3226 =  ( n3137 ) ? ( iram_210 ) : ( n3225 ) ;
assign n3227 =  ( n3136 ) ? ( iram_209 ) : ( n3226 ) ;
assign n3228 =  ( n3135 ) ? ( iram_208 ) : ( n3227 ) ;
assign n3229 =  ( n3134 ) ? ( iram_207 ) : ( n3228 ) ;
assign n3230 =  ( n3133 ) ? ( iram_206 ) : ( n3229 ) ;
assign n3231 =  ( n3132 ) ? ( iram_205 ) : ( n3230 ) ;
assign n3232 =  ( n3131 ) ? ( iram_204 ) : ( n3231 ) ;
assign n3233 =  ( n3130 ) ? ( iram_203 ) : ( n3232 ) ;
assign n3234 =  ( n3129 ) ? ( iram_202 ) : ( n3233 ) ;
assign n3235 =  ( n3128 ) ? ( iram_201 ) : ( n3234 ) ;
assign n3236 =  ( n3127 ) ? ( iram_200 ) : ( n3235 ) ;
assign n3237 =  ( n3126 ) ? ( iram_199 ) : ( n3236 ) ;
assign n3238 =  ( n3125 ) ? ( iram_198 ) : ( n3237 ) ;
assign n3239 =  ( n3124 ) ? ( iram_197 ) : ( n3238 ) ;
assign n3240 =  ( n3123 ) ? ( iram_196 ) : ( n3239 ) ;
assign n3241 =  ( n3122 ) ? ( iram_195 ) : ( n3240 ) ;
assign n3242 =  ( n3121 ) ? ( iram_194 ) : ( n3241 ) ;
assign n3243 =  ( n3120 ) ? ( iram_193 ) : ( n3242 ) ;
assign n3244 =  ( n3119 ) ? ( iram_192 ) : ( n3243 ) ;
assign n3245 =  ( n3118 ) ? ( iram_191 ) : ( n3244 ) ;
assign n3246 =  ( n3117 ) ? ( iram_190 ) : ( n3245 ) ;
assign n3247 =  ( n3116 ) ? ( iram_189 ) : ( n3246 ) ;
assign n3248 =  ( n3115 ) ? ( iram_188 ) : ( n3247 ) ;
assign n3249 =  ( n3114 ) ? ( iram_187 ) : ( n3248 ) ;
assign n3250 =  ( n3113 ) ? ( iram_186 ) : ( n3249 ) ;
assign n3251 =  ( n3112 ) ? ( iram_185 ) : ( n3250 ) ;
assign n3252 =  ( n3111 ) ? ( iram_184 ) : ( n3251 ) ;
assign n3253 =  ( n3110 ) ? ( iram_183 ) : ( n3252 ) ;
assign n3254 =  ( n3109 ) ? ( iram_182 ) : ( n3253 ) ;
assign n3255 =  ( n3108 ) ? ( iram_181 ) : ( n3254 ) ;
assign n3256 =  ( n3107 ) ? ( iram_180 ) : ( n3255 ) ;
assign n3257 =  ( n3106 ) ? ( iram_179 ) : ( n3256 ) ;
assign n3258 =  ( n3105 ) ? ( iram_178 ) : ( n3257 ) ;
assign n3259 =  ( n3104 ) ? ( iram_177 ) : ( n3258 ) ;
assign n3260 =  ( n3103 ) ? ( iram_176 ) : ( n3259 ) ;
assign n3261 =  ( n3102 ) ? ( iram_175 ) : ( n3260 ) ;
assign n3262 =  ( n3101 ) ? ( iram_174 ) : ( n3261 ) ;
assign n3263 =  ( n3100 ) ? ( iram_173 ) : ( n3262 ) ;
assign n3264 =  ( n3099 ) ? ( iram_172 ) : ( n3263 ) ;
assign n3265 =  ( n3098 ) ? ( iram_171 ) : ( n3264 ) ;
assign n3266 =  ( n3097 ) ? ( iram_170 ) : ( n3265 ) ;
assign n3267 =  ( n3096 ) ? ( iram_169 ) : ( n3266 ) ;
assign n3268 =  ( n3095 ) ? ( iram_168 ) : ( n3267 ) ;
assign n3269 =  ( n3094 ) ? ( iram_167 ) : ( n3268 ) ;
assign n3270 =  ( n3093 ) ? ( iram_166 ) : ( n3269 ) ;
assign n3271 =  ( n3092 ) ? ( iram_165 ) : ( n3270 ) ;
assign n3272 =  ( n3091 ) ? ( iram_164 ) : ( n3271 ) ;
assign n3273 =  ( n3090 ) ? ( iram_163 ) : ( n3272 ) ;
assign n3274 =  ( n3089 ) ? ( iram_162 ) : ( n3273 ) ;
assign n3275 =  ( n3088 ) ? ( iram_161 ) : ( n3274 ) ;
assign n3276 =  ( n3087 ) ? ( iram_160 ) : ( n3275 ) ;
assign n3277 =  ( n3086 ) ? ( iram_159 ) : ( n3276 ) ;
assign n3278 =  ( n3085 ) ? ( iram_158 ) : ( n3277 ) ;
assign n3279 =  ( n3084 ) ? ( iram_157 ) : ( n3278 ) ;
assign n3280 =  ( n3083 ) ? ( iram_156 ) : ( n3279 ) ;
assign n3281 =  ( n3082 ) ? ( iram_155 ) : ( n3280 ) ;
assign n3282 =  ( n3081 ) ? ( iram_154 ) : ( n3281 ) ;
assign n3283 =  ( n3080 ) ? ( iram_153 ) : ( n3282 ) ;
assign n3284 =  ( n3079 ) ? ( iram_152 ) : ( n3283 ) ;
assign n3285 =  ( n3078 ) ? ( iram_151 ) : ( n3284 ) ;
assign n3286 =  ( n3077 ) ? ( iram_150 ) : ( n3285 ) ;
assign n3287 =  ( n3076 ) ? ( iram_149 ) : ( n3286 ) ;
assign n3288 =  ( n3075 ) ? ( iram_148 ) : ( n3287 ) ;
assign n3289 =  ( n3074 ) ? ( iram_147 ) : ( n3288 ) ;
assign n3290 =  ( n3073 ) ? ( iram_146 ) : ( n3289 ) ;
assign n3291 =  ( n3072 ) ? ( iram_145 ) : ( n3290 ) ;
assign n3292 =  ( n3071 ) ? ( iram_144 ) : ( n3291 ) ;
assign n3293 =  ( n3070 ) ? ( iram_143 ) : ( n3292 ) ;
assign n3294 =  ( n3069 ) ? ( iram_142 ) : ( n3293 ) ;
assign n3295 =  ( n3068 ) ? ( iram_141 ) : ( n3294 ) ;
assign n3296 =  ( n3067 ) ? ( iram_140 ) : ( n3295 ) ;
assign n3297 =  ( n3066 ) ? ( iram_139 ) : ( n3296 ) ;
assign n3298 =  ( n3065 ) ? ( iram_138 ) : ( n3297 ) ;
assign n3299 =  ( n3064 ) ? ( iram_137 ) : ( n3298 ) ;
assign n3300 =  ( n3063 ) ? ( iram_136 ) : ( n3299 ) ;
assign n3301 =  ( n3062 ) ? ( iram_135 ) : ( n3300 ) ;
assign n3302 =  ( n3061 ) ? ( iram_134 ) : ( n3301 ) ;
assign n3303 =  ( n3060 ) ? ( iram_133 ) : ( n3302 ) ;
assign n3304 =  ( n3059 ) ? ( iram_132 ) : ( n3303 ) ;
assign n3305 =  ( n3058 ) ? ( iram_131 ) : ( n3304 ) ;
assign n3306 =  ( n3057 ) ? ( iram_130 ) : ( n3305 ) ;
assign n3307 =  ( n3056 ) ? ( iram_129 ) : ( n3306 ) ;
assign n3308 =  ( n3055 ) ? ( iram_128 ) : ( n3307 ) ;
assign n3309 =  ( n3054 ) ? ( iram_127 ) : ( n3308 ) ;
assign n3310 =  ( n3053 ) ? ( iram_126 ) : ( n3309 ) ;
assign n3311 =  ( n3052 ) ? ( iram_125 ) : ( n3310 ) ;
assign n3312 =  ( n3051 ) ? ( iram_124 ) : ( n3311 ) ;
assign n3313 =  ( n3050 ) ? ( iram_123 ) : ( n3312 ) ;
assign n3314 =  ( n3049 ) ? ( iram_122 ) : ( n3313 ) ;
assign n3315 =  ( n3048 ) ? ( iram_121 ) : ( n3314 ) ;
assign n3316 =  ( n3047 ) ? ( iram_120 ) : ( n3315 ) ;
assign n3317 =  ( n3046 ) ? ( iram_119 ) : ( n3316 ) ;
assign n3318 =  ( n3045 ) ? ( iram_118 ) : ( n3317 ) ;
assign n3319 =  ( n3044 ) ? ( iram_117 ) : ( n3318 ) ;
assign n3320 =  ( n3043 ) ? ( iram_116 ) : ( n3319 ) ;
assign n3321 =  ( n3042 ) ? ( iram_115 ) : ( n3320 ) ;
assign n3322 =  ( n3041 ) ? ( iram_114 ) : ( n3321 ) ;
assign n3323 =  ( n3040 ) ? ( iram_113 ) : ( n3322 ) ;
assign n3324 =  ( n3039 ) ? ( iram_112 ) : ( n3323 ) ;
assign n3325 =  ( n3038 ) ? ( iram_111 ) : ( n3324 ) ;
assign n3326 =  ( n3037 ) ? ( iram_110 ) : ( n3325 ) ;
assign n3327 =  ( n3036 ) ? ( iram_109 ) : ( n3326 ) ;
assign n3328 =  ( n3035 ) ? ( iram_108 ) : ( n3327 ) ;
assign n3329 =  ( n3034 ) ? ( iram_107 ) : ( n3328 ) ;
assign n3330 =  ( n3033 ) ? ( iram_106 ) : ( n3329 ) ;
assign n3331 =  ( n3032 ) ? ( iram_105 ) : ( n3330 ) ;
assign n3332 =  ( n3031 ) ? ( iram_104 ) : ( n3331 ) ;
assign n3333 =  ( n3030 ) ? ( iram_103 ) : ( n3332 ) ;
assign n3334 =  ( n3029 ) ? ( iram_102 ) : ( n3333 ) ;
assign n3335 =  ( n3028 ) ? ( iram_101 ) : ( n3334 ) ;
assign n3336 =  ( n3027 ) ? ( iram_100 ) : ( n3335 ) ;
assign n3337 =  ( n3026 ) ? ( iram_99 ) : ( n3336 ) ;
assign n3338 =  ( n3025 ) ? ( iram_98 ) : ( n3337 ) ;
assign n3339 =  ( n3024 ) ? ( iram_97 ) : ( n3338 ) ;
assign n3340 =  ( n3023 ) ? ( iram_96 ) : ( n3339 ) ;
assign n3341 =  ( n3022 ) ? ( iram_95 ) : ( n3340 ) ;
assign n3342 =  ( n3021 ) ? ( iram_94 ) : ( n3341 ) ;
assign n3343 =  ( n3020 ) ? ( iram_93 ) : ( n3342 ) ;
assign n3344 =  ( n3019 ) ? ( iram_92 ) : ( n3343 ) ;
assign n3345 =  ( n3018 ) ? ( iram_91 ) : ( n3344 ) ;
assign n3346 =  ( n3017 ) ? ( iram_90 ) : ( n3345 ) ;
assign n3347 =  ( n3016 ) ? ( iram_89 ) : ( n3346 ) ;
assign n3348 =  ( n3015 ) ? ( iram_88 ) : ( n3347 ) ;
assign n3349 =  ( n3014 ) ? ( iram_87 ) : ( n3348 ) ;
assign n3350 =  ( n3013 ) ? ( iram_86 ) : ( n3349 ) ;
assign n3351 =  ( n3012 ) ? ( iram_85 ) : ( n3350 ) ;
assign n3352 =  ( n3011 ) ? ( iram_84 ) : ( n3351 ) ;
assign n3353 =  ( n3010 ) ? ( iram_83 ) : ( n3352 ) ;
assign n3354 =  ( n3009 ) ? ( iram_82 ) : ( n3353 ) ;
assign n3355 =  ( n3008 ) ? ( iram_81 ) : ( n3354 ) ;
assign n3356 =  ( n3007 ) ? ( iram_80 ) : ( n3355 ) ;
assign n3357 =  ( n3006 ) ? ( iram_79 ) : ( n3356 ) ;
assign n3358 =  ( n3005 ) ? ( iram_78 ) : ( n3357 ) ;
assign n3359 =  ( n3004 ) ? ( iram_77 ) : ( n3358 ) ;
assign n3360 =  ( n3003 ) ? ( iram_76 ) : ( n3359 ) ;
assign n3361 =  ( n3002 ) ? ( iram_75 ) : ( n3360 ) ;
assign n3362 =  ( n3001 ) ? ( iram_74 ) : ( n3361 ) ;
assign n3363 =  ( n3000 ) ? ( iram_73 ) : ( n3362 ) ;
assign n3364 =  ( n2999 ) ? ( iram_72 ) : ( n3363 ) ;
assign n3365 =  ( n2998 ) ? ( iram_71 ) : ( n3364 ) ;
assign n3366 =  ( n2997 ) ? ( iram_70 ) : ( n3365 ) ;
assign n3367 =  ( n2996 ) ? ( iram_69 ) : ( n3366 ) ;
assign n3368 =  ( n2995 ) ? ( iram_68 ) : ( n3367 ) ;
assign n3369 =  ( n2994 ) ? ( iram_67 ) : ( n3368 ) ;
assign n3370 =  ( n2993 ) ? ( iram_66 ) : ( n3369 ) ;
assign n3371 =  ( n2992 ) ? ( iram_65 ) : ( n3370 ) ;
assign n3372 =  ( n2991 ) ? ( iram_64 ) : ( n3371 ) ;
assign n3373 =  ( n2990 ) ? ( iram_63 ) : ( n3372 ) ;
assign n3374 =  ( n2989 ) ? ( iram_62 ) : ( n3373 ) ;
assign n3375 =  ( n2988 ) ? ( iram_61 ) : ( n3374 ) ;
assign n3376 =  ( n2987 ) ? ( iram_60 ) : ( n3375 ) ;
assign n3377 =  ( n2986 ) ? ( iram_59 ) : ( n3376 ) ;
assign n3378 =  ( n2985 ) ? ( iram_58 ) : ( n3377 ) ;
assign n3379 =  ( n2984 ) ? ( iram_57 ) : ( n3378 ) ;
assign n3380 =  ( n2983 ) ? ( iram_56 ) : ( n3379 ) ;
assign n3381 =  ( n2982 ) ? ( iram_55 ) : ( n3380 ) ;
assign n3382 =  ( n2981 ) ? ( iram_54 ) : ( n3381 ) ;
assign n3383 =  ( n2980 ) ? ( iram_53 ) : ( n3382 ) ;
assign n3384 =  ( n2979 ) ? ( iram_52 ) : ( n3383 ) ;
assign n3385 =  ( n2978 ) ? ( iram_51 ) : ( n3384 ) ;
assign n3386 =  ( n2977 ) ? ( iram_50 ) : ( n3385 ) ;
assign n3387 =  ( n2976 ) ? ( iram_49 ) : ( n3386 ) ;
assign n3388 =  ( n2975 ) ? ( iram_48 ) : ( n3387 ) ;
assign n3389 =  ( n2974 ) ? ( iram_47 ) : ( n3388 ) ;
assign n3390 =  ( n2973 ) ? ( iram_46 ) : ( n3389 ) ;
assign n3391 =  ( n2972 ) ? ( iram_45 ) : ( n3390 ) ;
assign n3392 =  ( n2971 ) ? ( iram_44 ) : ( n3391 ) ;
assign n3393 =  ( n2970 ) ? ( iram_43 ) : ( n3392 ) ;
assign n3394 =  ( n2969 ) ? ( iram_42 ) : ( n3393 ) ;
assign n3395 =  ( n2968 ) ? ( iram_41 ) : ( n3394 ) ;
assign n3396 =  ( n2967 ) ? ( iram_40 ) : ( n3395 ) ;
assign n3397 =  ( n2966 ) ? ( iram_39 ) : ( n3396 ) ;
assign n3398 =  ( n2965 ) ? ( iram_38 ) : ( n3397 ) ;
assign n3399 =  ( n2964 ) ? ( iram_37 ) : ( n3398 ) ;
assign n3400 =  ( n2963 ) ? ( iram_36 ) : ( n3399 ) ;
assign n3401 =  ( n2962 ) ? ( iram_35 ) : ( n3400 ) ;
assign n3402 =  ( n2961 ) ? ( iram_34 ) : ( n3401 ) ;
assign n3403 =  ( n2960 ) ? ( iram_33 ) : ( n3402 ) ;
assign n3404 =  ( n2959 ) ? ( iram_32 ) : ( n3403 ) ;
assign n3405 =  ( n2958 ) ? ( iram_31 ) : ( n3404 ) ;
assign n3406 =  ( n2957 ) ? ( iram_30 ) : ( n3405 ) ;
assign n3407 =  ( n2956 ) ? ( iram_29 ) : ( n3406 ) ;
assign n3408 =  ( n2955 ) ? ( iram_28 ) : ( n3407 ) ;
assign n3409 =  ( n2954 ) ? ( iram_27 ) : ( n3408 ) ;
assign n3410 =  ( n2953 ) ? ( iram_26 ) : ( n3409 ) ;
assign n3411 =  ( n2952 ) ? ( iram_25 ) : ( n3410 ) ;
assign n3412 =  ( n2951 ) ? ( iram_24 ) : ( n3411 ) ;
assign n3413 =  ( n2950 ) ? ( iram_23 ) : ( n3412 ) ;
assign n3414 =  ( n2949 ) ? ( iram_22 ) : ( n3413 ) ;
assign n3415 =  ( n2948 ) ? ( iram_21 ) : ( n3414 ) ;
assign n3416 =  ( n2947 ) ? ( iram_20 ) : ( n3415 ) ;
assign n3417 =  ( n2946 ) ? ( iram_19 ) : ( n3416 ) ;
assign n3418 =  ( n2945 ) ? ( iram_18 ) : ( n3417 ) ;
assign n3419 =  ( n2944 ) ? ( iram_17 ) : ( n3418 ) ;
assign n3420 =  ( n2943 ) ? ( iram_16 ) : ( n3419 ) ;
assign n3421 =  ( n2942 ) ? ( iram_15 ) : ( n3420 ) ;
assign n3422 =  ( n2941 ) ? ( iram_14 ) : ( n3421 ) ;
assign n3423 =  ( n2940 ) ? ( iram_13 ) : ( n3422 ) ;
assign n3424 =  ( n2939 ) ? ( iram_12 ) : ( n3423 ) ;
assign n3425 =  ( n2938 ) ? ( iram_11 ) : ( n3424 ) ;
assign n3426 =  ( n2937 ) ? ( iram_10 ) : ( n3425 ) ;
assign n3427 =  ( n2936 ) ? ( iram_9 ) : ( n3426 ) ;
assign n3428 =  ( n2935 ) ? ( iram_8 ) : ( n3427 ) ;
assign n3429 =  ( n2934 ) ? ( iram_7 ) : ( n3428 ) ;
assign n3430 =  ( n2933 ) ? ( iram_6 ) : ( n3429 ) ;
assign n3431 =  ( n2932 ) ? ( iram_5 ) : ( n3430 ) ;
assign n3432 =  ( n2931 ) ? ( iram_4 ) : ( n3431 ) ;
assign n3433 =  ( n2930 ) ? ( iram_3 ) : ( n3432 ) ;
assign n3434 =  ( n2929 ) ? ( iram_2 ) : ( n3433 ) ;
assign n3435 =  ( n2928 ) ? ( iram_1 ) : ( n3434 ) ;
assign n3436 =  ( n2927 ) ? ( iram_0 ) : ( n3435 ) ;
assign n3437 =  ( n2925 ) ? ( ram_rd_data ) : ( n3436 ) ;
assign n3438 = rd_addr[7:3] ;
assign n3439 =  { ( n3438 ) , ( bv_3_0_n46 ) }  ;
assign n3440 =  ( n3439 ) == ( bv_8_224_n517 )  ;
assign n3441 =  ( n3439 ) == ( bv_8_240_n549 )  ;
assign n3442 =  ( n3439 ) == ( bv_8_208_n485 )  ;
assign n3443 =  { ( psw ) , ( p ) }  ;
assign n3444 =  ( n3439 ) == ( bv_8_129_n327 )  ;
assign n3445 =  ( n3439 ) == ( bv_8_130_n329 )  ;
assign n3446 =  ( n3439 ) == ( bv_8_131_n331 )  ;
assign n3447 =  ( n3439 ) == ( bv_8_128_n325 )  ;
assign n3448 =  ( n3439 ) == ( bv_8_144_n357 )  ;
assign n3449 =  ( n3439 ) == ( bv_8_160_n389 )  ;
assign n3450 =  ( n3439 ) == ( bv_8_176_n421 )  ;
assign n3451 =  ( n3439 ) == ( bv_8_184_n437 )  ;
assign n3452 =  ( n3439 ) == ( bv_8_168_n405 )  ;
assign n3453 =  ( n3439 ) == ( bv_8_136_n341 )  ;
assign n3454 =  ( n3439 ) == ( bv_8_152_n373 )  ;
assign n3455 =  ( n3454 ) ? ( scon ) : ( bv_8_0_n69 ) ;
assign n3456 =  ( n3453 ) ? ( tcon ) : ( n3455 ) ;
assign n3457 =  ( n3452 ) ? ( ie ) : ( n3456 ) ;
assign n3458 =  ( n3451 ) ? ( ip ) : ( n3457 ) ;
assign n3459 =  ( n3450 ) ? ( p3 ) : ( n3458 ) ;
assign n3460 =  ( n3449 ) ? ( p2 ) : ( n3459 ) ;
assign n3461 =  ( n3448 ) ? ( p1 ) : ( n3460 ) ;
assign n3462 =  ( n3447 ) ? ( p0 ) : ( n3461 ) ;
assign n3463 =  ( n3446 ) ? ( dptr_hi ) : ( n3462 ) ;
assign n3464 =  ( n3445 ) ? ( dptr_lo ) : ( n3463 ) ;
assign n3465 =  ( n3444 ) ? ( sp ) : ( n3464 ) ;
assign n3466 =  ( n3442 ) ? ( n3443 ) : ( n3465 ) ;
assign n3467 =  ( n3441 ) ? ( b_reg ) : ( n3466 ) ;
assign n3468 =  ( n3440 ) ? ( acc ) : ( n3467 ) ;
assign n3469 =  ( rd_addr ) == ( bv_8_224_n517 )  ;
assign n3470 =  ( rd_addr ) == ( bv_8_240_n549 )  ;
assign n3471 =  ( rd_addr ) == ( bv_8_208_n485 )  ;
assign n3472 =  { ( psw ) , ( p ) }  ;
assign n3473 =  ( rd_addr ) == ( bv_8_129_n327 )  ;
assign n3474 =  ( rd_addr ) == ( bv_8_130_n329 )  ;
assign n3475 =  ( rd_addr ) == ( bv_8_131_n331 )  ;
assign n3476 =  ( rd_addr ) == ( bv_8_128_n325 )  ;
assign n3477 =  ( rd_addr ) == ( bv_8_144_n357 )  ;
assign n3478 =  ( rd_addr ) == ( bv_8_160_n389 )  ;
assign n3479 =  ( rd_addr ) == ( bv_8_176_n421 )  ;
assign n3480 =  ( rd_addr ) == ( bv_8_184_n437 )  ;
assign n3481 =  ( rd_addr ) == ( bv_8_168_n405 )  ;
assign n3482 =  ( n3481 ) ? ( ie ) : ( bv_8_0_n69 ) ;
assign n3483 =  ( n3480 ) ? ( ip ) : ( n3482 ) ;
assign n3484 =  ( n3479 ) ? ( p3 ) : ( n3483 ) ;
assign n3485 =  ( n3478 ) ? ( p2 ) : ( n3484 ) ;
assign n3486 =  ( n3477 ) ? ( p1 ) : ( n3485 ) ;
assign n3487 =  ( n3476 ) ? ( p0 ) : ( n3486 ) ;
assign n3488 =  ( n3475 ) ? ( dptr_hi ) : ( n3487 ) ;
assign n3489 =  ( n3474 ) ? ( dptr_lo ) : ( n3488 ) ;
assign n3490 =  ( n3473 ) ? ( sp ) : ( n3489 ) ;
assign n3491 =  ( n3471 ) ? ( n3472 ) : ( n3490 ) ;
assign n3492 =  ( n3470 ) ? ( b_reg ) : ( n3491 ) ;
assign n3493 =  ( n3469 ) ? ( acc ) : ( n3492 ) ;
assign n3494 =  ( bit_addr ) ? ( n3468 ) : ( n3493 ) ;
assign bv_2_3_n3495 = 2'h3 ;
assign n3496 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n3497 =  ( rd_addr ) == ( bv_8_130_n329 )  ;
assign n3498 =  ( n3496 ) & (n3497 )  ;
assign n3500 = nondet_des_acc_func_n3499 ;
assign bv_2_1_n3501 = 2'h1 ;
assign n3502 =  ( wr_sfr ) == ( bv_2_1_n3501 )  ;
assign n3503 =  ( rd_addr ) == ( bv_8_224_n517 )  ;
assign n3504 =  ( n3502 ) & (n3503 )  ;
assign bv_2_2_n3505 = 2'h2 ;
assign n3506 =  ( wr_sfr ) == ( bv_2_2_n3505 )  ;
assign n3507 =  ( rd_addr ) == ( bv_8_224_n517 )  ;
assign n3508 =  ( n3506 ) & (n3507 )  ;
assign n3509 =  ( n3504 ) | ( n3508 )  ;
assign n3510 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n3511 =  ( rd_addr ) == ( bv_8_131_n331 )  ;
assign n3512 =  ( n3510 ) & (n3511 )  ;
assign n3513 =  ( n3509 ) | ( n3512 )  ;
assign n3514 =  ( wait_data ) == ( 1'b0 )  ;
assign n3515 =  ( n3513 ) & (n3514 )  ;
assign n3516 =  ( rd_addr ) == ( bv_8_129_n327 )  ;
assign bv_3_3_n3517 = 3'h3 ;
assign n3518 =  ( ram_wr_sel ) == ( bv_3_3_n3517 )  ;
assign n3519 =  ( sp ) + ( bv_8_1_n71 )  ;
assign bv_7_0_n3520 = 7'h0 ;
assign n3521 =  ( pop ) ? ( bv_1_1_n34 ) : ( bv_1_0_n53 ) ;
assign n3522 =  { ( bv_7_0_n3520 ) , ( n3521 ) }  ;
assign n3523 =  ( sp ) - ( n3522 )  ;
assign n3524 =  ( n3518 ) ? ( n3519 ) : ( n3523 ) ;
assign n3525 =  ( n3516 ) ? ( n3524 ) : ( n3493 ) ;
assign n3526 =  ( n3515 ) ? ( sfr_rd_data ) : ( n3525 ) ;
assign n3527 =  ( n3498 ) ? ( n3500 ) : ( n3526 ) ;
assign n3528 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n3529 =  ( rd_addr ) == ( bv_8_130_n329 )  ;
assign n3530 =  ( n3528 ) & (n3529 )  ;
assign n3531 =  ( wr_sfr ) == ( bv_2_1_n3501 )  ;
assign n3532 =  ( rd_addr ) == ( bv_8_224_n517 )  ;
assign n3533 =  ( n3531 ) & (n3532 )  ;
assign n3534 =  ( wr_sfr ) == ( bv_2_2_n3505 )  ;
assign n3535 =  ( rd_addr ) == ( bv_8_224_n517 )  ;
assign n3536 =  ( n3534 ) & (n3535 )  ;
assign n3537 =  ( n3533 ) | ( n3536 )  ;
assign n3538 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n3539 =  ( rd_addr ) == ( bv_8_131_n331 )  ;
assign n3540 =  ( n3538 ) & (n3539 )  ;
assign n3541 =  ( n3537 ) | ( n3540 )  ;
assign n3542 = wr_addr[7:7] ;
assign n3543 =  ( n3542 ) == ( bv_1_1_n34 )  ;
assign n3544 =  ( rd_addr ) == ( wr_addr )  ;
assign n3545 =  ( n3543 ) & (n3544 )  ;
assign n3546 =  ( wr_bit_r ) == ( 1'b0 )  ;
assign n3547 =  ( n3545 ) & (n3546 )  ;
assign n3548 =  ( n3541 ) | ( n3547 )  ;
assign n3549 = wr_addr[7:7] ;
assign n3550 =  ( n3549 ) == ( bv_1_1_n34 )  ;
assign n3551 = rd_addr[7:3] ;
assign n3552 = wr_addr[7:3] ;
assign n3553 =  ( n3551 ) == ( n3552 )  ;
assign n3554 =  ( n3550 ) & (n3553 )  ;
assign n3555 =  ( n3554 ) & (wr_bit_r )  ;
assign n3556 = rd_addr[2:0] ;
assign bv_3_7_n3557 = 3'h7 ;
assign n3558 =  ( n3556 ) == ( bv_3_7_n3557 )  ;
assign n3559 = ~ ( n3558 )  ;
assign n3560 =  ( n3555 ) & (n3559 )  ;
assign n3561 =  ( n3548 ) | ( n3560 )  ;
assign n3562 =  ( wait_data ) == ( 1'b0 )  ;
assign n3563 =  ( n3561 ) & (n3562 )  ;
assign n3564 =  ( rd_addr ) == ( bv_8_129_n327 )  ;
assign n3565 =  ( ram_wr_sel ) == ( bv_3_3_n3517 )  ;
assign n3566 =  ( sp ) + ( bv_8_1_n71 )  ;
assign n3567 =  ( pop ) ? ( bv_1_1_n34 ) : ( bv_1_0_n53 ) ;
assign n3568 =  { ( bv_7_0_n3520 ) , ( n3567 ) }  ;
assign n3569 =  ( sp ) - ( n3568 )  ;
assign n3570 =  ( n3565 ) ? ( n3566 ) : ( n3569 ) ;
assign n3571 =  ( n3564 ) ? ( n3570 ) : ( n3493 ) ;
assign n3572 =  ( n3563 ) ? ( sfr_rd_data ) : ( n3571 ) ;
assign n3573 =  ( n3530 ) ? ( n3500 ) : ( n3572 ) ;
assign n3574 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n3575 =  ( rd_addr ) == ( bv_8_130_n329 )  ;
assign n3576 =  ( n3574 ) & (n3575 )  ;
assign n3577 =  ( wr_sfr ) == ( bv_2_1_n3501 )  ;
assign n3578 =  ( rd_addr ) == ( bv_8_224_n517 )  ;
assign n3579 =  ( n3577 ) & (n3578 )  ;
assign n3580 =  ( wr_sfr ) == ( bv_2_2_n3505 )  ;
assign n3581 =  ( rd_addr ) == ( bv_8_224_n517 )  ;
assign n3582 =  ( n3580 ) & (n3581 )  ;
assign n3583 =  ( n3579 ) | ( n3582 )  ;
assign n3584 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n3585 =  ( rd_addr ) == ( bv_8_131_n331 )  ;
assign n3586 =  ( n3584 ) & (n3585 )  ;
assign n3587 =  ( n3583 ) | ( n3586 )  ;
assign n3588 =  ( wait_data ) == ( 1'b0 )  ;
assign n3589 =  ( n3587 ) & (n3588 )  ;
assign n3590 =  ( rd_addr ) == ( bv_8_129_n327 )  ;
assign n3591 =  ( ram_wr_sel ) == ( bv_3_3_n3517 )  ;
assign n3592 =  ( sp ) + ( bv_8_1_n71 )  ;
assign n3593 =  ( pop ) ? ( bv_1_1_n34 ) : ( bv_1_0_n53 ) ;
assign n3594 =  { ( bv_7_0_n3520 ) , ( n3593 ) }  ;
assign n3595 =  ( sp ) - ( n3594 )  ;
assign n3596 =  ( n3591 ) ? ( n3592 ) : ( n3595 ) ;
assign n3597 =  ( n3590 ) ? ( n3596 ) : ( n3493 ) ;
assign n3598 =  ( n3589 ) ? ( sfr_rd_data ) : ( n3597 ) ;
assign n3599 =  ( n3576 ) ? ( n3500 ) : ( n3598 ) ;
assign n3600 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n3601 =  ( rd_addr ) == ( bv_8_130_n329 )  ;
assign n3602 =  ( n3600 ) & (n3601 )  ;
assign n3603 =  ( wr_sfr ) == ( bv_2_1_n3501 )  ;
assign n3604 =  ( rd_addr ) == ( bv_8_224_n517 )  ;
assign n3605 =  ( n3603 ) & (n3604 )  ;
assign n3606 =  ( wr_sfr ) == ( bv_2_2_n3505 )  ;
assign n3607 =  ( rd_addr ) == ( bv_8_224_n517 )  ;
assign n3608 =  ( n3606 ) & (n3607 )  ;
assign n3609 =  ( n3605 ) | ( n3608 )  ;
assign n3610 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n3611 =  ( rd_addr ) == ( bv_8_131_n331 )  ;
assign n3612 =  ( n3610 ) & (n3611 )  ;
assign n3613 =  ( n3609 ) | ( n3612 )  ;
assign n3614 = wr_addr[7:7] ;
assign n3615 =  ( n3614 ) == ( bv_1_1_n34 )  ;
assign n3616 =  ( rd_addr ) == ( wr_addr )  ;
assign n3617 =  ( n3615 ) & (n3616 )  ;
assign n3618 =  ( wr_bit_r ) == ( 1'b0 )  ;
assign n3619 =  ( n3617 ) & (n3618 )  ;
assign n3620 =  ( n3613 ) | ( n3619 )  ;
assign n3621 = wr_addr[7:7] ;
assign n3622 =  ( n3621 ) == ( bv_1_1_n34 )  ;
assign n3623 = rd_addr[7:3] ;
assign n3624 = wr_addr[7:3] ;
assign n3625 =  ( n3623 ) == ( n3624 )  ;
assign n3626 =  ( n3622 ) & (n3625 )  ;
assign n3627 =  ( n3626 ) & (wr_bit_r )  ;
assign n3628 = rd_addr[2:0] ;
assign n3629 =  ( n3628 ) == ( bv_3_7_n3557 )  ;
assign n3630 = ~ ( n3629 )  ;
assign n3631 =  ( n3627 ) & (n3630 )  ;
assign n3632 =  ( n3620 ) | ( n3631 )  ;
assign n3633 =  ( wait_data ) == ( 1'b0 )  ;
assign n3634 =  ( n3632 ) & (n3633 )  ;
assign n3635 =  ( rd_addr ) == ( bv_8_129_n327 )  ;
assign n3636 =  ( ram_wr_sel ) == ( bv_3_3_n3517 )  ;
assign n3637 =  ( sp ) + ( bv_8_1_n71 )  ;
assign n3638 =  ( pop ) ? ( bv_1_1_n34 ) : ( bv_1_0_n53 ) ;
assign n3639 =  { ( bv_7_0_n3520 ) , ( n3638 ) }  ;
assign n3640 =  ( sp ) - ( n3639 )  ;
assign n3641 =  ( n3636 ) ? ( n3637 ) : ( n3640 ) ;
assign n3642 =  ( n3635 ) ? ( n3641 ) : ( n3493 ) ;
assign n3643 =  ( n3634 ) ? ( sfr_rd_data ) : ( n3642 ) ;
assign n3644 =  ( n3602 ) ? ( n3500 ) : ( n3643 ) ;
assign n3645 =  ( wr_sfr ) == ( bv_2_1_n3501 )  ;
assign n3646 = rd_addr[7:3] ;
assign bv_5_28_n3647 = 5'h1c ;
assign n3648 =  ( n3646 ) == ( bv_5_28_n3647 )  ;
assign n3649 =  ( n3645 ) & (n3648 )  ;
assign n3650 = rd_addr[2:0] ;
assign n3651 =  ( n3650 ) == ( bv_3_7_n3557 )  ;
assign n3652 = n3500[7:7] ;
assign bv_3_6_n3653 = 3'h6 ;
assign n3654 =  ( n3650 ) == ( bv_3_6_n3653 )  ;
assign n3655 = n3500[6:6] ;
assign bv_3_5_n3656 = 3'h5 ;
assign n3657 =  ( n3650 ) == ( bv_3_5_n3656 )  ;
assign n3658 = n3500[5:5] ;
assign bv_3_4_n3659 = 3'h4 ;
assign n3660 =  ( n3650 ) == ( bv_3_4_n3659 )  ;
assign n3661 = n3500[4:4] ;
assign n3662 =  ( n3650 ) == ( bv_3_3_n3517 )  ;
assign n3663 = n3500[3:3] ;
assign bv_3_2_n3664 = 3'h2 ;
assign n3665 =  ( n3650 ) == ( bv_3_2_n3664 )  ;
assign n3666 = n3500[2:2] ;
assign bv_3_1_n3667 = 3'h1 ;
assign n3668 =  ( n3650 ) == ( bv_3_1_n3667 )  ;
assign n3669 = n3500[1:1] ;
assign n3670 = n3500[0:0] ;
assign n3671 =  ( n3668 ) ? ( n3669 ) : ( n3670 ) ;
assign n3672 =  ( n3665 ) ? ( n3666 ) : ( n3671 ) ;
assign n3673 =  ( n3662 ) ? ( n3663 ) : ( n3672 ) ;
assign n3674 =  ( n3660 ) ? ( n3661 ) : ( n3673 ) ;
assign n3675 =  ( n3657 ) ? ( n3658 ) : ( n3674 ) ;
assign n3676 =  ( n3654 ) ? ( n3655 ) : ( n3675 ) ;
assign n3677 =  ( n3651 ) ? ( n3652 ) : ( n3676 ) ;
assign n3678 =  ( n3646 ) == ( bv_5_28_n3647 )  ;
assign n3679 =  ( n3650 ) == ( bv_3_7_n3557 )  ;
assign n3680 = acc[7:7] ;
assign n3681 =  ( n3650 ) == ( bv_3_6_n3653 )  ;
assign n3682 = acc[6:6] ;
assign n3683 =  ( n3650 ) == ( bv_3_5_n3656 )  ;
assign n3684 = acc[5:5] ;
assign n3685 =  ( n3650 ) == ( bv_3_4_n3659 )  ;
assign n3686 = acc[4:4] ;
assign n3687 =  ( n3650 ) == ( bv_3_3_n3517 )  ;
assign n3688 = acc[3:3] ;
assign n3689 =  ( n3650 ) == ( bv_3_2_n3664 )  ;
assign n3690 = acc[2:2] ;
assign n3691 =  ( n3650 ) == ( bv_3_1_n3667 )  ;
assign n3692 = acc[1:1] ;
assign n3693 = acc[0:0] ;
assign n3694 =  ( n3691 ) ? ( n3692 ) : ( n3693 ) ;
assign n3695 =  ( n3689 ) ? ( n3690 ) : ( n3694 ) ;
assign n3696 =  ( n3687 ) ? ( n3688 ) : ( n3695 ) ;
assign n3697 =  ( n3685 ) ? ( n3686 ) : ( n3696 ) ;
assign n3698 =  ( n3683 ) ? ( n3684 ) : ( n3697 ) ;
assign n3699 =  ( n3681 ) ? ( n3682 ) : ( n3698 ) ;
assign n3700 =  ( n3679 ) ? ( n3680 ) : ( n3699 ) ;
assign bv_5_26_n3701 = 5'h1a ;
assign n3702 =  ( n3646 ) == ( bv_5_26_n3701 )  ;
assign n3703 =  ( n3650 ) == ( bv_3_7_n3557 )  ;
assign n3705 = nondet_psw_next_func_n3704 ;
assign n3706 = n3705[7:7] ;
assign n3707 =  ( n3650 ) == ( bv_3_6_n3653 )  ;
assign n3708 = n3705[6:6] ;
assign n3709 =  ( n3650 ) == ( bv_3_5_n3656 )  ;
assign n3710 = n3705[5:5] ;
assign n3711 =  ( n3650 ) == ( bv_3_4_n3659 )  ;
assign n3712 = n3705[4:4] ;
assign n3713 =  ( n3650 ) == ( bv_3_3_n3517 )  ;
assign n3714 = n3705[3:3] ;
assign n3715 =  ( n3650 ) == ( bv_3_2_n3664 )  ;
assign n3716 = n3705[2:2] ;
assign n3717 =  ( n3650 ) == ( bv_3_1_n3667 )  ;
assign n3718 = n3705[1:1] ;
assign n3719 = n3705[0:0] ;
assign n3720 =  ( n3717 ) ? ( n3718 ) : ( n3719 ) ;
assign n3721 =  ( n3715 ) ? ( n3716 ) : ( n3720 ) ;
assign n3722 =  ( n3713 ) ? ( n3714 ) : ( n3721 ) ;
assign n3723 =  ( n3711 ) ? ( n3712 ) : ( n3722 ) ;
assign n3724 =  ( n3709 ) ? ( n3710 ) : ( n3723 ) ;
assign n3725 =  ( n3707 ) ? ( n3708 ) : ( n3724 ) ;
assign n3726 =  ( n3703 ) ? ( n3706 ) : ( n3725 ) ;
assign bv_5_16_n3727 = 5'h10 ;
assign n3728 =  ( n3646 ) == ( bv_5_16_n3727 )  ;
assign n3729 =  ( n3650 ) == ( bv_3_7_n3557 )  ;
assign n3730 = p0[7:7] ;
assign n3731 =  ( n3650 ) == ( bv_3_6_n3653 )  ;
assign n3732 = p0[6:6] ;
assign n3733 =  ( n3650 ) == ( bv_3_5_n3656 )  ;
assign n3734 = p0[5:5] ;
assign n3735 =  ( n3650 ) == ( bv_3_4_n3659 )  ;
assign n3736 = p0[4:4] ;
assign n3737 =  ( n3650 ) == ( bv_3_3_n3517 )  ;
assign n3738 = p0[3:3] ;
assign n3739 =  ( n3650 ) == ( bv_3_2_n3664 )  ;
assign n3740 = p0[2:2] ;
assign n3741 =  ( n3650 ) == ( bv_3_1_n3667 )  ;
assign n3742 = p0[1:1] ;
assign n3743 = p0[0:0] ;
assign n3744 =  ( n3741 ) ? ( n3742 ) : ( n3743 ) ;
assign n3745 =  ( n3739 ) ? ( n3740 ) : ( n3744 ) ;
assign n3746 =  ( n3737 ) ? ( n3738 ) : ( n3745 ) ;
assign n3747 =  ( n3735 ) ? ( n3736 ) : ( n3746 ) ;
assign n3748 =  ( n3733 ) ? ( n3734 ) : ( n3747 ) ;
assign n3749 =  ( n3731 ) ? ( n3732 ) : ( n3748 ) ;
assign n3750 =  ( n3729 ) ? ( n3730 ) : ( n3749 ) ;
assign bv_5_18_n3751 = 5'h12 ;
assign n3752 =  ( n3646 ) == ( bv_5_18_n3751 )  ;
assign n3753 =  ( n3650 ) == ( bv_3_7_n3557 )  ;
assign n3754 = p1[7:7] ;
assign n3755 =  ( n3650 ) == ( bv_3_6_n3653 )  ;
assign n3756 = p1[6:6] ;
assign n3757 =  ( n3650 ) == ( bv_3_5_n3656 )  ;
assign n3758 = p1[5:5] ;
assign n3759 =  ( n3650 ) == ( bv_3_4_n3659 )  ;
assign n3760 = p1[4:4] ;
assign n3761 =  ( n3650 ) == ( bv_3_3_n3517 )  ;
assign n3762 = p1[3:3] ;
assign n3763 =  ( n3650 ) == ( bv_3_2_n3664 )  ;
assign n3764 = p1[2:2] ;
assign n3765 =  ( n3650 ) == ( bv_3_1_n3667 )  ;
assign n3766 = p1[1:1] ;
assign n3767 = p1[0:0] ;
assign n3768 =  ( n3765 ) ? ( n3766 ) : ( n3767 ) ;
assign n3769 =  ( n3763 ) ? ( n3764 ) : ( n3768 ) ;
assign n3770 =  ( n3761 ) ? ( n3762 ) : ( n3769 ) ;
assign n3771 =  ( n3759 ) ? ( n3760 ) : ( n3770 ) ;
assign n3772 =  ( n3757 ) ? ( n3758 ) : ( n3771 ) ;
assign n3773 =  ( n3755 ) ? ( n3756 ) : ( n3772 ) ;
assign n3774 =  ( n3753 ) ? ( n3754 ) : ( n3773 ) ;
assign bv_5_20_n3775 = 5'h14 ;
assign n3776 =  ( n3646 ) == ( bv_5_20_n3775 )  ;
assign n3777 =  ( n3650 ) == ( bv_3_7_n3557 )  ;
assign n3778 = p2[7:7] ;
assign n3779 =  ( n3650 ) == ( bv_3_6_n3653 )  ;
assign n3780 = p2[6:6] ;
assign n3781 =  ( n3650 ) == ( bv_3_5_n3656 )  ;
assign n3782 = p2[5:5] ;
assign n3783 =  ( n3650 ) == ( bv_3_4_n3659 )  ;
assign n3784 = p2[4:4] ;
assign n3785 =  ( n3650 ) == ( bv_3_3_n3517 )  ;
assign n3786 = p2[3:3] ;
assign n3787 =  ( n3650 ) == ( bv_3_2_n3664 )  ;
assign n3788 = p2[2:2] ;
assign n3789 =  ( n3650 ) == ( bv_3_1_n3667 )  ;
assign n3790 = p2[1:1] ;
assign n3791 = p2[0:0] ;
assign n3792 =  ( n3789 ) ? ( n3790 ) : ( n3791 ) ;
assign n3793 =  ( n3787 ) ? ( n3788 ) : ( n3792 ) ;
assign n3794 =  ( n3785 ) ? ( n3786 ) : ( n3793 ) ;
assign n3795 =  ( n3783 ) ? ( n3784 ) : ( n3794 ) ;
assign n3796 =  ( n3781 ) ? ( n3782 ) : ( n3795 ) ;
assign n3797 =  ( n3779 ) ? ( n3780 ) : ( n3796 ) ;
assign n3798 =  ( n3777 ) ? ( n3778 ) : ( n3797 ) ;
assign bv_5_22_n3799 = 5'h16 ;
assign n3800 =  ( n3646 ) == ( bv_5_22_n3799 )  ;
assign n3801 =  ( n3650 ) == ( bv_3_7_n3557 )  ;
assign n3802 = p3[7:7] ;
assign n3803 =  ( n3650 ) == ( bv_3_6_n3653 )  ;
assign n3804 = p3[6:6] ;
assign n3805 =  ( n3650 ) == ( bv_3_5_n3656 )  ;
assign n3806 = p3[5:5] ;
assign n3807 =  ( n3650 ) == ( bv_3_4_n3659 )  ;
assign n3808 = p3[4:4] ;
assign n3809 =  ( n3650 ) == ( bv_3_3_n3517 )  ;
assign n3810 = p3[3:3] ;
assign n3811 =  ( n3650 ) == ( bv_3_2_n3664 )  ;
assign n3812 = p3[2:2] ;
assign n3813 =  ( n3650 ) == ( bv_3_1_n3667 )  ;
assign n3814 = p3[1:1] ;
assign n3815 = p3[0:0] ;
assign n3816 =  ( n3813 ) ? ( n3814 ) : ( n3815 ) ;
assign n3817 =  ( n3811 ) ? ( n3812 ) : ( n3816 ) ;
assign n3818 =  ( n3809 ) ? ( n3810 ) : ( n3817 ) ;
assign n3819 =  ( n3807 ) ? ( n3808 ) : ( n3818 ) ;
assign n3820 =  ( n3805 ) ? ( n3806 ) : ( n3819 ) ;
assign n3821 =  ( n3803 ) ? ( n3804 ) : ( n3820 ) ;
assign n3822 =  ( n3801 ) ? ( n3802 ) : ( n3821 ) ;
assign bv_5_30_n3823 = 5'h1e ;
assign n3824 =  ( n3646 ) == ( bv_5_30_n3823 )  ;
assign n3825 =  ( n3650 ) == ( bv_3_7_n3557 )  ;
assign n3826 = b_reg[7:7] ;
assign n3827 =  ( n3650 ) == ( bv_3_6_n3653 )  ;
assign n3828 = b_reg[6:6] ;
assign n3829 =  ( n3650 ) == ( bv_3_5_n3656 )  ;
assign n3830 = b_reg[5:5] ;
assign n3831 =  ( n3650 ) == ( bv_3_4_n3659 )  ;
assign n3832 = b_reg[4:4] ;
assign n3833 =  ( n3650 ) == ( bv_3_3_n3517 )  ;
assign n3834 = b_reg[3:3] ;
assign n3835 =  ( n3650 ) == ( bv_3_2_n3664 )  ;
assign n3836 = b_reg[2:2] ;
assign n3837 =  ( n3650 ) == ( bv_3_1_n3667 )  ;
assign n3838 = b_reg[1:1] ;
assign n3839 = b_reg[0:0] ;
assign n3840 =  ( n3837 ) ? ( n3838 ) : ( n3839 ) ;
assign n3841 =  ( n3835 ) ? ( n3836 ) : ( n3840 ) ;
assign n3842 =  ( n3833 ) ? ( n3834 ) : ( n3841 ) ;
assign n3843 =  ( n3831 ) ? ( n3832 ) : ( n3842 ) ;
assign n3844 =  ( n3829 ) ? ( n3830 ) : ( n3843 ) ;
assign n3845 =  ( n3827 ) ? ( n3828 ) : ( n3844 ) ;
assign n3846 =  ( n3825 ) ? ( n3826 ) : ( n3845 ) ;
assign bv_5_23_n3847 = 5'h17 ;
assign n3848 =  ( n3646 ) == ( bv_5_23_n3847 )  ;
assign n3849 =  ( n3650 ) == ( bv_3_7_n3557 )  ;
assign n3850 = ip[7:7] ;
assign n3851 =  ( n3650 ) == ( bv_3_6_n3653 )  ;
assign n3852 = ip[6:6] ;
assign n3853 =  ( n3650 ) == ( bv_3_5_n3656 )  ;
assign n3854 = ip[5:5] ;
assign n3855 =  ( n3650 ) == ( bv_3_4_n3659 )  ;
assign n3856 = ip[4:4] ;
assign n3857 =  ( n3650 ) == ( bv_3_3_n3517 )  ;
assign n3858 = ip[3:3] ;
assign n3859 =  ( n3650 ) == ( bv_3_2_n3664 )  ;
assign n3860 = ip[2:2] ;
assign n3861 =  ( n3650 ) == ( bv_3_1_n3667 )  ;
assign n3862 = ip[1:1] ;
assign n3863 = ip[0:0] ;
assign n3864 =  ( n3861 ) ? ( n3862 ) : ( n3863 ) ;
assign n3865 =  ( n3859 ) ? ( n3860 ) : ( n3864 ) ;
assign n3866 =  ( n3857 ) ? ( n3858 ) : ( n3865 ) ;
assign n3867 =  ( n3855 ) ? ( n3856 ) : ( n3866 ) ;
assign n3868 =  ( n3853 ) ? ( n3854 ) : ( n3867 ) ;
assign n3869 =  ( n3851 ) ? ( n3852 ) : ( n3868 ) ;
assign n3870 =  ( n3849 ) ? ( n3850 ) : ( n3869 ) ;
assign bv_5_21_n3871 = 5'h15 ;
assign n3872 =  ( n3646 ) == ( bv_5_21_n3871 )  ;
assign n3873 =  ( n3650 ) == ( bv_3_7_n3557 )  ;
assign n3874 = ie[7:7] ;
assign n3875 =  ( n3650 ) == ( bv_3_6_n3653 )  ;
assign n3876 = ie[6:6] ;
assign n3877 =  ( n3650 ) == ( bv_3_5_n3656 )  ;
assign n3878 = ie[5:5] ;
assign n3879 =  ( n3650 ) == ( bv_3_4_n3659 )  ;
assign n3880 = ie[4:4] ;
assign n3881 =  ( n3650 ) == ( bv_3_3_n3517 )  ;
assign n3882 = ie[3:3] ;
assign n3883 =  ( n3650 ) == ( bv_3_2_n3664 )  ;
assign n3884 = ie[2:2] ;
assign n3885 =  ( n3650 ) == ( bv_3_1_n3667 )  ;
assign n3886 = ie[1:1] ;
assign n3887 = ie[0:0] ;
assign n3888 =  ( n3885 ) ? ( n3886 ) : ( n3887 ) ;
assign n3889 =  ( n3883 ) ? ( n3884 ) : ( n3888 ) ;
assign n3890 =  ( n3881 ) ? ( n3882 ) : ( n3889 ) ;
assign n3891 =  ( n3879 ) ? ( n3880 ) : ( n3890 ) ;
assign n3892 =  ( n3877 ) ? ( n3878 ) : ( n3891 ) ;
assign n3893 =  ( n3875 ) ? ( n3876 ) : ( n3892 ) ;
assign n3894 =  ( n3873 ) ? ( n3874 ) : ( n3893 ) ;
assign n3895 =  ( n3872 ) ? ( n3894 ) : ( bv_1_0_n53 ) ;
assign n3896 =  ( n3848 ) ? ( n3870 ) : ( n3895 ) ;
assign n3897 =  ( n3824 ) ? ( n3846 ) : ( n3896 ) ;
assign n3898 =  ( n3800 ) ? ( n3822 ) : ( n3897 ) ;
assign n3899 =  ( n3776 ) ? ( n3798 ) : ( n3898 ) ;
assign n3900 =  ( n3752 ) ? ( n3774 ) : ( n3899 ) ;
assign n3901 =  ( n3728 ) ? ( n3750 ) : ( n3900 ) ;
assign n3902 =  ( n3702 ) ? ( n3726 ) : ( n3901 ) ;
assign n3903 =  ( n3678 ) ? ( n3700 ) : ( n3902 ) ;
assign n3904 =  ( n3649 ) ? ( n3677 ) : ( n3903 ) ;
assign n3905 = rd_addr[7:3] ;
assign n3906 = wr_addr[7:3] ;
assign n3907 =  ( n3905 ) == ( n3906 )  ;
assign n3908 =  ( wr_bit_r ) == ( 1'b0 )  ;
assign n3909 =  ( n3907 ) & (n3908 )  ;
assign n3910 = wr_addr[2:0] ;
assign n3911 =  ( n3910 ) == ( bv_3_0_n46 )  ;
assign n3912 =  ( n3909 ) & (n3911 )  ;
assign n3913 = rd_addr[7:3] ;
assign n3914 =  ( n3913 ) == ( bv_5_28_n3647 )  ;
assign n3915 = rd_addr[7:3] ;
assign n3916 =  ( n3915 ) == ( bv_5_26_n3701 )  ;
assign n3917 =  ( n3914 ) | ( n3916 )  ;
assign n3918 = rd_addr[7:3] ;
assign n3919 =  ( n3918 ) == ( bv_5_30_n3823 )  ;
assign n3920 =  ( n3917 ) | ( n3919 )  ;
assign n3921 = rd_addr[7:3] ;
assign n3922 =  ( n3921 ) == ( bv_5_16_n3727 )  ;
assign n3923 =  ( n3920 ) | ( n3922 )  ;
assign n3924 = rd_addr[7:3] ;
assign n3925 =  ( n3924 ) == ( bv_5_18_n3751 )  ;
assign n3926 =  ( n3923 ) | ( n3925 )  ;
assign n3927 = rd_addr[7:3] ;
assign n3928 =  ( n3927 ) == ( bv_5_20_n3775 )  ;
assign n3929 =  ( n3926 ) | ( n3928 )  ;
assign n3930 = rd_addr[7:3] ;
assign n3931 =  ( n3930 ) == ( bv_5_22_n3799 )  ;
assign n3932 =  ( n3929 ) | ( n3931 )  ;
assign n3933 =  ( n3912 ) & (n3932 )  ;
assign n3934 = rd_addr[2:0] ;
assign n3935 =  ( n3934 ) == ( bv_3_7_n3557 )  ;
assign n3937 = nondet_des1_func_n3936 ;
assign n3938 = n3937[7:7] ;
assign n3939 =  ( n3934 ) == ( bv_3_6_n3653 )  ;
assign n3940 = n3937[6:6] ;
assign n3941 =  ( n3934 ) == ( bv_3_5_n3656 )  ;
assign n3942 = n3937[5:5] ;
assign n3943 =  ( n3934 ) == ( bv_3_4_n3659 )  ;
assign n3944 = n3937[4:4] ;
assign n3945 =  ( n3934 ) == ( bv_3_3_n3517 )  ;
assign n3946 = n3937[3:3] ;
assign n3947 =  ( n3934 ) == ( bv_3_2_n3664 )  ;
assign n3948 = n3937[2:2] ;
assign n3949 =  ( n3934 ) == ( bv_3_1_n3667 )  ;
assign n3950 = n3937[1:1] ;
assign n3951 = n3937[0:0] ;
assign n3952 =  ( n3949 ) ? ( n3950 ) : ( n3951 ) ;
assign n3953 =  ( n3947 ) ? ( n3948 ) : ( n3952 ) ;
assign n3954 =  ( n3945 ) ? ( n3946 ) : ( n3953 ) ;
assign n3955 =  ( n3943 ) ? ( n3944 ) : ( n3954 ) ;
assign n3956 =  ( n3941 ) ? ( n3942 ) : ( n3955 ) ;
assign n3957 =  ( n3939 ) ? ( n3940 ) : ( n3956 ) ;
assign n3958 =  ( n3935 ) ? ( n3938 ) : ( n3957 ) ;
assign n3959 =  ( wr_sfr ) == ( bv_2_1_n3501 )  ;
assign n3960 = rd_addr[7:3] ;
assign n3961 =  ( n3960 ) == ( bv_5_28_n3647 )  ;
assign n3962 =  ( n3959 ) & (n3961 )  ;
assign n3963 =  ( n3934 ) == ( bv_3_7_n3557 )  ;
assign n3964 = n3500[7:7] ;
assign n3965 =  ( n3934 ) == ( bv_3_6_n3653 )  ;
assign n3966 = n3500[6:6] ;
assign n3967 =  ( n3934 ) == ( bv_3_5_n3656 )  ;
assign n3968 = n3500[5:5] ;
assign n3969 =  ( n3934 ) == ( bv_3_4_n3659 )  ;
assign n3970 = n3500[4:4] ;
assign n3971 =  ( n3934 ) == ( bv_3_3_n3517 )  ;
assign n3972 = n3500[3:3] ;
assign n3973 =  ( n3934 ) == ( bv_3_2_n3664 )  ;
assign n3974 = n3500[2:2] ;
assign n3975 =  ( n3934 ) == ( bv_3_1_n3667 )  ;
assign n3976 = n3500[1:1] ;
assign n3977 = n3500[0:0] ;
assign n3978 =  ( n3975 ) ? ( n3976 ) : ( n3977 ) ;
assign n3979 =  ( n3973 ) ? ( n3974 ) : ( n3978 ) ;
assign n3980 =  ( n3971 ) ? ( n3972 ) : ( n3979 ) ;
assign n3981 =  ( n3969 ) ? ( n3970 ) : ( n3980 ) ;
assign n3982 =  ( n3967 ) ? ( n3968 ) : ( n3981 ) ;
assign n3983 =  ( n3965 ) ? ( n3966 ) : ( n3982 ) ;
assign n3984 =  ( n3963 ) ? ( n3964 ) : ( n3983 ) ;
assign n3985 =  ( rd_addr ) == ( wr_addr )  ;
assign n3986 =  ( n3985 ) & (wr_bit_r )  ;
assign n3987 =  ( n3986 ) & (n3932 )  ;
assign n3989 = nondet_desCy_func_n3988 ;
assign n3990 =  ( n3960 ) == ( bv_5_28_n3647 )  ;
assign n3991 =  ( n3934 ) == ( bv_3_7_n3557 )  ;
assign n3992 = acc[7:7] ;
assign n3993 =  ( n3934 ) == ( bv_3_6_n3653 )  ;
assign n3994 = acc[6:6] ;
assign n3995 =  ( n3934 ) == ( bv_3_5_n3656 )  ;
assign n3996 = acc[5:5] ;
assign n3997 =  ( n3934 ) == ( bv_3_4_n3659 )  ;
assign n3998 = acc[4:4] ;
assign n3999 =  ( n3934 ) == ( bv_3_3_n3517 )  ;
assign n4000 = acc[3:3] ;
assign n4001 =  ( n3934 ) == ( bv_3_2_n3664 )  ;
assign n4002 = acc[2:2] ;
assign n4003 =  ( n3934 ) == ( bv_3_1_n3667 )  ;
assign n4004 = acc[1:1] ;
assign n4005 = acc[0:0] ;
assign n4006 =  ( n4003 ) ? ( n4004 ) : ( n4005 ) ;
assign n4007 =  ( n4001 ) ? ( n4002 ) : ( n4006 ) ;
assign n4008 =  ( n3999 ) ? ( n4000 ) : ( n4007 ) ;
assign n4009 =  ( n3997 ) ? ( n3998 ) : ( n4008 ) ;
assign n4010 =  ( n3995 ) ? ( n3996 ) : ( n4009 ) ;
assign n4011 =  ( n3993 ) ? ( n3994 ) : ( n4010 ) ;
assign n4012 =  ( n3991 ) ? ( n3992 ) : ( n4011 ) ;
assign n4013 =  ( n3960 ) == ( bv_5_26_n3701 )  ;
assign n4014 =  ( n3934 ) == ( bv_3_7_n3557 )  ;
assign n4015 = n3705[7:7] ;
assign n4016 =  ( n3934 ) == ( bv_3_6_n3653 )  ;
assign n4017 = n3705[6:6] ;
assign n4018 =  ( n3934 ) == ( bv_3_5_n3656 )  ;
assign n4019 = n3705[5:5] ;
assign n4020 =  ( n3934 ) == ( bv_3_4_n3659 )  ;
assign n4021 = n3705[4:4] ;
assign n4022 =  ( n3934 ) == ( bv_3_3_n3517 )  ;
assign n4023 = n3705[3:3] ;
assign n4024 =  ( n3934 ) == ( bv_3_2_n3664 )  ;
assign n4025 = n3705[2:2] ;
assign n4026 =  ( n3934 ) == ( bv_3_1_n3667 )  ;
assign n4027 = n3705[1:1] ;
assign n4028 = n3705[0:0] ;
assign n4029 =  ( n4026 ) ? ( n4027 ) : ( n4028 ) ;
assign n4030 =  ( n4024 ) ? ( n4025 ) : ( n4029 ) ;
assign n4031 =  ( n4022 ) ? ( n4023 ) : ( n4030 ) ;
assign n4032 =  ( n4020 ) ? ( n4021 ) : ( n4031 ) ;
assign n4033 =  ( n4018 ) ? ( n4019 ) : ( n4032 ) ;
assign n4034 =  ( n4016 ) ? ( n4017 ) : ( n4033 ) ;
assign n4035 =  ( n4014 ) ? ( n4015 ) : ( n4034 ) ;
assign n4036 =  ( n3960 ) == ( bv_5_16_n3727 )  ;
assign n4037 =  ( n3934 ) == ( bv_3_7_n3557 )  ;
assign n4038 = p0[7:7] ;
assign n4039 =  ( n3934 ) == ( bv_3_6_n3653 )  ;
assign n4040 = p0[6:6] ;
assign n4041 =  ( n3934 ) == ( bv_3_5_n3656 )  ;
assign n4042 = p0[5:5] ;
assign n4043 =  ( n3934 ) == ( bv_3_4_n3659 )  ;
assign n4044 = p0[4:4] ;
assign n4045 =  ( n3934 ) == ( bv_3_3_n3517 )  ;
assign n4046 = p0[3:3] ;
assign n4047 =  ( n3934 ) == ( bv_3_2_n3664 )  ;
assign n4048 = p0[2:2] ;
assign n4049 =  ( n3934 ) == ( bv_3_1_n3667 )  ;
assign n4050 = p0[1:1] ;
assign n4051 = p0[0:0] ;
assign n4052 =  ( n4049 ) ? ( n4050 ) : ( n4051 ) ;
assign n4053 =  ( n4047 ) ? ( n4048 ) : ( n4052 ) ;
assign n4054 =  ( n4045 ) ? ( n4046 ) : ( n4053 ) ;
assign n4055 =  ( n4043 ) ? ( n4044 ) : ( n4054 ) ;
assign n4056 =  ( n4041 ) ? ( n4042 ) : ( n4055 ) ;
assign n4057 =  ( n4039 ) ? ( n4040 ) : ( n4056 ) ;
assign n4058 =  ( n4037 ) ? ( n4038 ) : ( n4057 ) ;
assign n4059 =  ( n3960 ) == ( bv_5_18_n3751 )  ;
assign n4060 =  ( n3934 ) == ( bv_3_7_n3557 )  ;
assign n4061 = p1[7:7] ;
assign n4062 =  ( n3934 ) == ( bv_3_6_n3653 )  ;
assign n4063 = p1[6:6] ;
assign n4064 =  ( n3934 ) == ( bv_3_5_n3656 )  ;
assign n4065 = p1[5:5] ;
assign n4066 =  ( n3934 ) == ( bv_3_4_n3659 )  ;
assign n4067 = p1[4:4] ;
assign n4068 =  ( n3934 ) == ( bv_3_3_n3517 )  ;
assign n4069 = p1[3:3] ;
assign n4070 =  ( n3934 ) == ( bv_3_2_n3664 )  ;
assign n4071 = p1[2:2] ;
assign n4072 =  ( n3934 ) == ( bv_3_1_n3667 )  ;
assign n4073 = p1[1:1] ;
assign n4074 = p1[0:0] ;
assign n4075 =  ( n4072 ) ? ( n4073 ) : ( n4074 ) ;
assign n4076 =  ( n4070 ) ? ( n4071 ) : ( n4075 ) ;
assign n4077 =  ( n4068 ) ? ( n4069 ) : ( n4076 ) ;
assign n4078 =  ( n4066 ) ? ( n4067 ) : ( n4077 ) ;
assign n4079 =  ( n4064 ) ? ( n4065 ) : ( n4078 ) ;
assign n4080 =  ( n4062 ) ? ( n4063 ) : ( n4079 ) ;
assign n4081 =  ( n4060 ) ? ( n4061 ) : ( n4080 ) ;
assign n4082 =  ( n3960 ) == ( bv_5_20_n3775 )  ;
assign n4083 =  ( n3934 ) == ( bv_3_7_n3557 )  ;
assign n4084 = p2[7:7] ;
assign n4085 =  ( n3934 ) == ( bv_3_6_n3653 )  ;
assign n4086 = p2[6:6] ;
assign n4087 =  ( n3934 ) == ( bv_3_5_n3656 )  ;
assign n4088 = p2[5:5] ;
assign n4089 =  ( n3934 ) == ( bv_3_4_n3659 )  ;
assign n4090 = p2[4:4] ;
assign n4091 =  ( n3934 ) == ( bv_3_3_n3517 )  ;
assign n4092 = p2[3:3] ;
assign n4093 =  ( n3934 ) == ( bv_3_2_n3664 )  ;
assign n4094 = p2[2:2] ;
assign n4095 =  ( n3934 ) == ( bv_3_1_n3667 )  ;
assign n4096 = p2[1:1] ;
assign n4097 = p2[0:0] ;
assign n4098 =  ( n4095 ) ? ( n4096 ) : ( n4097 ) ;
assign n4099 =  ( n4093 ) ? ( n4094 ) : ( n4098 ) ;
assign n4100 =  ( n4091 ) ? ( n4092 ) : ( n4099 ) ;
assign n4101 =  ( n4089 ) ? ( n4090 ) : ( n4100 ) ;
assign n4102 =  ( n4087 ) ? ( n4088 ) : ( n4101 ) ;
assign n4103 =  ( n4085 ) ? ( n4086 ) : ( n4102 ) ;
assign n4104 =  ( n4083 ) ? ( n4084 ) : ( n4103 ) ;
assign n4105 =  ( n3960 ) == ( bv_5_22_n3799 )  ;
assign n4106 =  ( n3934 ) == ( bv_3_7_n3557 )  ;
assign n4107 = p3[7:7] ;
assign n4108 =  ( n3934 ) == ( bv_3_6_n3653 )  ;
assign n4109 = p3[6:6] ;
assign n4110 =  ( n3934 ) == ( bv_3_5_n3656 )  ;
assign n4111 = p3[5:5] ;
assign n4112 =  ( n3934 ) == ( bv_3_4_n3659 )  ;
assign n4113 = p3[4:4] ;
assign n4114 =  ( n3934 ) == ( bv_3_3_n3517 )  ;
assign n4115 = p3[3:3] ;
assign n4116 =  ( n3934 ) == ( bv_3_2_n3664 )  ;
assign n4117 = p3[2:2] ;
assign n4118 =  ( n3934 ) == ( bv_3_1_n3667 )  ;
assign n4119 = p3[1:1] ;
assign n4120 = p3[0:0] ;
assign n4121 =  ( n4118 ) ? ( n4119 ) : ( n4120 ) ;
assign n4122 =  ( n4116 ) ? ( n4117 ) : ( n4121 ) ;
assign n4123 =  ( n4114 ) ? ( n4115 ) : ( n4122 ) ;
assign n4124 =  ( n4112 ) ? ( n4113 ) : ( n4123 ) ;
assign n4125 =  ( n4110 ) ? ( n4111 ) : ( n4124 ) ;
assign n4126 =  ( n4108 ) ? ( n4109 ) : ( n4125 ) ;
assign n4127 =  ( n4106 ) ? ( n4107 ) : ( n4126 ) ;
assign n4128 =  ( n3960 ) == ( bv_5_30_n3823 )  ;
assign n4129 =  ( n3934 ) == ( bv_3_7_n3557 )  ;
assign n4130 = b_reg[7:7] ;
assign n4131 =  ( n3934 ) == ( bv_3_6_n3653 )  ;
assign n4132 = b_reg[6:6] ;
assign n4133 =  ( n3934 ) == ( bv_3_5_n3656 )  ;
assign n4134 = b_reg[5:5] ;
assign n4135 =  ( n3934 ) == ( bv_3_4_n3659 )  ;
assign n4136 = b_reg[4:4] ;
assign n4137 =  ( n3934 ) == ( bv_3_3_n3517 )  ;
assign n4138 = b_reg[3:3] ;
assign n4139 =  ( n3934 ) == ( bv_3_2_n3664 )  ;
assign n4140 = b_reg[2:2] ;
assign n4141 =  ( n3934 ) == ( bv_3_1_n3667 )  ;
assign n4142 = b_reg[1:1] ;
assign n4143 = b_reg[0:0] ;
assign n4144 =  ( n4141 ) ? ( n4142 ) : ( n4143 ) ;
assign n4145 =  ( n4139 ) ? ( n4140 ) : ( n4144 ) ;
assign n4146 =  ( n4137 ) ? ( n4138 ) : ( n4145 ) ;
assign n4147 =  ( n4135 ) ? ( n4136 ) : ( n4146 ) ;
assign n4148 =  ( n4133 ) ? ( n4134 ) : ( n4147 ) ;
assign n4149 =  ( n4131 ) ? ( n4132 ) : ( n4148 ) ;
assign n4150 =  ( n4129 ) ? ( n4130 ) : ( n4149 ) ;
assign n4151 =  ( n3960 ) == ( bv_5_23_n3847 )  ;
assign n4152 =  ( n3934 ) == ( bv_3_7_n3557 )  ;
assign n4153 = ip[7:7] ;
assign n4154 =  ( n3934 ) == ( bv_3_6_n3653 )  ;
assign n4155 = ip[6:6] ;
assign n4156 =  ( n3934 ) == ( bv_3_5_n3656 )  ;
assign n4157 = ip[5:5] ;
assign n4158 =  ( n3934 ) == ( bv_3_4_n3659 )  ;
assign n4159 = ip[4:4] ;
assign n4160 =  ( n3934 ) == ( bv_3_3_n3517 )  ;
assign n4161 = ip[3:3] ;
assign n4162 =  ( n3934 ) == ( bv_3_2_n3664 )  ;
assign n4163 = ip[2:2] ;
assign n4164 =  ( n3934 ) == ( bv_3_1_n3667 )  ;
assign n4165 = ip[1:1] ;
assign n4166 = ip[0:0] ;
assign n4167 =  ( n4164 ) ? ( n4165 ) : ( n4166 ) ;
assign n4168 =  ( n4162 ) ? ( n4163 ) : ( n4167 ) ;
assign n4169 =  ( n4160 ) ? ( n4161 ) : ( n4168 ) ;
assign n4170 =  ( n4158 ) ? ( n4159 ) : ( n4169 ) ;
assign n4171 =  ( n4156 ) ? ( n4157 ) : ( n4170 ) ;
assign n4172 =  ( n4154 ) ? ( n4155 ) : ( n4171 ) ;
assign n4173 =  ( n4152 ) ? ( n4153 ) : ( n4172 ) ;
assign n4174 =  ( n3960 ) == ( bv_5_21_n3871 )  ;
assign n4175 =  ( n3934 ) == ( bv_3_7_n3557 )  ;
assign n4176 = ie[7:7] ;
assign n4177 =  ( n3934 ) == ( bv_3_6_n3653 )  ;
assign n4178 = ie[6:6] ;
assign n4179 =  ( n3934 ) == ( bv_3_5_n3656 )  ;
assign n4180 = ie[5:5] ;
assign n4181 =  ( n3934 ) == ( bv_3_4_n3659 )  ;
assign n4182 = ie[4:4] ;
assign n4183 =  ( n3934 ) == ( bv_3_3_n3517 )  ;
assign n4184 = ie[3:3] ;
assign n4185 =  ( n3934 ) == ( bv_3_2_n3664 )  ;
assign n4186 = ie[2:2] ;
assign n4187 =  ( n3934 ) == ( bv_3_1_n3667 )  ;
assign n4188 = ie[1:1] ;
assign n4189 = ie[0:0] ;
assign n4190 =  ( n4187 ) ? ( n4188 ) : ( n4189 ) ;
assign n4191 =  ( n4185 ) ? ( n4186 ) : ( n4190 ) ;
assign n4192 =  ( n4183 ) ? ( n4184 ) : ( n4191 ) ;
assign n4193 =  ( n4181 ) ? ( n4182 ) : ( n4192 ) ;
assign n4194 =  ( n4179 ) ? ( n4180 ) : ( n4193 ) ;
assign n4195 =  ( n4177 ) ? ( n4178 ) : ( n4194 ) ;
assign n4196 =  ( n4175 ) ? ( n4176 ) : ( n4195 ) ;
assign n4197 =  ( n4174 ) ? ( n4196 ) : ( bv_1_0_n53 ) ;
assign n4198 =  ( n4151 ) ? ( n4173 ) : ( n4197 ) ;
assign n4199 =  ( n4128 ) ? ( n4150 ) : ( n4198 ) ;
assign n4200 =  ( n4105 ) ? ( n4127 ) : ( n4199 ) ;
assign n4201 =  ( n4082 ) ? ( n4104 ) : ( n4200 ) ;
assign n4202 =  ( n4059 ) ? ( n4081 ) : ( n4201 ) ;
assign n4203 =  ( n4036 ) ? ( n4058 ) : ( n4202 ) ;
assign n4204 =  ( n4013 ) ? ( n4035 ) : ( n4203 ) ;
assign n4205 =  ( n3990 ) ? ( n4012 ) : ( n4204 ) ;
assign n4206 =  ( n3987 ) ? ( n3989 ) : ( n4205 ) ;
assign n4207 =  ( n3962 ) ? ( n3984 ) : ( n4206 ) ;
assign n4208 =  ( n3933 ) ? ( n3958 ) : ( n4207 ) ;
assign n4209 =  ( wr_sfr ) == ( bv_2_1_n3501 )  ;
assign n4210 = rd_addr[7:3] ;
assign n4211 =  ( n4210 ) == ( bv_5_28_n3647 )  ;
assign n4212 =  ( n4209 ) & (n4211 )  ;
assign n4213 = rd_addr[2:0] ;
assign n4214 =  ( n4213 ) == ( bv_3_7_n3557 )  ;
assign n4215 = n3500[7:7] ;
assign n4216 =  ( n4213 ) == ( bv_3_6_n3653 )  ;
assign n4217 = n3500[6:6] ;
assign n4218 =  ( n4213 ) == ( bv_3_5_n3656 )  ;
assign n4219 = n3500[5:5] ;
assign n4220 =  ( n4213 ) == ( bv_3_4_n3659 )  ;
assign n4221 = n3500[4:4] ;
assign n4222 =  ( n4213 ) == ( bv_3_3_n3517 )  ;
assign n4223 = n3500[3:3] ;
assign n4224 =  ( n4213 ) == ( bv_3_2_n3664 )  ;
assign n4225 = n3500[2:2] ;
assign n4226 =  ( n4213 ) == ( bv_3_1_n3667 )  ;
assign n4227 = n3500[1:1] ;
assign n4228 = n3500[0:0] ;
assign n4229 =  ( n4226 ) ? ( n4227 ) : ( n4228 ) ;
assign n4230 =  ( n4224 ) ? ( n4225 ) : ( n4229 ) ;
assign n4231 =  ( n4222 ) ? ( n4223 ) : ( n4230 ) ;
assign n4232 =  ( n4220 ) ? ( n4221 ) : ( n4231 ) ;
assign n4233 =  ( n4218 ) ? ( n4219 ) : ( n4232 ) ;
assign n4234 =  ( n4216 ) ? ( n4217 ) : ( n4233 ) ;
assign n4235 =  ( n4214 ) ? ( n4215 ) : ( n4234 ) ;
assign n4236 =  ( n4210 ) == ( bv_5_28_n3647 )  ;
assign n4237 =  ( n4213 ) == ( bv_3_7_n3557 )  ;
assign n4238 = acc[7:7] ;
assign n4239 =  ( n4213 ) == ( bv_3_6_n3653 )  ;
assign n4240 = acc[6:6] ;
assign n4241 =  ( n4213 ) == ( bv_3_5_n3656 )  ;
assign n4242 = acc[5:5] ;
assign n4243 =  ( n4213 ) == ( bv_3_4_n3659 )  ;
assign n4244 = acc[4:4] ;
assign n4245 =  ( n4213 ) == ( bv_3_3_n3517 )  ;
assign n4246 = acc[3:3] ;
assign n4247 =  ( n4213 ) == ( bv_3_2_n3664 )  ;
assign n4248 = acc[2:2] ;
assign n4249 =  ( n4213 ) == ( bv_3_1_n3667 )  ;
assign n4250 = acc[1:1] ;
assign n4251 = acc[0:0] ;
assign n4252 =  ( n4249 ) ? ( n4250 ) : ( n4251 ) ;
assign n4253 =  ( n4247 ) ? ( n4248 ) : ( n4252 ) ;
assign n4254 =  ( n4245 ) ? ( n4246 ) : ( n4253 ) ;
assign n4255 =  ( n4243 ) ? ( n4244 ) : ( n4254 ) ;
assign n4256 =  ( n4241 ) ? ( n4242 ) : ( n4255 ) ;
assign n4257 =  ( n4239 ) ? ( n4240 ) : ( n4256 ) ;
assign n4258 =  ( n4237 ) ? ( n4238 ) : ( n4257 ) ;
assign n4259 =  ( n4210 ) == ( bv_5_26_n3701 )  ;
assign n4260 =  ( n4213 ) == ( bv_3_7_n3557 )  ;
assign n4261 = n3705[7:7] ;
assign n4262 =  ( n4213 ) == ( bv_3_6_n3653 )  ;
assign n4263 = n3705[6:6] ;
assign n4264 =  ( n4213 ) == ( bv_3_5_n3656 )  ;
assign n4265 = n3705[5:5] ;
assign n4266 =  ( n4213 ) == ( bv_3_4_n3659 )  ;
assign n4267 = n3705[4:4] ;
assign n4268 =  ( n4213 ) == ( bv_3_3_n3517 )  ;
assign n4269 = n3705[3:3] ;
assign n4270 =  ( n4213 ) == ( bv_3_2_n3664 )  ;
assign n4271 = n3705[2:2] ;
assign n4272 =  ( n4213 ) == ( bv_3_1_n3667 )  ;
assign n4273 = n3705[1:1] ;
assign n4274 = n3705[0:0] ;
assign n4275 =  ( n4272 ) ? ( n4273 ) : ( n4274 ) ;
assign n4276 =  ( n4270 ) ? ( n4271 ) : ( n4275 ) ;
assign n4277 =  ( n4268 ) ? ( n4269 ) : ( n4276 ) ;
assign n4278 =  ( n4266 ) ? ( n4267 ) : ( n4277 ) ;
assign n4279 =  ( n4264 ) ? ( n4265 ) : ( n4278 ) ;
assign n4280 =  ( n4262 ) ? ( n4263 ) : ( n4279 ) ;
assign n4281 =  ( n4260 ) ? ( n4261 ) : ( n4280 ) ;
assign n4282 =  ( n4210 ) == ( bv_5_16_n3727 )  ;
assign n4283 =  ( n4213 ) == ( bv_3_7_n3557 )  ;
assign n4284 = p0[7:7] ;
assign n4285 =  ( n4213 ) == ( bv_3_6_n3653 )  ;
assign n4286 = p0[6:6] ;
assign n4287 =  ( n4213 ) == ( bv_3_5_n3656 )  ;
assign n4288 = p0[5:5] ;
assign n4289 =  ( n4213 ) == ( bv_3_4_n3659 )  ;
assign n4290 = p0[4:4] ;
assign n4291 =  ( n4213 ) == ( bv_3_3_n3517 )  ;
assign n4292 = p0[3:3] ;
assign n4293 =  ( n4213 ) == ( bv_3_2_n3664 )  ;
assign n4294 = p0[2:2] ;
assign n4295 =  ( n4213 ) == ( bv_3_1_n3667 )  ;
assign n4296 = p0[1:1] ;
assign n4297 = p0[0:0] ;
assign n4298 =  ( n4295 ) ? ( n4296 ) : ( n4297 ) ;
assign n4299 =  ( n4293 ) ? ( n4294 ) : ( n4298 ) ;
assign n4300 =  ( n4291 ) ? ( n4292 ) : ( n4299 ) ;
assign n4301 =  ( n4289 ) ? ( n4290 ) : ( n4300 ) ;
assign n4302 =  ( n4287 ) ? ( n4288 ) : ( n4301 ) ;
assign n4303 =  ( n4285 ) ? ( n4286 ) : ( n4302 ) ;
assign n4304 =  ( n4283 ) ? ( n4284 ) : ( n4303 ) ;
assign n4305 =  ( n4210 ) == ( bv_5_18_n3751 )  ;
assign n4306 =  ( n4213 ) == ( bv_3_7_n3557 )  ;
assign n4307 = p1[7:7] ;
assign n4308 =  ( n4213 ) == ( bv_3_6_n3653 )  ;
assign n4309 = p1[6:6] ;
assign n4310 =  ( n4213 ) == ( bv_3_5_n3656 )  ;
assign n4311 = p1[5:5] ;
assign n4312 =  ( n4213 ) == ( bv_3_4_n3659 )  ;
assign n4313 = p1[4:4] ;
assign n4314 =  ( n4213 ) == ( bv_3_3_n3517 )  ;
assign n4315 = p1[3:3] ;
assign n4316 =  ( n4213 ) == ( bv_3_2_n3664 )  ;
assign n4317 = p1[2:2] ;
assign n4318 =  ( n4213 ) == ( bv_3_1_n3667 )  ;
assign n4319 = p1[1:1] ;
assign n4320 = p1[0:0] ;
assign n4321 =  ( n4318 ) ? ( n4319 ) : ( n4320 ) ;
assign n4322 =  ( n4316 ) ? ( n4317 ) : ( n4321 ) ;
assign n4323 =  ( n4314 ) ? ( n4315 ) : ( n4322 ) ;
assign n4324 =  ( n4312 ) ? ( n4313 ) : ( n4323 ) ;
assign n4325 =  ( n4310 ) ? ( n4311 ) : ( n4324 ) ;
assign n4326 =  ( n4308 ) ? ( n4309 ) : ( n4325 ) ;
assign n4327 =  ( n4306 ) ? ( n4307 ) : ( n4326 ) ;
assign n4328 =  ( n4210 ) == ( bv_5_20_n3775 )  ;
assign n4329 =  ( n4213 ) == ( bv_3_7_n3557 )  ;
assign n4330 = p2[7:7] ;
assign n4331 =  ( n4213 ) == ( bv_3_6_n3653 )  ;
assign n4332 = p2[6:6] ;
assign n4333 =  ( n4213 ) == ( bv_3_5_n3656 )  ;
assign n4334 = p2[5:5] ;
assign n4335 =  ( n4213 ) == ( bv_3_4_n3659 )  ;
assign n4336 = p2[4:4] ;
assign n4337 =  ( n4213 ) == ( bv_3_3_n3517 )  ;
assign n4338 = p2[3:3] ;
assign n4339 =  ( n4213 ) == ( bv_3_2_n3664 )  ;
assign n4340 = p2[2:2] ;
assign n4341 =  ( n4213 ) == ( bv_3_1_n3667 )  ;
assign n4342 = p2[1:1] ;
assign n4343 = p2[0:0] ;
assign n4344 =  ( n4341 ) ? ( n4342 ) : ( n4343 ) ;
assign n4345 =  ( n4339 ) ? ( n4340 ) : ( n4344 ) ;
assign n4346 =  ( n4337 ) ? ( n4338 ) : ( n4345 ) ;
assign n4347 =  ( n4335 ) ? ( n4336 ) : ( n4346 ) ;
assign n4348 =  ( n4333 ) ? ( n4334 ) : ( n4347 ) ;
assign n4349 =  ( n4331 ) ? ( n4332 ) : ( n4348 ) ;
assign n4350 =  ( n4329 ) ? ( n4330 ) : ( n4349 ) ;
assign n4351 =  ( n4210 ) == ( bv_5_22_n3799 )  ;
assign n4352 =  ( n4213 ) == ( bv_3_7_n3557 )  ;
assign n4353 = p3[7:7] ;
assign n4354 =  ( n4213 ) == ( bv_3_6_n3653 )  ;
assign n4355 = p3[6:6] ;
assign n4356 =  ( n4213 ) == ( bv_3_5_n3656 )  ;
assign n4357 = p3[5:5] ;
assign n4358 =  ( n4213 ) == ( bv_3_4_n3659 )  ;
assign n4359 = p3[4:4] ;
assign n4360 =  ( n4213 ) == ( bv_3_3_n3517 )  ;
assign n4361 = p3[3:3] ;
assign n4362 =  ( n4213 ) == ( bv_3_2_n3664 )  ;
assign n4363 = p3[2:2] ;
assign n4364 =  ( n4213 ) == ( bv_3_1_n3667 )  ;
assign n4365 = p3[1:1] ;
assign n4366 = p3[0:0] ;
assign n4367 =  ( n4364 ) ? ( n4365 ) : ( n4366 ) ;
assign n4368 =  ( n4362 ) ? ( n4363 ) : ( n4367 ) ;
assign n4369 =  ( n4360 ) ? ( n4361 ) : ( n4368 ) ;
assign n4370 =  ( n4358 ) ? ( n4359 ) : ( n4369 ) ;
assign n4371 =  ( n4356 ) ? ( n4357 ) : ( n4370 ) ;
assign n4372 =  ( n4354 ) ? ( n4355 ) : ( n4371 ) ;
assign n4373 =  ( n4352 ) ? ( n4353 ) : ( n4372 ) ;
assign n4374 =  ( n4210 ) == ( bv_5_30_n3823 )  ;
assign n4375 =  ( n4213 ) == ( bv_3_7_n3557 )  ;
assign n4376 = b_reg[7:7] ;
assign n4377 =  ( n4213 ) == ( bv_3_6_n3653 )  ;
assign n4378 = b_reg[6:6] ;
assign n4379 =  ( n4213 ) == ( bv_3_5_n3656 )  ;
assign n4380 = b_reg[5:5] ;
assign n4381 =  ( n4213 ) == ( bv_3_4_n3659 )  ;
assign n4382 = b_reg[4:4] ;
assign n4383 =  ( n4213 ) == ( bv_3_3_n3517 )  ;
assign n4384 = b_reg[3:3] ;
assign n4385 =  ( n4213 ) == ( bv_3_2_n3664 )  ;
assign n4386 = b_reg[2:2] ;
assign n4387 =  ( n4213 ) == ( bv_3_1_n3667 )  ;
assign n4388 = b_reg[1:1] ;
assign n4389 = b_reg[0:0] ;
assign n4390 =  ( n4387 ) ? ( n4388 ) : ( n4389 ) ;
assign n4391 =  ( n4385 ) ? ( n4386 ) : ( n4390 ) ;
assign n4392 =  ( n4383 ) ? ( n4384 ) : ( n4391 ) ;
assign n4393 =  ( n4381 ) ? ( n4382 ) : ( n4392 ) ;
assign n4394 =  ( n4379 ) ? ( n4380 ) : ( n4393 ) ;
assign n4395 =  ( n4377 ) ? ( n4378 ) : ( n4394 ) ;
assign n4396 =  ( n4375 ) ? ( n4376 ) : ( n4395 ) ;
assign n4397 =  ( n4210 ) == ( bv_5_23_n3847 )  ;
assign n4398 =  ( n4213 ) == ( bv_3_7_n3557 )  ;
assign n4399 = ip[7:7] ;
assign n4400 =  ( n4213 ) == ( bv_3_6_n3653 )  ;
assign n4401 = ip[6:6] ;
assign n4402 =  ( n4213 ) == ( bv_3_5_n3656 )  ;
assign n4403 = ip[5:5] ;
assign n4404 =  ( n4213 ) == ( bv_3_4_n3659 )  ;
assign n4405 = ip[4:4] ;
assign n4406 =  ( n4213 ) == ( bv_3_3_n3517 )  ;
assign n4407 = ip[3:3] ;
assign n4408 =  ( n4213 ) == ( bv_3_2_n3664 )  ;
assign n4409 = ip[2:2] ;
assign n4410 =  ( n4213 ) == ( bv_3_1_n3667 )  ;
assign n4411 = ip[1:1] ;
assign n4412 = ip[0:0] ;
assign n4413 =  ( n4410 ) ? ( n4411 ) : ( n4412 ) ;
assign n4414 =  ( n4408 ) ? ( n4409 ) : ( n4413 ) ;
assign n4415 =  ( n4406 ) ? ( n4407 ) : ( n4414 ) ;
assign n4416 =  ( n4404 ) ? ( n4405 ) : ( n4415 ) ;
assign n4417 =  ( n4402 ) ? ( n4403 ) : ( n4416 ) ;
assign n4418 =  ( n4400 ) ? ( n4401 ) : ( n4417 ) ;
assign n4419 =  ( n4398 ) ? ( n4399 ) : ( n4418 ) ;
assign n4420 =  ( n4210 ) == ( bv_5_21_n3871 )  ;
assign n4421 =  ( n4213 ) == ( bv_3_7_n3557 )  ;
assign n4422 = ie[7:7] ;
assign n4423 =  ( n4213 ) == ( bv_3_6_n3653 )  ;
assign n4424 = ie[6:6] ;
assign n4425 =  ( n4213 ) == ( bv_3_5_n3656 )  ;
assign n4426 = ie[5:5] ;
assign n4427 =  ( n4213 ) == ( bv_3_4_n3659 )  ;
assign n4428 = ie[4:4] ;
assign n4429 =  ( n4213 ) == ( bv_3_3_n3517 )  ;
assign n4430 = ie[3:3] ;
assign n4431 =  ( n4213 ) == ( bv_3_2_n3664 )  ;
assign n4432 = ie[2:2] ;
assign n4433 =  ( n4213 ) == ( bv_3_1_n3667 )  ;
assign n4434 = ie[1:1] ;
assign n4435 = ie[0:0] ;
assign n4436 =  ( n4433 ) ? ( n4434 ) : ( n4435 ) ;
assign n4437 =  ( n4431 ) ? ( n4432 ) : ( n4436 ) ;
assign n4438 =  ( n4429 ) ? ( n4430 ) : ( n4437 ) ;
assign n4439 =  ( n4427 ) ? ( n4428 ) : ( n4438 ) ;
assign n4440 =  ( n4425 ) ? ( n4426 ) : ( n4439 ) ;
assign n4441 =  ( n4423 ) ? ( n4424 ) : ( n4440 ) ;
assign n4442 =  ( n4421 ) ? ( n4422 ) : ( n4441 ) ;
assign n4443 =  ( n4420 ) ? ( n4442 ) : ( bv_1_0_n53 ) ;
assign n4444 =  ( n4397 ) ? ( n4419 ) : ( n4443 ) ;
assign n4445 =  ( n4374 ) ? ( n4396 ) : ( n4444 ) ;
assign n4446 =  ( n4351 ) ? ( n4373 ) : ( n4445 ) ;
assign n4447 =  ( n4328 ) ? ( n4350 ) : ( n4446 ) ;
assign n4448 =  ( n4305 ) ? ( n4327 ) : ( n4447 ) ;
assign n4449 =  ( n4282 ) ? ( n4304 ) : ( n4448 ) ;
assign n4450 =  ( n4259 ) ? ( n4281 ) : ( n4449 ) ;
assign n4451 =  ( n4236 ) ? ( n4258 ) : ( n4450 ) ;
assign n4452 =  ( n4212 ) ? ( n4235 ) : ( n4451 ) ;
assign n4453 = rd_addr[7:3] ;
assign n4454 = wr_addr[7:3] ;
assign n4455 =  ( n4453 ) == ( n4454 )  ;
assign n4456 =  ( wr_bit_r ) == ( 1'b0 )  ;
assign n4457 =  ( n4455 ) & (n4456 )  ;
assign n4458 = wr_addr[2:0] ;
assign n4459 =  ( n4458 ) == ( bv_3_0_n46 )  ;
assign n4460 =  ( n4457 ) & (n4459 )  ;
assign n4461 =  ( n4460 ) & (n3932 )  ;
assign n4462 = rd_addr[2:0] ;
assign n4463 =  ( n4462 ) == ( bv_3_7_n3557 )  ;
assign n4464 = n3937[7:7] ;
assign n4465 =  ( n4462 ) == ( bv_3_6_n3653 )  ;
assign n4466 = n3937[6:6] ;
assign n4467 =  ( n4462 ) == ( bv_3_5_n3656 )  ;
assign n4468 = n3937[5:5] ;
assign n4469 =  ( n4462 ) == ( bv_3_4_n3659 )  ;
assign n4470 = n3937[4:4] ;
assign n4471 =  ( n4462 ) == ( bv_3_3_n3517 )  ;
assign n4472 = n3937[3:3] ;
assign n4473 =  ( n4462 ) == ( bv_3_2_n3664 )  ;
assign n4474 = n3937[2:2] ;
assign n4475 =  ( n4462 ) == ( bv_3_1_n3667 )  ;
assign n4476 = n3937[1:1] ;
assign n4477 = n3937[0:0] ;
assign n4478 =  ( n4475 ) ? ( n4476 ) : ( n4477 ) ;
assign n4479 =  ( n4473 ) ? ( n4474 ) : ( n4478 ) ;
assign n4480 =  ( n4471 ) ? ( n4472 ) : ( n4479 ) ;
assign n4481 =  ( n4469 ) ? ( n4470 ) : ( n4480 ) ;
assign n4482 =  ( n4467 ) ? ( n4468 ) : ( n4481 ) ;
assign n4483 =  ( n4465 ) ? ( n4466 ) : ( n4482 ) ;
assign n4484 =  ( n4463 ) ? ( n4464 ) : ( n4483 ) ;
assign n4485 =  ( wr_sfr ) == ( bv_2_1_n3501 )  ;
assign n4486 = rd_addr[7:3] ;
assign n4487 =  ( n4486 ) == ( bv_5_28_n3647 )  ;
assign n4488 =  ( n4485 ) & (n4487 )  ;
assign n4489 =  ( n4462 ) == ( bv_3_7_n3557 )  ;
assign n4490 = n3500[7:7] ;
assign n4491 =  ( n4462 ) == ( bv_3_6_n3653 )  ;
assign n4492 = n3500[6:6] ;
assign n4493 =  ( n4462 ) == ( bv_3_5_n3656 )  ;
assign n4494 = n3500[5:5] ;
assign n4495 =  ( n4462 ) == ( bv_3_4_n3659 )  ;
assign n4496 = n3500[4:4] ;
assign n4497 =  ( n4462 ) == ( bv_3_3_n3517 )  ;
assign n4498 = n3500[3:3] ;
assign n4499 =  ( n4462 ) == ( bv_3_2_n3664 )  ;
assign n4500 = n3500[2:2] ;
assign n4501 =  ( n4462 ) == ( bv_3_1_n3667 )  ;
assign n4502 = n3500[1:1] ;
assign n4503 = n3500[0:0] ;
assign n4504 =  ( n4501 ) ? ( n4502 ) : ( n4503 ) ;
assign n4505 =  ( n4499 ) ? ( n4500 ) : ( n4504 ) ;
assign n4506 =  ( n4497 ) ? ( n4498 ) : ( n4505 ) ;
assign n4507 =  ( n4495 ) ? ( n4496 ) : ( n4506 ) ;
assign n4508 =  ( n4493 ) ? ( n4494 ) : ( n4507 ) ;
assign n4509 =  ( n4491 ) ? ( n4492 ) : ( n4508 ) ;
assign n4510 =  ( n4489 ) ? ( n4490 ) : ( n4509 ) ;
assign n4511 =  ( rd_addr ) == ( wr_addr )  ;
assign n4512 =  ( n4511 ) & (wr_bit_r )  ;
assign n4513 =  ( n4512 ) & (n3932 )  ;
assign n4514 =  ( n4486 ) == ( bv_5_28_n3647 )  ;
assign n4515 =  ( n4462 ) == ( bv_3_7_n3557 )  ;
assign n4516 = acc[7:7] ;
assign n4517 =  ( n4462 ) == ( bv_3_6_n3653 )  ;
assign n4518 = acc[6:6] ;
assign n4519 =  ( n4462 ) == ( bv_3_5_n3656 )  ;
assign n4520 = acc[5:5] ;
assign n4521 =  ( n4462 ) == ( bv_3_4_n3659 )  ;
assign n4522 = acc[4:4] ;
assign n4523 =  ( n4462 ) == ( bv_3_3_n3517 )  ;
assign n4524 = acc[3:3] ;
assign n4525 =  ( n4462 ) == ( bv_3_2_n3664 )  ;
assign n4526 = acc[2:2] ;
assign n4527 =  ( n4462 ) == ( bv_3_1_n3667 )  ;
assign n4528 = acc[1:1] ;
assign n4529 = acc[0:0] ;
assign n4530 =  ( n4527 ) ? ( n4528 ) : ( n4529 ) ;
assign n4531 =  ( n4525 ) ? ( n4526 ) : ( n4530 ) ;
assign n4532 =  ( n4523 ) ? ( n4524 ) : ( n4531 ) ;
assign n4533 =  ( n4521 ) ? ( n4522 ) : ( n4532 ) ;
assign n4534 =  ( n4519 ) ? ( n4520 ) : ( n4533 ) ;
assign n4535 =  ( n4517 ) ? ( n4518 ) : ( n4534 ) ;
assign n4536 =  ( n4515 ) ? ( n4516 ) : ( n4535 ) ;
assign n4537 =  ( n4486 ) == ( bv_5_26_n3701 )  ;
assign n4538 =  ( n4462 ) == ( bv_3_7_n3557 )  ;
assign n4539 = n3705[7:7] ;
assign n4540 =  ( n4462 ) == ( bv_3_6_n3653 )  ;
assign n4541 = n3705[6:6] ;
assign n4542 =  ( n4462 ) == ( bv_3_5_n3656 )  ;
assign n4543 = n3705[5:5] ;
assign n4544 =  ( n4462 ) == ( bv_3_4_n3659 )  ;
assign n4545 = n3705[4:4] ;
assign n4546 =  ( n4462 ) == ( bv_3_3_n3517 )  ;
assign n4547 = n3705[3:3] ;
assign n4548 =  ( n4462 ) == ( bv_3_2_n3664 )  ;
assign n4549 = n3705[2:2] ;
assign n4550 =  ( n4462 ) == ( bv_3_1_n3667 )  ;
assign n4551 = n3705[1:1] ;
assign n4552 = n3705[0:0] ;
assign n4553 =  ( n4550 ) ? ( n4551 ) : ( n4552 ) ;
assign n4554 =  ( n4548 ) ? ( n4549 ) : ( n4553 ) ;
assign n4555 =  ( n4546 ) ? ( n4547 ) : ( n4554 ) ;
assign n4556 =  ( n4544 ) ? ( n4545 ) : ( n4555 ) ;
assign n4557 =  ( n4542 ) ? ( n4543 ) : ( n4556 ) ;
assign n4558 =  ( n4540 ) ? ( n4541 ) : ( n4557 ) ;
assign n4559 =  ( n4538 ) ? ( n4539 ) : ( n4558 ) ;
assign n4560 =  ( n4486 ) == ( bv_5_16_n3727 )  ;
assign n4561 =  ( n4462 ) == ( bv_3_7_n3557 )  ;
assign n4562 = p0[7:7] ;
assign n4563 =  ( n4462 ) == ( bv_3_6_n3653 )  ;
assign n4564 = p0[6:6] ;
assign n4565 =  ( n4462 ) == ( bv_3_5_n3656 )  ;
assign n4566 = p0[5:5] ;
assign n4567 =  ( n4462 ) == ( bv_3_4_n3659 )  ;
assign n4568 = p0[4:4] ;
assign n4569 =  ( n4462 ) == ( bv_3_3_n3517 )  ;
assign n4570 = p0[3:3] ;
assign n4571 =  ( n4462 ) == ( bv_3_2_n3664 )  ;
assign n4572 = p0[2:2] ;
assign n4573 =  ( n4462 ) == ( bv_3_1_n3667 )  ;
assign n4574 = p0[1:1] ;
assign n4575 = p0[0:0] ;
assign n4576 =  ( n4573 ) ? ( n4574 ) : ( n4575 ) ;
assign n4577 =  ( n4571 ) ? ( n4572 ) : ( n4576 ) ;
assign n4578 =  ( n4569 ) ? ( n4570 ) : ( n4577 ) ;
assign n4579 =  ( n4567 ) ? ( n4568 ) : ( n4578 ) ;
assign n4580 =  ( n4565 ) ? ( n4566 ) : ( n4579 ) ;
assign n4581 =  ( n4563 ) ? ( n4564 ) : ( n4580 ) ;
assign n4582 =  ( n4561 ) ? ( n4562 ) : ( n4581 ) ;
assign n4583 =  ( n4486 ) == ( bv_5_18_n3751 )  ;
assign n4584 =  ( n4462 ) == ( bv_3_7_n3557 )  ;
assign n4585 = p1[7:7] ;
assign n4586 =  ( n4462 ) == ( bv_3_6_n3653 )  ;
assign n4587 = p1[6:6] ;
assign n4588 =  ( n4462 ) == ( bv_3_5_n3656 )  ;
assign n4589 = p1[5:5] ;
assign n4590 =  ( n4462 ) == ( bv_3_4_n3659 )  ;
assign n4591 = p1[4:4] ;
assign n4592 =  ( n4462 ) == ( bv_3_3_n3517 )  ;
assign n4593 = p1[3:3] ;
assign n4594 =  ( n4462 ) == ( bv_3_2_n3664 )  ;
assign n4595 = p1[2:2] ;
assign n4596 =  ( n4462 ) == ( bv_3_1_n3667 )  ;
assign n4597 = p1[1:1] ;
assign n4598 = p1[0:0] ;
assign n4599 =  ( n4596 ) ? ( n4597 ) : ( n4598 ) ;
assign n4600 =  ( n4594 ) ? ( n4595 ) : ( n4599 ) ;
assign n4601 =  ( n4592 ) ? ( n4593 ) : ( n4600 ) ;
assign n4602 =  ( n4590 ) ? ( n4591 ) : ( n4601 ) ;
assign n4603 =  ( n4588 ) ? ( n4589 ) : ( n4602 ) ;
assign n4604 =  ( n4586 ) ? ( n4587 ) : ( n4603 ) ;
assign n4605 =  ( n4584 ) ? ( n4585 ) : ( n4604 ) ;
assign n4606 =  ( n4486 ) == ( bv_5_20_n3775 )  ;
assign n4607 =  ( n4462 ) == ( bv_3_7_n3557 )  ;
assign n4608 = p2[7:7] ;
assign n4609 =  ( n4462 ) == ( bv_3_6_n3653 )  ;
assign n4610 = p2[6:6] ;
assign n4611 =  ( n4462 ) == ( bv_3_5_n3656 )  ;
assign n4612 = p2[5:5] ;
assign n4613 =  ( n4462 ) == ( bv_3_4_n3659 )  ;
assign n4614 = p2[4:4] ;
assign n4615 =  ( n4462 ) == ( bv_3_3_n3517 )  ;
assign n4616 = p2[3:3] ;
assign n4617 =  ( n4462 ) == ( bv_3_2_n3664 )  ;
assign n4618 = p2[2:2] ;
assign n4619 =  ( n4462 ) == ( bv_3_1_n3667 )  ;
assign n4620 = p2[1:1] ;
assign n4621 = p2[0:0] ;
assign n4622 =  ( n4619 ) ? ( n4620 ) : ( n4621 ) ;
assign n4623 =  ( n4617 ) ? ( n4618 ) : ( n4622 ) ;
assign n4624 =  ( n4615 ) ? ( n4616 ) : ( n4623 ) ;
assign n4625 =  ( n4613 ) ? ( n4614 ) : ( n4624 ) ;
assign n4626 =  ( n4611 ) ? ( n4612 ) : ( n4625 ) ;
assign n4627 =  ( n4609 ) ? ( n4610 ) : ( n4626 ) ;
assign n4628 =  ( n4607 ) ? ( n4608 ) : ( n4627 ) ;
assign n4629 =  ( n4486 ) == ( bv_5_22_n3799 )  ;
assign n4630 =  ( n4462 ) == ( bv_3_7_n3557 )  ;
assign n4631 = p3[7:7] ;
assign n4632 =  ( n4462 ) == ( bv_3_6_n3653 )  ;
assign n4633 = p3[6:6] ;
assign n4634 =  ( n4462 ) == ( bv_3_5_n3656 )  ;
assign n4635 = p3[5:5] ;
assign n4636 =  ( n4462 ) == ( bv_3_4_n3659 )  ;
assign n4637 = p3[4:4] ;
assign n4638 =  ( n4462 ) == ( bv_3_3_n3517 )  ;
assign n4639 = p3[3:3] ;
assign n4640 =  ( n4462 ) == ( bv_3_2_n3664 )  ;
assign n4641 = p3[2:2] ;
assign n4642 =  ( n4462 ) == ( bv_3_1_n3667 )  ;
assign n4643 = p3[1:1] ;
assign n4644 = p3[0:0] ;
assign n4645 =  ( n4642 ) ? ( n4643 ) : ( n4644 ) ;
assign n4646 =  ( n4640 ) ? ( n4641 ) : ( n4645 ) ;
assign n4647 =  ( n4638 ) ? ( n4639 ) : ( n4646 ) ;
assign n4648 =  ( n4636 ) ? ( n4637 ) : ( n4647 ) ;
assign n4649 =  ( n4634 ) ? ( n4635 ) : ( n4648 ) ;
assign n4650 =  ( n4632 ) ? ( n4633 ) : ( n4649 ) ;
assign n4651 =  ( n4630 ) ? ( n4631 ) : ( n4650 ) ;
assign n4652 =  ( n4486 ) == ( bv_5_30_n3823 )  ;
assign n4653 =  ( n4462 ) == ( bv_3_7_n3557 )  ;
assign n4654 = b_reg[7:7] ;
assign n4655 =  ( n4462 ) == ( bv_3_6_n3653 )  ;
assign n4656 = b_reg[6:6] ;
assign n4657 =  ( n4462 ) == ( bv_3_5_n3656 )  ;
assign n4658 = b_reg[5:5] ;
assign n4659 =  ( n4462 ) == ( bv_3_4_n3659 )  ;
assign n4660 = b_reg[4:4] ;
assign n4661 =  ( n4462 ) == ( bv_3_3_n3517 )  ;
assign n4662 = b_reg[3:3] ;
assign n4663 =  ( n4462 ) == ( bv_3_2_n3664 )  ;
assign n4664 = b_reg[2:2] ;
assign n4665 =  ( n4462 ) == ( bv_3_1_n3667 )  ;
assign n4666 = b_reg[1:1] ;
assign n4667 = b_reg[0:0] ;
assign n4668 =  ( n4665 ) ? ( n4666 ) : ( n4667 ) ;
assign n4669 =  ( n4663 ) ? ( n4664 ) : ( n4668 ) ;
assign n4670 =  ( n4661 ) ? ( n4662 ) : ( n4669 ) ;
assign n4671 =  ( n4659 ) ? ( n4660 ) : ( n4670 ) ;
assign n4672 =  ( n4657 ) ? ( n4658 ) : ( n4671 ) ;
assign n4673 =  ( n4655 ) ? ( n4656 ) : ( n4672 ) ;
assign n4674 =  ( n4653 ) ? ( n4654 ) : ( n4673 ) ;
assign n4675 =  ( n4486 ) == ( bv_5_23_n3847 )  ;
assign n4676 =  ( n4462 ) == ( bv_3_7_n3557 )  ;
assign n4677 = ip[7:7] ;
assign n4678 =  ( n4462 ) == ( bv_3_6_n3653 )  ;
assign n4679 = ip[6:6] ;
assign n4680 =  ( n4462 ) == ( bv_3_5_n3656 )  ;
assign n4681 = ip[5:5] ;
assign n4682 =  ( n4462 ) == ( bv_3_4_n3659 )  ;
assign n4683 = ip[4:4] ;
assign n4684 =  ( n4462 ) == ( bv_3_3_n3517 )  ;
assign n4685 = ip[3:3] ;
assign n4686 =  ( n4462 ) == ( bv_3_2_n3664 )  ;
assign n4687 = ip[2:2] ;
assign n4688 =  ( n4462 ) == ( bv_3_1_n3667 )  ;
assign n4689 = ip[1:1] ;
assign n4690 = ip[0:0] ;
assign n4691 =  ( n4688 ) ? ( n4689 ) : ( n4690 ) ;
assign n4692 =  ( n4686 ) ? ( n4687 ) : ( n4691 ) ;
assign n4693 =  ( n4684 ) ? ( n4685 ) : ( n4692 ) ;
assign n4694 =  ( n4682 ) ? ( n4683 ) : ( n4693 ) ;
assign n4695 =  ( n4680 ) ? ( n4681 ) : ( n4694 ) ;
assign n4696 =  ( n4678 ) ? ( n4679 ) : ( n4695 ) ;
assign n4697 =  ( n4676 ) ? ( n4677 ) : ( n4696 ) ;
assign n4698 =  ( n4486 ) == ( bv_5_21_n3871 )  ;
assign n4699 =  ( n4462 ) == ( bv_3_7_n3557 )  ;
assign n4700 = ie[7:7] ;
assign n4701 =  ( n4462 ) == ( bv_3_6_n3653 )  ;
assign n4702 = ie[6:6] ;
assign n4703 =  ( n4462 ) == ( bv_3_5_n3656 )  ;
assign n4704 = ie[5:5] ;
assign n4705 =  ( n4462 ) == ( bv_3_4_n3659 )  ;
assign n4706 = ie[4:4] ;
assign n4707 =  ( n4462 ) == ( bv_3_3_n3517 )  ;
assign n4708 = ie[3:3] ;
assign n4709 =  ( n4462 ) == ( bv_3_2_n3664 )  ;
assign n4710 = ie[2:2] ;
assign n4711 =  ( n4462 ) == ( bv_3_1_n3667 )  ;
assign n4712 = ie[1:1] ;
assign n4713 = ie[0:0] ;
assign n4714 =  ( n4711 ) ? ( n4712 ) : ( n4713 ) ;
assign n4715 =  ( n4709 ) ? ( n4710 ) : ( n4714 ) ;
assign n4716 =  ( n4707 ) ? ( n4708 ) : ( n4715 ) ;
assign n4717 =  ( n4705 ) ? ( n4706 ) : ( n4716 ) ;
assign n4718 =  ( n4703 ) ? ( n4704 ) : ( n4717 ) ;
assign n4719 =  ( n4701 ) ? ( n4702 ) : ( n4718 ) ;
assign n4720 =  ( n4699 ) ? ( n4700 ) : ( n4719 ) ;
assign n4721 =  ( n4698 ) ? ( n4720 ) : ( bv_1_0_n53 ) ;
assign n4722 =  ( n4675 ) ? ( n4697 ) : ( n4721 ) ;
assign n4723 =  ( n4652 ) ? ( n4674 ) : ( n4722 ) ;
assign n4724 =  ( n4629 ) ? ( n4651 ) : ( n4723 ) ;
assign n4725 =  ( n4606 ) ? ( n4628 ) : ( n4724 ) ;
assign n4726 =  ( n4583 ) ? ( n4605 ) : ( n4725 ) ;
assign n4727 =  ( n4560 ) ? ( n4582 ) : ( n4726 ) ;
assign n4728 =  ( n4537 ) ? ( n4559 ) : ( n4727 ) ;
assign n4729 =  ( n4514 ) ? ( n4536 ) : ( n4728 ) ;
assign n4730 =  ( n4513 ) ? ( n3989 ) : ( n4729 ) ;
assign n4731 =  ( n4488 ) ? ( n4510 ) : ( n4730 ) ;
assign n4732 =  ( n4461 ) ? ( n4484 ) : ( n4731 ) ;
assign n4733 = rd_addr[7:7] ;
assign n4734 = rd_addr[7:7] ;
assign n4735 = rd_addr[7:7] ;
assign n4736 = rd_addr[7:7] ;
assign n4737 = rd_addr[7:7] ;
assign n4738 =  ( ram_rd_sel ) == ( bv_3_1_n3667 )  ;
assign n4739 =  ( ram_rd_sel ) == ( bv_3_1_n3667 )  ;
assign n4740 =  ( ram_rd_sel ) == ( bv_3_3_n3517 )  ;
assign n4741 =  ( n4739 ) | ( n4740 )  ;
assign n4742 =  ( ram_rd_sel ) == ( bv_3_1_n3667 )  ;
assign n4743 =  ( ram_rd_sel ) == ( bv_3_3_n3517 )  ;
assign n4744 =  ( n4742 ) | ( n4743 )  ;
assign n4745 =  ( ram_rd_sel ) == ( bv_3_1_n3667 )  ;
assign n4746 =  ( ram_rd_sel ) == ( bv_3_3_n3517 )  ;
assign n4747 =  ( n4745 ) | ( n4746 )  ;
assign n4748 =  ( ram_rd_sel ) == ( bv_3_1_n3667 )  ;
assign n4749 =  ( ram_rd_sel ) == ( bv_3_3_n3517 )  ;
assign n4750 =  ( n4748 ) | ( n4749 )  ;
assign n4751 =  ( wr_sfr ) == ( bv_2_2_n3505 )  ;
assign n4752 =  ( wr_sfr ) == ( bv_2_1_n3501 )  ;
assign n4753 =  ( src_sel1 ) == ( bv_3_1_n3667 )  ;
assign n4754 =  ( src_sel1 ) == ( bv_3_0_n46 )  ;
assign n4755 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n4756 =  ( rd_ind ) == ( 1'b0 )  ;
assign n4757 =  ( n4755 ) & (n4756 )  ;
assign n4758 =  ( n4757 ) ? ( sfr_rd_data ) : ( ram_rd_data ) ;
assign n4759 =  ( src_sel1 ) == ( bv_3_2_n3664 )  ;
assign n4760 =  ( src_sel1 ) == ( bv_3_4_n3659 )  ;
assign n4761 = pc[15:8] ;
assign n4762 =  ( src_sel1 ) == ( bv_3_5_n3656 )  ;
assign n4763 = pc[7:0] ;
assign n4764 =  ( src_sel1 ) == ( bv_3_3_n3517 )  ;
assign n4765 =  ( n4764 ) ? ( acc ) : ( bv_8_0_n69 ) ;
assign n4766 =  ( n4762 ) ? ( n4763 ) : ( n4765 ) ;
assign n4767 =  ( n4760 ) ? ( n4761 ) : ( n4766 ) ;
assign n4768 =  ( n4759 ) ? ( op3_reg ) : ( n4767 ) ;
assign n4769 =  ( n4754 ) ? ( n4758 ) : ( n4768 ) ;
assign n4770 =  ( n4753 ) ? ( op2_reg ) : ( n4769 ) ;
assign bv_2_0_n4771 = 2'h0 ;
assign n4772 =  ( src_sel2 ) == ( bv_2_0_n4771 )  ;
assign n4773 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n4774 =  ( rd_ind ) == ( 1'b0 )  ;
assign n4775 =  ( n4773 ) & (n4774 )  ;
assign n4776 =  ( n4775 ) ? ( sfr_rd_data ) : ( ram_rd_data ) ;
assign n4777 =  ( src_sel2 ) == ( bv_2_2_n3505 )  ;
assign n4778 =  ( src_sel2 ) == ( bv_2_3_n3495 )  ;
assign n4779 =  ( n4778 ) ? ( op2_reg ) : ( acc ) ;
assign n4780 =  ( n4777 ) ? ( bv_8_0_n69 ) : ( n4779 ) ;
assign n4781 =  ( n4772 ) ? ( n4776 ) : ( n4780 ) ;
assign n4782 =  ( n4770 ) & ( n4781 )  ;
assign n4783 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n4784 =  ( n4783 ) & (wr )  ;
assign n4785 =  ( n4784 ) ? ( n4782 ) : ( acc ) ;
assign n4786 =  ( n4752 ) ? ( n4782 ) : ( n4785 ) ;
assign n4787 =  ( n4751 ) ? ( bv_8_0_n69 ) : ( n4786 ) ;
assign n4788 =  ( wr_sfr ) == ( bv_2_2_n3505 )  ;
assign n4789 =  ( cy_sel ) == ( bv_2_0_n4771 )  ;
assign n4790 =  ( cy_sel ) == ( bv_2_1_n3501 )  ;
assign n4791 = psw[6:6] ;
assign n4792 =  ( cy_sel ) == ( bv_2_2_n3505 )  ;
assign n4793 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n4794 =  ( rd_ind ) == ( 1'b0 )  ;
assign n4795 =  ( n4793 ) & (n4794 )  ;
assign n4796 =  ( n4795 ) ? ( sfr_bit_rd_data ) : ( ram_bit_rd_data ) ;
assign n4797 =  ( n4792 ) ? ( n4796 ) : ( bv_1_1_n34 ) ;
assign n4798 =  ( n4790 ) ? ( n4791 ) : ( n4797 ) ;
assign n4799 =  ( n4789 ) ? ( bv_1_0_n53 ) : ( n4798 ) ;
assign n4800 =  ( n4799 ) == ( bv_1_1_n34 )  ;
assign n4801 =  ( src_sel2 ) == ( bv_2_0_n4771 )  ;
assign n4802 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n4803 =  ( rd_ind ) == ( 1'b0 )  ;
assign n4804 =  ( n4802 ) & (n4803 )  ;
assign n4805 =  ( n4804 ) ? ( sfr_rd_data ) : ( ram_rd_data ) ;
assign n4806 =  ( src_sel2 ) == ( bv_2_2_n3505 )  ;
assign n4807 =  ( src_sel2 ) == ( bv_2_3_n3495 )  ;
assign n4808 =  ( n4807 ) ? ( op2_reg ) : ( acc ) ;
assign n4809 =  ( n4806 ) ? ( bv_8_0_n69 ) : ( n4808 ) ;
assign n4810 =  ( n4801 ) ? ( n4805 ) : ( n4809 ) ;
assign n4811 =  ( src_sel1 ) == ( bv_3_1_n3667 )  ;
assign n4812 =  ( src_sel1 ) == ( bv_3_0_n46 )  ;
assign n4813 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n4814 =  ( rd_ind ) == ( 1'b0 )  ;
assign n4815 =  ( n4813 ) & (n4814 )  ;
assign n4816 =  ( n4815 ) ? ( sfr_rd_data ) : ( ram_rd_data ) ;
assign n4817 =  ( src_sel1 ) == ( bv_3_2_n3664 )  ;
assign n4818 =  ( src_sel1 ) == ( bv_3_4_n3659 )  ;
assign n4819 = pc[15:8] ;
assign n4820 =  ( src_sel1 ) == ( bv_3_5_n3656 )  ;
assign n4821 = pc[7:0] ;
assign n4822 =  ( src_sel1 ) == ( bv_3_3_n3517 )  ;
assign n4823 =  ( n4822 ) ? ( acc ) : ( bv_8_0_n69 ) ;
assign n4824 =  ( n4820 ) ? ( n4821 ) : ( n4823 ) ;
assign n4825 =  ( n4818 ) ? ( n4819 ) : ( n4824 ) ;
assign n4826 =  ( n4817 ) ? ( op3_reg ) : ( n4825 ) ;
assign n4827 =  ( n4812 ) ? ( n4816 ) : ( n4826 ) ;
assign n4828 =  ( n4811 ) ? ( op2_reg ) : ( n4827 ) ;
assign n4829 =  { ( n4810 ) , ( n4828 ) }  ;
assign bv_16_1_n4830 = 16'h1 ;
assign n4831 =  ( n4829 ) - ( bv_16_1_n4830 )  ;
assign n4832 = n4831[15:8] ;
assign n4833 =  { ( n4810 ) , ( n4828 ) }  ;
assign n4834 =  ( n4833 ) + ( bv_16_1_n4830 )  ;
assign n4835 = n4834[15:8] ;
assign n4836 =  ( n4800 ) ? ( n4832 ) : ( n4835 ) ;
assign n4837 =  ( wr_sfr ) == ( bv_2_1_n3501 )  ;
assign n4838 =  ( n4799 ) == ( bv_1_1_n34 )  ;
assign n4839 = n4831[7:0] ;
assign n4840 = n4834[7:0] ;
assign n4841 =  ( n4838 ) ? ( n4839 ) : ( n4840 ) ;
assign n4842 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n4843 =  ( n4842 ) & (wr )  ;
assign n4844 =  ( n4843 ) ? ( n4841 ) : ( acc ) ;
assign n4845 =  ( n4837 ) ? ( n4841 ) : ( n4844 ) ;
assign n4846 =  ( n4788 ) ? ( n4836 ) : ( n4845 ) ;
assign n4847 =  ( wr_sfr ) == ( bv_2_2_n3505 )  ;
assign n4848 =  ( wr_sfr ) == ( bv_2_1_n3501 )  ;
assign n4849 =  ( src_sel1 ) == ( bv_3_1_n3667 )  ;
assign n4850 =  ( src_sel1 ) == ( bv_3_0_n46 )  ;
assign n4851 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n4852 =  ( rd_ind ) == ( 1'b0 )  ;
assign n4853 =  ( n4851 ) & (n4852 )  ;
assign n4854 =  ( n4853 ) ? ( sfr_rd_data ) : ( ram_rd_data ) ;
assign n4855 =  ( src_sel1 ) == ( bv_3_2_n3664 )  ;
assign n4856 =  ( src_sel1 ) == ( bv_3_4_n3659 )  ;
assign n4857 = pc[15:8] ;
assign n4858 =  ( src_sel1 ) == ( bv_3_5_n3656 )  ;
assign n4859 = pc[7:0] ;
assign n4860 =  ( src_sel1 ) == ( bv_3_3_n3517 )  ;
assign n4861 =  ( n4860 ) ? ( acc ) : ( bv_8_0_n69 ) ;
assign n4862 =  ( n4858 ) ? ( n4859 ) : ( n4861 ) ;
assign n4863 =  ( n4856 ) ? ( n4857 ) : ( n4862 ) ;
assign n4864 =  ( n4855 ) ? ( op3_reg ) : ( n4863 ) ;
assign n4865 =  ( n4850 ) ? ( n4854 ) : ( n4864 ) ;
assign n4866 =  ( n4849 ) ? ( op2_reg ) : ( n4865 ) ;
assign n4867 = ~ ( n4866 ) ;
assign n4868 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n4869 =  ( n4868 ) & (wr )  ;
assign n4870 =  ( n4869 ) ? ( n4867 ) : ( acc ) ;
assign n4871 =  ( n4848 ) ? ( n4867 ) : ( n4870 ) ;
assign n4872 =  ( n4847 ) ? ( bv_8_0_n69 ) : ( n4871 ) ;
assign n4873 =  ( wr_sfr ) == ( bv_2_2_n3505 )  ;
assign n4874 =  ( wr_sfr ) == ( bv_2_1_n3501 )  ;
assign n4875 =  ( cy_sel ) == ( bv_2_0_n4771 )  ;
assign n4876 =  ( cy_sel ) == ( bv_2_1_n3501 )  ;
assign n4877 = psw[6:6] ;
assign n4878 =  ( cy_sel ) == ( bv_2_2_n3505 )  ;
assign n4879 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n4880 =  ( rd_ind ) == ( 1'b0 )  ;
assign n4881 =  ( n4879 ) & (n4880 )  ;
assign n4882 =  ( n4881 ) ? ( sfr_bit_rd_data ) : ( ram_bit_rd_data ) ;
assign n4883 =  ( n4878 ) ? ( n4882 ) : ( bv_1_1_n34 ) ;
assign n4884 =  ( n4876 ) ? ( n4877 ) : ( n4883 ) ;
assign n4885 =  ( n4875 ) ? ( bv_1_0_n53 ) : ( n4884 ) ;
assign n4886 =  ( n4885 ) == ( bv_1_1_n34 )  ;
assign n4887 = psw[5:5] ;
assign n4888 =  ( n4887 ) == ( bv_1_1_n34 )  ;
assign n4889 =  ( src_sel1 ) == ( bv_3_1_n3667 )  ;
assign n4890 =  ( src_sel1 ) == ( bv_3_0_n46 )  ;
assign n4891 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n4892 =  ( rd_ind ) == ( 1'b0 )  ;
assign n4893 =  ( n4891 ) & (n4892 )  ;
assign n4894 =  ( n4893 ) ? ( sfr_rd_data ) : ( ram_rd_data ) ;
assign n4895 =  ( src_sel1 ) == ( bv_3_2_n3664 )  ;
assign n4896 =  ( src_sel1 ) == ( bv_3_4_n3659 )  ;
assign n4897 = pc[15:8] ;
assign n4898 =  ( src_sel1 ) == ( bv_3_5_n3656 )  ;
assign n4899 = pc[7:0] ;
assign n4900 =  ( src_sel1 ) == ( bv_3_3_n3517 )  ;
assign n4901 =  ( n4900 ) ? ( acc ) : ( bv_8_0_n69 ) ;
assign n4902 =  ( n4898 ) ? ( n4899 ) : ( n4901 ) ;
assign n4903 =  ( n4896 ) ? ( n4897 ) : ( n4902 ) ;
assign n4904 =  ( n4895 ) ? ( op3_reg ) : ( n4903 ) ;
assign n4905 =  ( n4890 ) ? ( n4894 ) : ( n4904 ) ;
assign n4906 =  ( n4889 ) ? ( op2_reg ) : ( n4905 ) ;
assign n4907 = n4906[3:0] ;
assign n4908 =  ( n4907 ) > ( bv_4_9_n14 )  ;
assign n4909 =  ( n4888 ) | ( n4908 )  ;
assign n4910 = n4906[3:0] ;
assign n4911 =  { ( bv_1_0_n53 ) , ( n4910 ) }  ;
assign bv_5_6_n4912 = 5'h6 ;
assign n4913 =  ( n4911 ) + ( bv_5_6_n4912 )  ;
assign n4914 = n4906[3:0] ;
assign n4915 =  { ( bv_1_0_n53 ) , ( n4914 ) }  ;
assign n4916 =  ( n4909 ) ? ( n4913 ) : ( n4915 ) ;
assign n4917 = n4916[4:4] ;
assign n4918 =  ( n4917 ) == ( bv_1_1_n34 )  ;
assign n4919 =  ( n4886 ) | ( n4918 )  ;
assign n4920 = n4906[7:4] ;
assign n4921 =  ( n4920 ) > ( bv_4_9_n14 )  ;
assign n4922 =  ( n4919 ) | ( n4921 )  ;
assign n4923 = n4906[7:4] ;
assign n4924 =  { ( n4885 ) , ( n4923 ) }  ;
assign n4925 =  ( n4924 ) + ( bv_5_6_n4912 )  ;
assign n4926 = n4916[4:4] ;
assign n4927 =  { ( bv_4_0_n30 ) , ( n4926 ) }  ;
assign n4928 =  ( n4925 ) + ( n4927 )  ;
assign n4929 = n4906[7:4] ;
assign n4930 =  { ( n4885 ) , ( n4929 ) }  ;
assign n4931 = n4916[4:4] ;
assign n4932 =  { ( bv_4_0_n30 ) , ( n4931 ) }  ;
assign n4933 =  ( n4930 ) + ( n4932 )  ;
assign n4934 =  ( n4922 ) ? ( n4928 ) : ( n4933 ) ;
assign n4935 = n4934[3:0] ;
assign n4936 = n4916[3:0] ;
assign n4937 =  { ( n4935 ) , ( n4936 ) }  ;
assign n4938 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n4939 =  ( n4938 ) & (wr )  ;
assign n4940 =  ( n4939 ) ? ( n4937 ) : ( acc ) ;
assign n4941 =  ( n4874 ) ? ( n4937 ) : ( n4940 ) ;
assign n4942 =  ( n4873 ) ? ( bv_8_0_n69 ) : ( n4941 ) ;
assign n4943 =  ( wr_sfr ) == ( bv_2_2_n3505 )  ;
assign n4945 = nondet_mul_des2_n4944 ;
assign n4946 =  ( wr_sfr ) == ( bv_2_1_n3501 )  ;
assign n4948 = nondet_mul_des1_n4947 ;
assign n4949 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n4950 =  ( n4949 ) & (wr )  ;
assign n4951 =  ( n4950 ) ? ( n4948 ) : ( acc ) ;
assign n4952 =  ( n4946 ) ? ( n4948 ) : ( n4951 ) ;
assign n4953 =  ( n4943 ) ? ( n4945 ) : ( n4952 ) ;
assign n4954 =  ( wr_sfr ) == ( bv_2_2_n3505 )  ;
assign n4956 = nondet_div_des2_n4955 ;
assign n4957 =  ( wr_sfr ) == ( bv_2_1_n3501 )  ;
assign n4959 = nondet_div_des1_n4958 ;
assign n4960 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n4961 =  ( n4960 ) & (wr )  ;
assign n4962 =  ( n4961 ) ? ( n4959 ) : ( acc ) ;
assign n4963 =  ( n4957 ) ? ( n4959 ) : ( n4962 ) ;
assign n4964 =  ( n4954 ) ? ( n4956 ) : ( n4963 ) ;
assign n4965 =  ( wr_sfr ) == ( bv_2_2_n3505 )  ;
assign n4966 =  ( wr_sfr ) == ( bv_2_1_n3501 )  ;
assign n4967 =  ( src_sel1 ) == ( bv_3_1_n3667 )  ;
assign n4968 =  ( src_sel1 ) == ( bv_3_0_n46 )  ;
assign n4969 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n4970 =  ( rd_ind ) == ( 1'b0 )  ;
assign n4971 =  ( n4969 ) & (n4970 )  ;
assign n4972 =  ( n4971 ) ? ( sfr_rd_data ) : ( ram_rd_data ) ;
assign n4973 =  ( src_sel1 ) == ( bv_3_2_n3664 )  ;
assign n4974 =  ( src_sel1 ) == ( bv_3_4_n3659 )  ;
assign n4975 = pc[15:8] ;
assign n4976 =  ( src_sel1 ) == ( bv_3_5_n3656 )  ;
assign n4977 = pc[7:0] ;
assign n4978 =  ( src_sel1 ) == ( bv_3_3_n3517 )  ;
assign n4979 =  ( n4978 ) ? ( acc ) : ( bv_8_0_n69 ) ;
assign n4980 =  ( n4976 ) ? ( n4977 ) : ( n4979 ) ;
assign n4981 =  ( n4974 ) ? ( n4975 ) : ( n4980 ) ;
assign n4982 =  ( n4973 ) ? ( op3_reg ) : ( n4981 ) ;
assign n4983 =  ( n4968 ) ? ( n4972 ) : ( n4982 ) ;
assign n4984 =  ( n4967 ) ? ( op2_reg ) : ( n4983 ) ;
assign n4985 = n4984[7:7] ;
assign n4986 =  { ( bv_1_1_n34 ) , ( n4985 ) }  ;
assign n4987 =  ( src_sel2 ) == ( bv_2_0_n4771 )  ;
assign n4988 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n4989 =  ( rd_ind ) == ( 1'b0 )  ;
assign n4990 =  ( n4988 ) & (n4989 )  ;
assign n4991 =  ( n4990 ) ? ( sfr_rd_data ) : ( ram_rd_data ) ;
assign n4992 =  ( src_sel2 ) == ( bv_2_2_n3505 )  ;
assign n4993 =  ( src_sel2 ) == ( bv_2_3_n3495 )  ;
assign n4994 =  ( n4993 ) ? ( op2_reg ) : ( acc ) ;
assign n4995 =  ( n4992 ) ? ( bv_8_0_n69 ) : ( n4994 ) ;
assign n4996 =  ( n4987 ) ? ( n4991 ) : ( n4995 ) ;
assign n4997 = n4996[7:7] ;
assign n4998 =  { ( bv_1_0_n53 ) , ( n4997 ) }  ;
assign n4999 =  ( n4986 ) - ( n4998 )  ;
assign n5000 = n4984[6:4] ;
assign n5001 =  { ( bv_1_1_n34 ) , ( n5000 ) }  ;
assign n5002 = n4996[6:4] ;
assign n5003 =  { ( bv_1_0_n53 ) , ( n5002 ) }  ;
assign n5004 =  ( n5001 ) - ( n5003 )  ;
assign n5005 = n4984[3:0] ;
assign n5006 =  { ( bv_1_1_n34 ) , ( n5005 ) }  ;
assign n5007 = n4996[3:0] ;
assign n5008 =  { ( bv_1_0_n53 ) , ( n5007 ) }  ;
assign n5009 =  ( n5006 ) - ( n5008 )  ;
assign n5010 =  ( cy_sel ) == ( bv_2_0_n4771 )  ;
assign n5011 =  ( cy_sel ) == ( bv_2_1_n3501 )  ;
assign n5012 = psw[6:6] ;
assign n5013 =  ( cy_sel ) == ( bv_2_2_n3505 )  ;
assign n5014 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n5015 =  ( rd_ind ) == ( 1'b0 )  ;
assign n5016 =  ( n5014 ) & (n5015 )  ;
assign n5017 =  ( n5016 ) ? ( sfr_bit_rd_data ) : ( ram_bit_rd_data ) ;
assign n5018 =  ( n5013 ) ? ( n5017 ) : ( bv_1_1_n34 ) ;
assign n5019 =  ( n5011 ) ? ( n5012 ) : ( n5018 ) ;
assign n5020 =  ( n5010 ) ? ( bv_1_0_n53 ) : ( n5019 ) ;
assign n5021 =  { ( bv_4_0_n30 ) , ( n5020 ) }  ;
assign n5022 =  ( n5009 ) - ( n5021 )  ;
assign n5023 = n5022[4:4] ;
assign n5024 = ~ ( n5023 ) ;
assign n5025 =  { ( bv_3_0_n46 ) , ( n5024 ) }  ;
assign n5026 =  ( n5004 ) - ( n5025 )  ;
assign n5027 = n5026[3:3] ;
assign n5028 = ~ ( n5027 ) ;
assign n5029 =  { ( bv_1_0_n53 ) , ( n5028 ) }  ;
assign n5030 =  ( n4999 ) - ( n5029 )  ;
assign n5031 = n5030[0:0] ;
assign n5032 = n5026[2:0] ;
assign n5033 =  { ( n5031 ) , ( n5032 ) }  ;
assign n5034 = n5022[3:0] ;
assign n5035 =  { ( n5033 ) , ( n5034 ) }  ;
assign n5036 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n5037 =  ( n5036 ) & (wr )  ;
assign n5038 =  ( n5037 ) ? ( n5035 ) : ( acc ) ;
assign n5039 =  ( n4966 ) ? ( n5035 ) : ( n5038 ) ;
assign n5040 =  ( n4965 ) ? ( bv_8_0_n69 ) : ( n5039 ) ;
assign n5041 =  ( wr_sfr ) == ( bv_2_2_n3505 )  ;
assign n5042 =  ( wr_sfr ) == ( bv_2_1_n3501 )  ;
assign n5043 =  ( src_sel1 ) == ( bv_3_1_n3667 )  ;
assign n5044 =  ( src_sel1 ) == ( bv_3_0_n46 )  ;
assign n5045 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n5046 =  ( rd_ind ) == ( 1'b0 )  ;
assign n5047 =  ( n5045 ) & (n5046 )  ;
assign n5048 =  ( n5047 ) ? ( sfr_rd_data ) : ( ram_rd_data ) ;
assign n5049 =  ( src_sel1 ) == ( bv_3_2_n3664 )  ;
assign n5050 =  ( src_sel1 ) == ( bv_3_4_n3659 )  ;
assign n5051 = pc[15:8] ;
assign n5052 =  ( src_sel1 ) == ( bv_3_5_n3656 )  ;
assign n5053 = pc[7:0] ;
assign n5054 =  ( src_sel1 ) == ( bv_3_3_n3517 )  ;
assign n5055 =  ( n5054 ) ? ( acc ) : ( bv_8_0_n69 ) ;
assign n5056 =  ( n5052 ) ? ( n5053 ) : ( n5055 ) ;
assign n5057 =  ( n5050 ) ? ( n5051 ) : ( n5056 ) ;
assign n5058 =  ( n5049 ) ? ( op3_reg ) : ( n5057 ) ;
assign n5059 =  ( n5044 ) ? ( n5048 ) : ( n5058 ) ;
assign n5060 =  ( n5043 ) ? ( op2_reg ) : ( n5059 ) ;
assign n5061 =  ( src_sel2 ) == ( bv_2_0_n4771 )  ;
assign n5062 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n5063 =  ( rd_ind ) == ( 1'b0 )  ;
assign n5064 =  ( n5062 ) & (n5063 )  ;
assign n5065 =  ( n5064 ) ? ( sfr_rd_data ) : ( ram_rd_data ) ;
assign n5066 =  ( src_sel2 ) == ( bv_2_2_n3505 )  ;
assign n5067 =  ( src_sel2 ) == ( bv_2_3_n3495 )  ;
assign n5068 =  ( n5067 ) ? ( op2_reg ) : ( acc ) ;
assign n5069 =  ( n5066 ) ? ( bv_8_0_n69 ) : ( n5068 ) ;
assign n5070 =  ( n5061 ) ? ( n5065 ) : ( n5069 ) ;
assign n5071 =  ( n5060 ) | ( n5070 )  ;
assign n5072 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n5073 =  ( n5072 ) & (wr )  ;
assign n5074 =  ( n5073 ) ? ( n5071 ) : ( acc ) ;
assign n5075 =  ( n5042 ) ? ( n5071 ) : ( n5074 ) ;
assign n5076 =  ( n5041 ) ? ( bv_8_0_n69 ) : ( n5075 ) ;
assign n5077 =  ( wr_sfr ) == ( bv_2_2_n3505 )  ;
assign n5078 =  ( wr_sfr ) == ( bv_2_1_n3501 )  ;
assign n5079 =  ( src_sel1 ) == ( bv_3_1_n3667 )  ;
assign n5080 =  ( src_sel1 ) == ( bv_3_0_n46 )  ;
assign n5081 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n5082 =  ( rd_ind ) == ( 1'b0 )  ;
assign n5083 =  ( n5081 ) & (n5082 )  ;
assign n5084 =  ( n5083 ) ? ( sfr_rd_data ) : ( ram_rd_data ) ;
assign n5085 =  ( src_sel1 ) == ( bv_3_2_n3664 )  ;
assign n5086 =  ( src_sel1 ) == ( bv_3_4_n3659 )  ;
assign n5087 = pc[15:8] ;
assign n5088 =  ( src_sel1 ) == ( bv_3_5_n3656 )  ;
assign n5089 = pc[7:0] ;
assign n5090 =  ( src_sel1 ) == ( bv_3_3_n3517 )  ;
assign n5091 =  ( n5090 ) ? ( acc ) : ( bv_8_0_n69 ) ;
assign n5092 =  ( n5088 ) ? ( n5089 ) : ( n5091 ) ;
assign n5093 =  ( n5086 ) ? ( n5087 ) : ( n5092 ) ;
assign n5094 =  ( n5085 ) ? ( op3_reg ) : ( n5093 ) ;
assign n5095 =  ( n5080 ) ? ( n5084 ) : ( n5094 ) ;
assign n5096 =  ( n5079 ) ? ( op2_reg ) : ( n5095 ) ;
assign n5097 = n5096[6:0] ;
assign n5098 = n5096[7:7] ;
assign n5099 =  { ( n5097 ) , ( n5098 ) }  ;
assign n5100 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n5101 =  ( n5100 ) & (wr )  ;
assign n5102 =  ( n5101 ) ? ( n5099 ) : ( acc ) ;
assign n5103 =  ( n5078 ) ? ( n5099 ) : ( n5102 ) ;
assign n5104 =  ( n5077 ) ? ( bv_8_0_n69 ) : ( n5103 ) ;
assign n5105 =  ( wr_sfr ) == ( bv_2_2_n3505 )  ;
assign n5106 =  ( src_sel1 ) == ( bv_3_1_n3667 )  ;
assign n5107 =  ( src_sel1 ) == ( bv_3_0_n46 )  ;
assign n5108 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n5109 =  ( rd_ind ) == ( 1'b0 )  ;
assign n5110 =  ( n5108 ) & (n5109 )  ;
assign n5111 =  ( n5110 ) ? ( sfr_rd_data ) : ( ram_rd_data ) ;
assign n5112 =  ( src_sel1 ) == ( bv_3_2_n3664 )  ;
assign n5113 =  ( src_sel1 ) == ( bv_3_4_n3659 )  ;
assign n5114 = pc[15:8] ;
assign n5115 =  ( src_sel1 ) == ( bv_3_5_n3656 )  ;
assign n5116 = pc[7:0] ;
assign n5117 =  ( src_sel1 ) == ( bv_3_3_n3517 )  ;
assign n5118 =  ( n5117 ) ? ( acc ) : ( bv_8_0_n69 ) ;
assign n5119 =  ( n5115 ) ? ( n5116 ) : ( n5118 ) ;
assign n5120 =  ( n5113 ) ? ( n5114 ) : ( n5119 ) ;
assign n5121 =  ( n5112 ) ? ( op3_reg ) : ( n5120 ) ;
assign n5122 =  ( n5107 ) ? ( n5111 ) : ( n5121 ) ;
assign n5123 =  ( n5106 ) ? ( op2_reg ) : ( n5122 ) ;
assign n5124 = n5123[3:0] ;
assign n5125 = n5123[7:4] ;
assign n5126 =  { ( n5124 ) , ( n5125 ) }  ;
assign n5127 =  ( wr_sfr ) == ( bv_2_1_n3501 )  ;
assign n5128 = n5123[6:0] ;
assign n5129 =  ( cy_sel ) == ( bv_2_0_n4771 )  ;
assign n5130 =  ( cy_sel ) == ( bv_2_1_n3501 )  ;
assign n5131 = psw[6:6] ;
assign n5132 =  ( cy_sel ) == ( bv_2_2_n3505 )  ;
assign n5133 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n5134 =  ( rd_ind ) == ( 1'b0 )  ;
assign n5135 =  ( n5133 ) & (n5134 )  ;
assign n5136 =  ( n5135 ) ? ( sfr_bit_rd_data ) : ( ram_bit_rd_data ) ;
assign n5137 =  ( n5132 ) ? ( n5136 ) : ( bv_1_1_n34 ) ;
assign n5138 =  ( n5130 ) ? ( n5131 ) : ( n5137 ) ;
assign n5139 =  ( n5129 ) ? ( bv_1_0_n53 ) : ( n5138 ) ;
assign n5140 =  { ( n5128 ) , ( n5139 ) }  ;
assign n5141 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n5142 =  ( n5141 ) & (wr )  ;
assign n5143 =  ( n5142 ) ? ( n5140 ) : ( acc ) ;
assign n5144 =  ( n5127 ) ? ( n5140 ) : ( n5143 ) ;
assign n5145 =  ( n5105 ) ? ( n5126 ) : ( n5144 ) ;
assign n5146 =  ( wr_sfr ) == ( bv_2_2_n3505 )  ;
assign n5147 =  ( wr_sfr ) == ( bv_2_1_n3501 )  ;
assign n5148 =  ( src_sel1 ) == ( bv_3_1_n3667 )  ;
assign n5149 =  ( src_sel1 ) == ( bv_3_0_n46 )  ;
assign n5150 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n5151 =  ( rd_ind ) == ( 1'b0 )  ;
assign n5152 =  ( n5150 ) & (n5151 )  ;
assign n5153 =  ( n5152 ) ? ( sfr_rd_data ) : ( ram_rd_data ) ;
assign n5154 =  ( src_sel1 ) == ( bv_3_2_n3664 )  ;
assign n5155 =  ( src_sel1 ) == ( bv_3_4_n3659 )  ;
assign n5156 = pc[15:8] ;
assign n5157 =  ( src_sel1 ) == ( bv_3_5_n3656 )  ;
assign n5158 = pc[7:0] ;
assign n5159 =  ( src_sel1 ) == ( bv_3_3_n3517 )  ;
assign n5160 =  ( n5159 ) ? ( acc ) : ( bv_8_0_n69 ) ;
assign n5161 =  ( n5157 ) ? ( n5158 ) : ( n5160 ) ;
assign n5162 =  ( n5155 ) ? ( n5156 ) : ( n5161 ) ;
assign n5163 =  ( n5154 ) ? ( op3_reg ) : ( n5162 ) ;
assign n5164 =  ( n5149 ) ? ( n5153 ) : ( n5163 ) ;
assign n5165 =  ( n5148 ) ? ( op2_reg ) : ( n5164 ) ;
assign n5166 = n5165[0:0] ;
assign n5167 = n5165[7:1] ;
assign n5168 =  { ( n5166 ) , ( n5167 ) }  ;
assign n5169 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n5170 =  ( n5169 ) & (wr )  ;
assign n5171 =  ( n5170 ) ? ( n5168 ) : ( acc ) ;
assign n5172 =  ( n5147 ) ? ( n5168 ) : ( n5171 ) ;
assign n5173 =  ( n5146 ) ? ( bv_8_0_n69 ) : ( n5172 ) ;
assign n5174 =  ( wr_sfr ) == ( bv_2_2_n3505 )  ;
assign n5175 =  ( wr_sfr ) == ( bv_2_1_n3501 )  ;
assign n5176 =  ( cy_sel ) == ( bv_2_0_n4771 )  ;
assign n5177 =  ( cy_sel ) == ( bv_2_1_n3501 )  ;
assign n5178 = psw[6:6] ;
assign n5179 =  ( cy_sel ) == ( bv_2_2_n3505 )  ;
assign n5180 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n5181 =  ( rd_ind ) == ( 1'b0 )  ;
assign n5182 =  ( n5180 ) & (n5181 )  ;
assign n5183 =  ( n5182 ) ? ( sfr_bit_rd_data ) : ( ram_bit_rd_data ) ;
assign n5184 =  ( n5179 ) ? ( n5183 ) : ( bv_1_1_n34 ) ;
assign n5185 =  ( n5177 ) ? ( n5178 ) : ( n5184 ) ;
assign n5186 =  ( n5176 ) ? ( bv_1_0_n53 ) : ( n5185 ) ;
assign n5187 =  ( src_sel1 ) == ( bv_3_1_n3667 )  ;
assign n5188 =  ( src_sel1 ) == ( bv_3_0_n46 )  ;
assign n5189 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n5190 =  ( rd_ind ) == ( 1'b0 )  ;
assign n5191 =  ( n5189 ) & (n5190 )  ;
assign n5192 =  ( n5191 ) ? ( sfr_rd_data ) : ( ram_rd_data ) ;
assign n5193 =  ( src_sel1 ) == ( bv_3_2_n3664 )  ;
assign n5194 =  ( src_sel1 ) == ( bv_3_4_n3659 )  ;
assign n5195 = pc[15:8] ;
assign n5196 =  ( src_sel1 ) == ( bv_3_5_n3656 )  ;
assign n5197 = pc[7:0] ;
assign n5198 =  ( src_sel1 ) == ( bv_3_3_n3517 )  ;
assign n5199 =  ( n5198 ) ? ( acc ) : ( bv_8_0_n69 ) ;
assign n5200 =  ( n5196 ) ? ( n5197 ) : ( n5199 ) ;
assign n5201 =  ( n5194 ) ? ( n5195 ) : ( n5200 ) ;
assign n5202 =  ( n5193 ) ? ( op3_reg ) : ( n5201 ) ;
assign n5203 =  ( n5188 ) ? ( n5192 ) : ( n5202 ) ;
assign n5204 =  ( n5187 ) ? ( op2_reg ) : ( n5203 ) ;
assign n5205 = n5204[7:1] ;
assign n5206 =  { ( n5186 ) , ( n5205 ) }  ;
assign n5207 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n5208 =  ( n5207 ) & (wr )  ;
assign n5209 =  ( n5208 ) ? ( n5206 ) : ( acc ) ;
assign n5210 =  ( n5175 ) ? ( n5206 ) : ( n5209 ) ;
assign n5211 =  ( n5174 ) ? ( bv_8_0_n69 ) : ( n5210 ) ;
assign n5212 =  ( wr_sfr ) == ( bv_2_2_n3505 )  ;
assign n5213 =  ( cy_sel ) == ( bv_2_0_n4771 )  ;
assign n5214 =  ( cy_sel ) == ( bv_2_1_n3501 )  ;
assign n5215 = psw[6:6] ;
assign n5216 =  ( cy_sel ) == ( bv_2_2_n3505 )  ;
assign n5217 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n5218 =  ( rd_ind ) == ( 1'b0 )  ;
assign n5219 =  ( n5217 ) & (n5218 )  ;
assign n5220 =  ( n5219 ) ? ( sfr_bit_rd_data ) : ( ram_bit_rd_data ) ;
assign n5221 =  ( n5216 ) ? ( n5220 ) : ( bv_1_1_n34 ) ;
assign n5222 =  ( n5214 ) ? ( n5215 ) : ( n5221 ) ;
assign n5223 =  ( n5213 ) ? ( bv_1_0_n53 ) : ( n5222 ) ;
assign n5224 =  ( n5223 ) == ( bv_1_1_n34 )  ;
assign n5225 =  ( src_sel1 ) == ( bv_3_1_n3667 )  ;
assign n5226 =  ( src_sel1 ) == ( bv_3_0_n46 )  ;
assign n5227 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n5228 =  ( rd_ind ) == ( 1'b0 )  ;
assign n5229 =  ( n5227 ) & (n5228 )  ;
assign n5230 =  ( n5229 ) ? ( sfr_rd_data ) : ( ram_rd_data ) ;
assign n5231 =  ( src_sel1 ) == ( bv_3_2_n3664 )  ;
assign n5232 =  ( src_sel1 ) == ( bv_3_4_n3659 )  ;
assign n5233 = pc[15:8] ;
assign n5234 =  ( src_sel1 ) == ( bv_3_5_n3656 )  ;
assign n5235 = pc[7:0] ;
assign n5236 =  ( src_sel1 ) == ( bv_3_3_n3517 )  ;
assign n5237 =  ( n5236 ) ? ( acc ) : ( bv_8_0_n69 ) ;
assign n5238 =  ( n5234 ) ? ( n5235 ) : ( n5237 ) ;
assign n5239 =  ( n5232 ) ? ( n5233 ) : ( n5238 ) ;
assign n5240 =  ( n5231 ) ? ( op3_reg ) : ( n5239 ) ;
assign n5241 =  ( n5226 ) ? ( n5230 ) : ( n5240 ) ;
assign n5242 =  ( n5225 ) ? ( op2_reg ) : ( n5241 ) ;
assign n5243 =  ( src_sel2 ) == ( bv_2_0_n4771 )  ;
assign n5244 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n5245 =  ( rd_ind ) == ( 1'b0 )  ;
assign n5246 =  ( n5244 ) & (n5245 )  ;
assign n5247 =  ( n5246 ) ? ( sfr_rd_data ) : ( ram_rd_data ) ;
assign n5248 =  ( src_sel2 ) == ( bv_2_2_n3505 )  ;
assign n5249 =  ( src_sel2 ) == ( bv_2_3_n3495 )  ;
assign n5250 =  ( n5249 ) ? ( op2_reg ) : ( acc ) ;
assign n5251 =  ( n5248 ) ? ( bv_8_0_n69 ) : ( n5250 ) ;
assign n5252 =  ( n5243 ) ? ( n5247 ) : ( n5251 ) ;
assign n5253 = n5252[7:4] ;
assign n5254 = n5242[3:0] ;
assign n5255 =  { ( n5253 ) , ( n5254 ) }  ;
assign n5256 =  ( n5224 ) ? ( n5242 ) : ( n5255 ) ;
assign n5257 =  ( wr_sfr ) == ( bv_2_1_n3501 )  ;
assign n5258 =  ( n5223 ) == ( bv_1_1_n34 )  ;
assign n5259 = n5242[7:4] ;
assign n5260 = n5252[3:0] ;
assign n5261 =  { ( n5259 ) , ( n5260 ) }  ;
assign n5262 =  ( n5258 ) ? ( n5252 ) : ( n5261 ) ;
assign n5263 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n5264 =  ( n5263 ) & (wr )  ;
assign n5265 =  ( n5264 ) ? ( n5262 ) : ( acc ) ;
assign n5266 =  ( n5257 ) ? ( n5262 ) : ( n5265 ) ;
assign n5267 =  ( n5212 ) ? ( n5256 ) : ( n5266 ) ;
assign n5268 =  ( wr_sfr ) == ( bv_2_2_n3505 )  ;
assign n5269 =  ( wr_sfr ) == ( bv_2_1_n3501 )  ;
assign n5270 =  ( src_sel1 ) == ( bv_3_1_n3667 )  ;
assign n5271 =  ( src_sel1 ) == ( bv_3_0_n46 )  ;
assign n5272 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n5273 =  ( rd_ind ) == ( 1'b0 )  ;
assign n5274 =  ( n5272 ) & (n5273 )  ;
assign n5275 =  ( n5274 ) ? ( sfr_rd_data ) : ( ram_rd_data ) ;
assign n5276 =  ( src_sel1 ) == ( bv_3_2_n3664 )  ;
assign n5277 =  ( src_sel1 ) == ( bv_3_4_n3659 )  ;
assign n5278 = pc[15:8] ;
assign n5279 =  ( src_sel1 ) == ( bv_3_5_n3656 )  ;
assign n5280 = pc[7:0] ;
assign n5281 =  ( src_sel1 ) == ( bv_3_3_n3517 )  ;
assign n5282 =  ( n5281 ) ? ( acc ) : ( bv_8_0_n69 ) ;
assign n5283 =  ( n5279 ) ? ( n5280 ) : ( n5282 ) ;
assign n5284 =  ( n5277 ) ? ( n5278 ) : ( n5283 ) ;
assign n5285 =  ( n5276 ) ? ( op3_reg ) : ( n5284 ) ;
assign n5286 =  ( n5271 ) ? ( n5275 ) : ( n5285 ) ;
assign n5287 =  ( n5270 ) ? ( op2_reg ) : ( n5286 ) ;
assign n5288 =  ( src_sel2 ) == ( bv_2_0_n4771 )  ;
assign n5289 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n5290 =  ( rd_ind ) == ( 1'b0 )  ;
assign n5291 =  ( n5289 ) & (n5290 )  ;
assign n5292 =  ( n5291 ) ? ( sfr_rd_data ) : ( ram_rd_data ) ;
assign n5293 =  ( src_sel2 ) == ( bv_2_2_n3505 )  ;
assign n5294 =  ( src_sel2 ) == ( bv_2_3_n3495 )  ;
assign n5295 =  ( n5294 ) ? ( op2_reg ) : ( acc ) ;
assign n5296 =  ( n5293 ) ? ( bv_8_0_n69 ) : ( n5295 ) ;
assign n5297 =  ( n5288 ) ? ( n5292 ) : ( n5296 ) ;
assign n5298 =  ( n5287 ) ^ ( n5297 )  ;
assign n5299 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n5300 =  ( n5299 ) & (wr )  ;
assign n5301 =  ( n5300 ) ? ( n5298 ) : ( acc ) ;
assign n5302 =  ( n5269 ) ? ( n5298 ) : ( n5301 ) ;
assign n5303 =  ( n5268 ) ? ( bv_8_0_n69 ) : ( n5302 ) ;
assign n5304 =  ( wr_sfr ) == ( bv_2_2_n3505 )  ;
assign n5305 =  ( src_sel3 ) == ( 1'b1 )  ;
assign n5306 = pc[15:8] ;
assign n5307 =  ( n5305 ) ? ( n5306 ) : ( dptr_hi ) ;
assign n5308 =  ( src_sel1 ) == ( bv_3_1_n3667 )  ;
assign n5309 =  ( src_sel1 ) == ( bv_3_0_n46 )  ;
assign n5310 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n5311 =  ( rd_ind ) == ( 1'b0 )  ;
assign n5312 =  ( n5310 ) & (n5311 )  ;
assign n5313 =  ( n5312 ) ? ( sfr_rd_data ) : ( ram_rd_data ) ;
assign n5314 =  ( src_sel1 ) == ( bv_3_2_n3664 )  ;
assign n5315 =  ( src_sel1 ) == ( bv_3_4_n3659 )  ;
assign n5316 = pc[15:8] ;
assign n5317 =  ( src_sel1 ) == ( bv_3_5_n3656 )  ;
assign n5318 = pc[7:0] ;
assign n5319 =  ( src_sel1 ) == ( bv_3_3_n3517 )  ;
assign n5320 =  ( n5319 ) ? ( acc ) : ( bv_8_0_n69 ) ;
assign n5321 =  ( n5317 ) ? ( n5318 ) : ( n5320 ) ;
assign n5322 =  ( n5315 ) ? ( n5316 ) : ( n5321 ) ;
assign n5323 =  ( n5314 ) ? ( op3_reg ) : ( n5322 ) ;
assign n5324 =  ( n5309 ) ? ( n5313 ) : ( n5323 ) ;
assign n5325 =  ( n5308 ) ? ( op2_reg ) : ( n5324 ) ;
assign n5326 = n5325[7:7] ;
assign n5327 =  { ( bv_1_0_n53 ) , ( n5326 ) }  ;
assign n5328 =  ( src_sel2 ) == ( bv_2_0_n4771 )  ;
assign n5329 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n5330 =  ( rd_ind ) == ( 1'b0 )  ;
assign n5331 =  ( n5329 ) & (n5330 )  ;
assign n5332 =  ( n5331 ) ? ( sfr_rd_data ) : ( ram_rd_data ) ;
assign n5333 =  ( src_sel2 ) == ( bv_2_2_n3505 )  ;
assign n5334 =  ( src_sel2 ) == ( bv_2_3_n3495 )  ;
assign n5335 =  ( n5334 ) ? ( op2_reg ) : ( acc ) ;
assign n5336 =  ( n5333 ) ? ( bv_8_0_n69 ) : ( n5335 ) ;
assign n5337 =  ( n5328 ) ? ( n5332 ) : ( n5336 ) ;
assign n5338 = n5337[7:7] ;
assign n5339 =  { ( bv_1_0_n53 ) , ( n5338 ) }  ;
assign n5340 =  ( n5327 ) + ( n5339 )  ;
assign n5341 = n5325[6:4] ;
assign n5342 =  { ( bv_1_0_n53 ) , ( n5341 ) }  ;
assign n5343 = n5337[6:4] ;
assign n5344 =  { ( bv_1_0_n53 ) , ( n5343 ) }  ;
assign n5345 =  ( n5342 ) + ( n5344 )  ;
assign n5346 = n5325[3:0] ;
assign n5347 =  { ( bv_1_0_n53 ) , ( n5346 ) }  ;
assign n5348 = n5337[3:0] ;
assign n5349 =  { ( bv_1_0_n53 ) , ( n5348 ) }  ;
assign n5350 =  ( n5347 ) + ( n5349 )  ;
assign n5351 =  ( cy_sel ) == ( bv_2_0_n4771 )  ;
assign n5352 =  ( cy_sel ) == ( bv_2_1_n3501 )  ;
assign n5353 = psw[6:6] ;
assign n5354 =  ( cy_sel ) == ( bv_2_2_n3505 )  ;
assign n5355 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n5356 =  ( rd_ind ) == ( 1'b0 )  ;
assign n5357 =  ( n5355 ) & (n5356 )  ;
assign n5358 =  ( n5357 ) ? ( sfr_bit_rd_data ) : ( ram_bit_rd_data ) ;
assign n5359 =  ( n5354 ) ? ( n5358 ) : ( bv_1_1_n34 ) ;
assign n5360 =  ( n5352 ) ? ( n5353 ) : ( n5359 ) ;
assign n5361 =  ( n5351 ) ? ( bv_1_0_n53 ) : ( n5360 ) ;
assign n5362 =  { ( bv_4_0_n30 ) , ( n5361 ) }  ;
assign n5363 =  ( n5350 ) + ( n5362 )  ;
assign n5364 = n5363[4:4] ;
assign n5365 =  { ( bv_3_0_n46 ) , ( n5364 ) }  ;
assign n5366 =  ( n5345 ) + ( n5365 )  ;
assign n5367 = n5366[3:3] ;
assign n5368 =  { ( bv_1_0_n53 ) , ( n5367 ) }  ;
assign n5369 =  ( n5340 ) + ( n5368 )  ;
assign n5370 = n5369[1:1] ;
assign n5371 =  { ( bv_7_0_n3520 ) , ( n5370 ) }  ;
assign n5372 =  ( n5307 ) + ( n5371 )  ;
assign n5373 =  ( wr_sfr ) == ( bv_2_1_n3501 )  ;
assign n5374 = n5369[0:0] ;
assign n5375 = n5366[2:0] ;
assign n5376 =  { ( n5374 ) , ( n5375 ) }  ;
assign n5377 = n5363[3:0] ;
assign n5378 =  { ( n5376 ) , ( n5377 ) }  ;
assign n5379 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n5380 =  ( n5379 ) & (wr )  ;
assign n5381 =  ( n5380 ) ? ( n5378 ) : ( acc ) ;
assign n5382 =  ( n5373 ) ? ( n5378 ) : ( n5381 ) ;
assign n5383 =  ( n5304 ) ? ( n5372 ) : ( n5382 ) ;
assign n5384 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n5385 =  ( n5384 ) & (wr )  ;
assign n5386 =  ( n5385 ) ? ( n4782 ) : ( b_reg ) ;
assign n5387 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n5388 =  ( n5387 ) & (wr )  ;
assign n5389 =  ( n5388 ) ? ( n4841 ) : ( b_reg ) ;
assign n5390 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n5391 =  ( n5390 ) & (wr )  ;
assign n5392 =  ( n5391 ) ? ( n4867 ) : ( b_reg ) ;
assign n5393 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n5394 =  ( n5393 ) & (wr )  ;
assign n5395 =  ( n5394 ) ? ( n4937 ) : ( b_reg ) ;
assign n5396 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n5397 =  ( n5396 ) & (wr )  ;
assign n5398 =  ( n5397 ) ? ( n4948 ) : ( b_reg ) ;
assign n5399 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n5400 =  ( n5399 ) & (wr )  ;
assign n5401 =  ( n5400 ) ? ( n4959 ) : ( b_reg ) ;
assign n5402 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n5403 =  ( n5402 ) & (wr )  ;
assign n5404 =  ( n5403 ) ? ( n5035 ) : ( b_reg ) ;
assign n5405 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n5406 =  ( n5405 ) & (wr )  ;
assign n5407 =  ( n5406 ) ? ( n5071 ) : ( b_reg ) ;
assign n5408 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n5409 =  ( n5408 ) & (wr )  ;
assign n5410 =  ( n5409 ) ? ( n5099 ) : ( b_reg ) ;
assign n5411 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n5412 =  ( n5411 ) & (wr )  ;
assign n5413 =  ( n5412 ) ? ( n5140 ) : ( b_reg ) ;
assign n5414 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n5415 =  ( n5414 ) & (wr )  ;
assign n5416 =  ( n5415 ) ? ( n5168 ) : ( b_reg ) ;
assign n5417 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n5418 =  ( n5417 ) & (wr )  ;
assign n5419 =  ( n5418 ) ? ( n5206 ) : ( b_reg ) ;
assign n5420 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n5421 =  ( n5420 ) & (wr )  ;
assign n5422 =  ( n5421 ) ? ( n5262 ) : ( b_reg ) ;
assign n5423 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n5424 =  ( n5423 ) & (wr )  ;
assign n5425 =  ( n5424 ) ? ( n5298 ) : ( b_reg ) ;
assign n5426 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n5427 =  ( n5426 ) & (wr )  ;
assign n5428 =  ( n5427 ) ? ( n5378 ) : ( b_reg ) ;
assign n5429 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n5430 =  ( n5429 ) & (wr )  ;
assign n5431 =  ( ram_wr_sel ) == ( bv_3_3_n3517 )  ;
assign n5432 =  ( sp ) + ( bv_8_1_n71 )  ;
assign n5433 =  ( pop ) ? ( bv_1_1_n34 ) : ( bv_1_0_n53 ) ;
assign n5434 =  { ( bv_7_0_n3520 ) , ( n5433 ) }  ;
assign n5435 =  ( sp ) - ( n5434 )  ;
assign n5436 =  ( n5431 ) ? ( n5432 ) : ( n5435 ) ;
assign n5437 =  ( n5430 ) ? ( n4782 ) : ( n5436 ) ;
assign n5438 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n5439 =  ( n5438 ) & (wr )  ;
assign n5440 =  ( ram_wr_sel ) == ( bv_3_3_n3517 )  ;
assign n5441 =  ( sp ) + ( bv_8_1_n71 )  ;
assign n5442 =  ( pop ) ? ( bv_1_1_n34 ) : ( bv_1_0_n53 ) ;
assign n5443 =  { ( bv_7_0_n3520 ) , ( n5442 ) }  ;
assign n5444 =  ( sp ) - ( n5443 )  ;
assign n5445 =  ( n5440 ) ? ( n5441 ) : ( n5444 ) ;
assign n5446 =  ( n5439 ) ? ( n4841 ) : ( n5445 ) ;
assign n5447 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n5448 =  ( n5447 ) & (wr )  ;
assign n5449 = ~ ( n4866 ) ;
assign n5450 =  ( ram_wr_sel ) == ( bv_3_3_n3517 )  ;
assign n5451 =  ( sp ) + ( bv_8_1_n71 )  ;
assign n5452 =  ( pop ) ? ( bv_1_1_n34 ) : ( bv_1_0_n53 ) ;
assign n5453 =  { ( bv_7_0_n3520 ) , ( n5452 ) }  ;
assign n5454 =  ( sp ) - ( n5453 )  ;
assign n5455 =  ( n5450 ) ? ( n5451 ) : ( n5454 ) ;
assign n5456 =  ( n5448 ) ? ( n5449 ) : ( n5455 ) ;
assign n5457 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n5458 =  ( n5457 ) & (wr )  ;
assign n5459 =  ( ram_wr_sel ) == ( bv_3_3_n3517 )  ;
assign n5460 =  ( sp ) + ( bv_8_1_n71 )  ;
assign n5461 =  ( pop ) ? ( bv_1_1_n34 ) : ( bv_1_0_n53 ) ;
assign n5462 =  { ( bv_7_0_n3520 ) , ( n5461 ) }  ;
assign n5463 =  ( sp ) - ( n5462 )  ;
assign n5464 =  ( n5459 ) ? ( n5460 ) : ( n5463 ) ;
assign n5465 =  ( n5458 ) ? ( n4906 ) : ( n5464 ) ;
assign n5466 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n5467 =  ( n5466 ) & (wr )  ;
assign n5468 =  ( src_sel1 ) == ( bv_3_1_n3667 )  ;
assign n5469 =  ( src_sel1 ) == ( bv_3_0_n46 )  ;
assign n5470 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n5471 =  ( rd_ind ) == ( 1'b0 )  ;
assign n5472 =  ( n5470 ) & (n5471 )  ;
assign n5473 =  ( n5472 ) ? ( sfr_rd_data ) : ( ram_rd_data ) ;
assign n5474 =  ( src_sel1 ) == ( bv_3_2_n3664 )  ;
assign n5475 =  ( src_sel1 ) == ( bv_3_4_n3659 )  ;
assign n5476 = pc[15:8] ;
assign n5477 =  ( src_sel1 ) == ( bv_3_5_n3656 )  ;
assign n5478 = pc[7:0] ;
assign n5479 =  ( src_sel1 ) == ( bv_3_3_n3517 )  ;
assign n5480 =  ( n5479 ) ? ( acc ) : ( bv_8_0_n69 ) ;
assign n5481 =  ( n5477 ) ? ( n5478 ) : ( n5480 ) ;
assign n5482 =  ( n5475 ) ? ( n5476 ) : ( n5481 ) ;
assign n5483 =  ( n5474 ) ? ( op3_reg ) : ( n5482 ) ;
assign n5484 =  ( n5469 ) ? ( n5473 ) : ( n5483 ) ;
assign n5485 =  ( n5468 ) ? ( op2_reg ) : ( n5484 ) ;
assign n5486 =  ( ram_wr_sel ) == ( bv_3_3_n3517 )  ;
assign n5487 =  ( sp ) + ( bv_8_1_n71 )  ;
assign n5488 =  ( pop ) ? ( bv_1_1_n34 ) : ( bv_1_0_n53 ) ;
assign n5489 =  { ( bv_7_0_n3520 ) , ( n5488 ) }  ;
assign n5490 =  ( sp ) - ( n5489 )  ;
assign n5491 =  ( n5486 ) ? ( n5487 ) : ( n5490 ) ;
assign n5492 =  ( n5467 ) ? ( n5485 ) : ( n5491 ) ;
assign n5493 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n5494 =  ( n5493 ) & (wr )  ;
assign n5495 =  ( src_sel1 ) == ( bv_3_1_n3667 )  ;
assign n5496 =  ( src_sel1 ) == ( bv_3_0_n46 )  ;
assign n5497 =  ( rd_addr_r ) == ( 1'b1 )  ;
assign n5498 =  ( rd_ind ) == ( 1'b0 )  ;
assign n5499 =  ( n5497 ) & (n5498 )  ;
assign n5500 =  ( n5499 ) ? ( sfr_rd_data ) : ( ram_rd_data ) ;
assign n5501 =  ( src_sel1 ) == ( bv_3_2_n3664 )  ;
assign n5502 =  ( src_sel1 ) == ( bv_3_4_n3659 )  ;
assign n5503 = pc[15:8] ;
assign n5504 =  ( src_sel1 ) == ( bv_3_5_n3656 )  ;
assign n5505 = pc[7:0] ;
assign n5506 =  ( src_sel1 ) == ( bv_3_3_n3517 )  ;
assign n5507 =  ( n5506 ) ? ( acc ) : ( bv_8_0_n69 ) ;
assign n5508 =  ( n5504 ) ? ( n5505 ) : ( n5507 ) ;
assign n5509 =  ( n5502 ) ? ( n5503 ) : ( n5508 ) ;
assign n5510 =  ( n5501 ) ? ( op3_reg ) : ( n5509 ) ;
assign n5511 =  ( n5496 ) ? ( n5500 ) : ( n5510 ) ;
assign n5512 =  ( n5495 ) ? ( op2_reg ) : ( n5511 ) ;
assign n5513 =  ( ram_wr_sel ) == ( bv_3_3_n3517 )  ;
assign n5514 =  ( sp ) + ( bv_8_1_n71 )  ;
assign n5515 =  ( pop ) ? ( bv_1_1_n34 ) : ( bv_1_0_n53 ) ;
assign n5516 =  { ( bv_7_0_n3520 ) , ( n5515 ) }  ;
assign n5517 =  ( sp ) - ( n5516 )  ;
assign n5518 =  ( n5513 ) ? ( n5514 ) : ( n5517 ) ;
assign n5519 =  ( n5494 ) ? ( n5512 ) : ( n5518 ) ;
assign n5520 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n5521 =  ( n5520 ) & (wr )  ;
assign n5522 =  ( ram_wr_sel ) == ( bv_3_3_n3517 )  ;
assign n5523 =  ( sp ) + ( bv_8_1_n71 )  ;
assign n5524 =  ( pop ) ? ( bv_1_1_n34 ) : ( bv_1_0_n53 ) ;
assign n5525 =  { ( bv_7_0_n3520 ) , ( n5524 ) }  ;
assign n5526 =  ( sp ) - ( n5525 )  ;
assign n5527 =  ( n5522 ) ? ( n5523 ) : ( n5526 ) ;
assign n5528 =  ( n5521 ) ? ( bv_8_0_n69 ) : ( n5527 ) ;
assign n5529 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n5530 =  ( n5529 ) & (wr )  ;
assign n5531 =  ( ram_wr_sel ) == ( bv_3_3_n3517 )  ;
assign n5532 =  ( sp ) + ( bv_8_1_n71 )  ;
assign n5533 =  ( pop ) ? ( bv_1_1_n34 ) : ( bv_1_0_n53 ) ;
assign n5534 =  { ( bv_7_0_n3520 ) , ( n5533 ) }  ;
assign n5535 =  ( sp ) - ( n5534 )  ;
assign n5536 =  ( n5531 ) ? ( n5532 ) : ( n5535 ) ;
assign n5537 =  ( n5530 ) ? ( n5071 ) : ( n5536 ) ;
assign n5538 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n5539 =  ( n5538 ) & (wr )  ;
assign n5540 =  ( ram_wr_sel ) == ( bv_3_3_n3517 )  ;
assign n5541 =  ( sp ) + ( bv_8_1_n71 )  ;
assign n5542 =  ( pop ) ? ( bv_1_1_n34 ) : ( bv_1_0_n53 ) ;
assign n5543 =  { ( bv_7_0_n3520 ) , ( n5542 ) }  ;
assign n5544 =  ( sp ) - ( n5543 )  ;
assign n5545 =  ( n5540 ) ? ( n5541 ) : ( n5544 ) ;
assign n5546 =  ( n5539 ) ? ( n5096 ) : ( n5545 ) ;
assign n5547 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n5548 =  ( n5547 ) & (wr )  ;
assign n5549 =  ( ram_wr_sel ) == ( bv_3_3_n3517 )  ;
assign n5550 =  ( sp ) + ( bv_8_1_n71 )  ;
assign n5551 =  ( pop ) ? ( bv_1_1_n34 ) : ( bv_1_0_n53 ) ;
assign n5552 =  { ( bv_7_0_n3520 ) , ( n5551 ) }  ;
assign n5553 =  ( sp ) - ( n5552 )  ;
assign n5554 =  ( n5549 ) ? ( n5550 ) : ( n5553 ) ;
assign n5555 =  ( n5548 ) ? ( n5123 ) : ( n5554 ) ;
assign n5556 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n5557 =  ( n5556 ) & (wr )  ;
assign n5558 =  ( ram_wr_sel ) == ( bv_3_3_n3517 )  ;
assign n5559 =  ( sp ) + ( bv_8_1_n71 )  ;
assign n5560 =  ( pop ) ? ( bv_1_1_n34 ) : ( bv_1_0_n53 ) ;
assign n5561 =  { ( bv_7_0_n3520 ) , ( n5560 ) }  ;
assign n5562 =  ( sp ) - ( n5561 )  ;
assign n5563 =  ( n5558 ) ? ( n5559 ) : ( n5562 ) ;
assign n5564 =  ( n5557 ) ? ( n5165 ) : ( n5563 ) ;
assign n5565 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n5566 =  ( n5565 ) & (wr )  ;
assign n5567 =  ( ram_wr_sel ) == ( bv_3_3_n3517 )  ;
assign n5568 =  ( sp ) + ( bv_8_1_n71 )  ;
assign n5569 =  ( pop ) ? ( bv_1_1_n34 ) : ( bv_1_0_n53 ) ;
assign n5570 =  { ( bv_7_0_n3520 ) , ( n5569 ) }  ;
assign n5571 =  ( sp ) - ( n5570 )  ;
assign n5572 =  ( n5567 ) ? ( n5568 ) : ( n5571 ) ;
assign n5573 =  ( n5566 ) ? ( n5204 ) : ( n5572 ) ;
assign n5574 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n5575 =  ( n5574 ) & (wr )  ;
assign n5576 =  ( ram_wr_sel ) == ( bv_3_3_n3517 )  ;
assign n5577 =  ( sp ) + ( bv_8_1_n71 )  ;
assign n5578 =  ( pop ) ? ( bv_1_1_n34 ) : ( bv_1_0_n53 ) ;
assign n5579 =  { ( bv_7_0_n3520 ) , ( n5578 ) }  ;
assign n5580 =  ( sp ) - ( n5579 )  ;
assign n5581 =  ( n5576 ) ? ( n5577 ) : ( n5580 ) ;
assign n5582 =  ( n5575 ) ? ( n5298 ) : ( n5581 ) ;
assign n5583 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n5584 =  ( n5583 ) & (wr )  ;
assign n5585 =  ( ram_wr_sel ) == ( bv_3_3_n3517 )  ;
assign n5586 =  ( sp ) + ( bv_8_1_n71 )  ;
assign n5587 =  ( pop ) ? ( bv_1_1_n34 ) : ( bv_1_0_n53 ) ;
assign n5588 =  { ( bv_7_0_n3520 ) , ( n5587 ) }  ;
assign n5589 =  ( sp ) - ( n5588 )  ;
assign n5590 =  ( n5585 ) ? ( n5586 ) : ( n5589 ) ;
assign n5591 =  ( n5584 ) ? ( n5325 ) : ( n5590 ) ;
assign n5592 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5593 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n5594 =  ( n5593 ) & (wr )  ;
assign n5595 =  ( n5594 ) ? ( n4782 ) : ( dptr_hi ) ;
assign n5596 =  ( n5592 ) ? ( bv_8_0_n69 ) : ( n5595 ) ;
assign n5597 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5598 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n5599 =  ( n5598 ) & (wr )  ;
assign n5600 =  ( n5599 ) ? ( n4841 ) : ( dptr_hi ) ;
assign n5601 =  ( n5597 ) ? ( n4836 ) : ( n5600 ) ;
assign n5602 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5603 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n5604 =  ( n5603 ) & (wr )  ;
assign n5605 =  ( n5604 ) ? ( n4867 ) : ( dptr_hi ) ;
assign n5606 =  ( n5602 ) ? ( bv_8_0_n69 ) : ( n5605 ) ;
assign n5607 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5608 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n5609 =  ( n5608 ) & (wr )  ;
assign n5610 =  ( n5609 ) ? ( n4937 ) : ( dptr_hi ) ;
assign n5611 =  ( n5607 ) ? ( bv_8_0_n69 ) : ( n5610 ) ;
assign n5612 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5613 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n5614 =  ( n5613 ) & (wr )  ;
assign n5615 =  ( n5614 ) ? ( n4948 ) : ( dptr_hi ) ;
assign n5616 =  ( n5612 ) ? ( n4945 ) : ( n5615 ) ;
assign n5617 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5618 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n5619 =  ( n5618 ) & (wr )  ;
assign n5620 =  ( n5619 ) ? ( n4959 ) : ( dptr_hi ) ;
assign n5621 =  ( n5617 ) ? ( n4956 ) : ( n5620 ) ;
assign n5622 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5623 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n5624 =  ( n5623 ) & (wr )  ;
assign n5625 =  ( n5624 ) ? ( n5035 ) : ( dptr_hi ) ;
assign n5626 =  ( n5622 ) ? ( bv_8_0_n69 ) : ( n5625 ) ;
assign n5627 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5628 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n5629 =  ( n5628 ) & (wr )  ;
assign n5630 =  ( n5629 ) ? ( n5071 ) : ( dptr_hi ) ;
assign n5631 =  ( n5627 ) ? ( bv_8_0_n69 ) : ( n5630 ) ;
assign n5632 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5633 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n5634 =  ( n5633 ) & (wr )  ;
assign n5635 =  ( n5634 ) ? ( n5099 ) : ( dptr_hi ) ;
assign n5636 =  ( n5632 ) ? ( bv_8_0_n69 ) : ( n5635 ) ;
assign n5637 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5638 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n5639 =  ( n5638 ) & (wr )  ;
assign n5640 =  ( n5639 ) ? ( n5140 ) : ( dptr_hi ) ;
assign n5641 =  ( n5637 ) ? ( n5126 ) : ( n5640 ) ;
assign n5642 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5643 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n5644 =  ( n5643 ) & (wr )  ;
assign n5645 =  ( n5644 ) ? ( n5168 ) : ( dptr_hi ) ;
assign n5646 =  ( n5642 ) ? ( bv_8_0_n69 ) : ( n5645 ) ;
assign n5647 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5648 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n5649 =  ( n5648 ) & (wr )  ;
assign n5650 =  ( n5649 ) ? ( n5206 ) : ( dptr_hi ) ;
assign n5651 =  ( n5647 ) ? ( bv_8_0_n69 ) : ( n5650 ) ;
assign n5652 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5653 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n5654 =  ( n5653 ) & (wr )  ;
assign n5655 =  ( n5654 ) ? ( n5262 ) : ( dptr_hi ) ;
assign n5656 =  ( n5652 ) ? ( n5256 ) : ( n5655 ) ;
assign n5657 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5658 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n5659 =  ( n5658 ) & (wr )  ;
assign n5660 =  ( n5659 ) ? ( n5298 ) : ( dptr_hi ) ;
assign n5661 =  ( n5657 ) ? ( bv_8_0_n69 ) : ( n5660 ) ;
assign n5662 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5663 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n5664 =  ( n5663 ) & (wr )  ;
assign n5665 =  ( n5664 ) ? ( n5378 ) : ( dptr_hi ) ;
assign n5666 =  ( n5662 ) ? ( n5372 ) : ( n5665 ) ;
assign n5667 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5668 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n5669 =  ( n5668 ) & (wr )  ;
assign n5670 =  ( n5669 ) ? ( n4782 ) : ( dptr_lo ) ;
assign n5671 =  ( n5667 ) ? ( n4782 ) : ( n5670 ) ;
assign n5672 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5673 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n5674 =  ( n5673 ) & (wr )  ;
assign n5675 =  ( n5674 ) ? ( n4841 ) : ( dptr_lo ) ;
assign n5676 =  ( n5672 ) ? ( n4841 ) : ( n5675 ) ;
assign n5677 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5678 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n5679 =  ( n5678 ) & (wr )  ;
assign n5680 =  ( n5679 ) ? ( n4867 ) : ( dptr_lo ) ;
assign n5681 =  ( n5677 ) ? ( n4867 ) : ( n5680 ) ;
assign n5682 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5683 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n5684 =  ( n5683 ) & (wr )  ;
assign n5685 =  ( n5684 ) ? ( n4937 ) : ( dptr_lo ) ;
assign n5686 =  ( n5682 ) ? ( n4937 ) : ( n5685 ) ;
assign n5687 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5688 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n5689 =  ( n5688 ) & (wr )  ;
assign n5690 =  ( n5689 ) ? ( n4948 ) : ( dptr_lo ) ;
assign n5691 =  ( n5687 ) ? ( n4948 ) : ( n5690 ) ;
assign n5692 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5693 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n5694 =  ( n5693 ) & (wr )  ;
assign n5695 =  ( n5694 ) ? ( n4959 ) : ( dptr_lo ) ;
assign n5696 =  ( n5692 ) ? ( n4959 ) : ( n5695 ) ;
assign n5697 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5698 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n5699 =  ( n5698 ) & (wr )  ;
assign n5700 =  ( n5699 ) ? ( n5035 ) : ( dptr_lo ) ;
assign n5701 =  ( n5697 ) ? ( n5035 ) : ( n5700 ) ;
assign n5702 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5703 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n5704 =  ( n5703 ) & (wr )  ;
assign n5705 =  ( n5704 ) ? ( n5071 ) : ( dptr_lo ) ;
assign n5706 =  ( n5702 ) ? ( n5071 ) : ( n5705 ) ;
assign n5707 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5708 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n5709 =  ( n5708 ) & (wr )  ;
assign n5710 =  ( n5709 ) ? ( n5099 ) : ( dptr_lo ) ;
assign n5711 =  ( n5707 ) ? ( n5099 ) : ( n5710 ) ;
assign n5712 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5713 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n5714 =  ( n5713 ) & (wr )  ;
assign n5715 =  ( n5714 ) ? ( n5140 ) : ( dptr_lo ) ;
assign n5716 =  ( n5712 ) ? ( n5140 ) : ( n5715 ) ;
assign n5717 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5718 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n5719 =  ( n5718 ) & (wr )  ;
assign n5720 =  ( n5719 ) ? ( n5168 ) : ( dptr_lo ) ;
assign n5721 =  ( n5717 ) ? ( n5168 ) : ( n5720 ) ;
assign n5722 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5723 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n5724 =  ( n5723 ) & (wr )  ;
assign n5725 =  ( n5724 ) ? ( n5206 ) : ( dptr_lo ) ;
assign n5726 =  ( n5722 ) ? ( n5206 ) : ( n5725 ) ;
assign n5727 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5728 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n5729 =  ( n5728 ) & (wr )  ;
assign n5730 =  ( n5729 ) ? ( n5262 ) : ( dptr_lo ) ;
assign n5731 =  ( n5727 ) ? ( n5262 ) : ( n5730 ) ;
assign n5732 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5733 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n5734 =  ( n5733 ) & (wr )  ;
assign n5735 =  ( n5734 ) ? ( n5298 ) : ( dptr_lo ) ;
assign n5736 =  ( n5732 ) ? ( n5298 ) : ( n5735 ) ;
assign n5737 =  ( wr_sfr ) == ( bv_2_3_n3495 )  ;
assign n5738 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n5739 =  ( n5738 ) & (wr )  ;
assign n5740 =  ( n5739 ) ? ( n5378 ) : ( dptr_lo ) ;
assign n5741 =  ( n5737 ) ? ( n5378 ) : ( n5740 ) ;
assign n5742 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n5743 =  ( n5742 ) & (wr )  ;
assign n5744 =  ( n5743 ) ? ( n4782 ) : ( p0 ) ;
assign n5745 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n5746 =  ( n5745 ) & (wr )  ;
assign n5747 =  ( n5746 ) ? ( n4841 ) : ( p0 ) ;
assign n5748 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n5749 =  ( n5748 ) & (wr )  ;
assign n5750 =  ( n5749 ) ? ( n5449 ) : ( p0 ) ;
assign n5751 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n5752 =  ( n5751 ) & (wr )  ;
assign n5753 =  ( n5752 ) ? ( n4906 ) : ( p0 ) ;
assign n5754 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n5755 =  ( n5754 ) & (wr )  ;
assign n5756 =  ( n5755 ) ? ( n5485 ) : ( p0 ) ;
assign n5757 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n5758 =  ( n5757 ) & (wr )  ;
assign n5759 =  ( n5758 ) ? ( n5512 ) : ( p0 ) ;
assign n5760 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n5761 =  ( n5760 ) & (wr )  ;
assign n5762 =  ( n5761 ) ? ( bv_8_0_n69 ) : ( p0 ) ;
assign n5763 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n5764 =  ( n5763 ) & (wr )  ;
assign n5765 =  ( n5764 ) ? ( n5071 ) : ( p0 ) ;
assign n5766 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n5767 =  ( n5766 ) & (wr )  ;
assign n5768 =  ( n5767 ) ? ( n5096 ) : ( p0 ) ;
assign n5769 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n5770 =  ( n5769 ) & (wr )  ;
assign n5771 =  ( n5770 ) ? ( n5123 ) : ( p0 ) ;
assign n5772 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n5773 =  ( n5772 ) & (wr )  ;
assign n5774 =  ( n5773 ) ? ( n5165 ) : ( p0 ) ;
assign n5775 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n5776 =  ( n5775 ) & (wr )  ;
assign n5777 =  ( n5776 ) ? ( n5204 ) : ( p0 ) ;
assign n5778 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n5779 =  ( n5778 ) & (wr )  ;
assign n5780 =  ( n5779 ) ? ( n5262 ) : ( p0 ) ;
assign n5781 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n5782 =  ( n5781 ) & (wr )  ;
assign n5783 =  ( n5782 ) ? ( n5298 ) : ( p0 ) ;
assign n5784 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n5785 =  ( n5784 ) & (wr )  ;
assign n5786 =  ( n5785 ) ? ( n5325 ) : ( p0 ) ;
assign n5787 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n5788 =  ( n5787 ) & (wr )  ;
assign n5789 =  ( n5788 ) ? ( n4782 ) : ( p1 ) ;
assign n5790 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n5791 =  ( n5790 ) & (wr )  ;
assign n5792 =  ( n5791 ) ? ( n4841 ) : ( p1 ) ;
assign n5793 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n5794 =  ( n5793 ) & (wr )  ;
assign n5795 =  ( n5794 ) ? ( n5449 ) : ( p1 ) ;
assign n5796 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n5797 =  ( n5796 ) & (wr )  ;
assign n5798 =  ( n5797 ) ? ( n4906 ) : ( p1 ) ;
assign n5799 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n5800 =  ( n5799 ) & (wr )  ;
assign n5801 =  ( n5800 ) ? ( n5485 ) : ( p1 ) ;
assign n5802 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n5803 =  ( n5802 ) & (wr )  ;
assign n5804 =  ( n5803 ) ? ( n5512 ) : ( p1 ) ;
assign n5805 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n5806 =  ( n5805 ) & (wr )  ;
assign n5807 =  ( n5806 ) ? ( bv_8_0_n69 ) : ( p1 ) ;
assign n5808 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n5809 =  ( n5808 ) & (wr )  ;
assign n5810 =  ( n5809 ) ? ( n5071 ) : ( p1 ) ;
assign n5811 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n5812 =  ( n5811 ) & (wr )  ;
assign n5813 =  ( n5812 ) ? ( n5096 ) : ( p1 ) ;
assign n5814 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n5815 =  ( n5814 ) & (wr )  ;
assign n5816 =  ( n5815 ) ? ( n5123 ) : ( p1 ) ;
assign n5817 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n5818 =  ( n5817 ) & (wr )  ;
assign n5819 =  ( n5818 ) ? ( n5165 ) : ( p1 ) ;
assign n5820 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n5821 =  ( n5820 ) & (wr )  ;
assign n5822 =  ( n5821 ) ? ( n5204 ) : ( p1 ) ;
assign n5823 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n5824 =  ( n5823 ) & (wr )  ;
assign n5825 =  ( n5824 ) ? ( n5262 ) : ( p1 ) ;
assign n5826 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n5827 =  ( n5826 ) & (wr )  ;
assign n5828 =  ( n5827 ) ? ( n5298 ) : ( p1 ) ;
assign n5829 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n5830 =  ( n5829 ) & (wr )  ;
assign n5831 =  ( n5830 ) ? ( n5325 ) : ( p1 ) ;
assign n5832 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n5833 =  ( n5832 ) & (wr )  ;
assign n5834 =  ( n5833 ) ? ( n4782 ) : ( p2 ) ;
assign n5835 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n5836 =  ( n5835 ) & (wr )  ;
assign n5837 =  ( n5836 ) ? ( n4841 ) : ( p2 ) ;
assign n5838 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n5839 =  ( n5838 ) & (wr )  ;
assign n5840 =  ( n5839 ) ? ( n5449 ) : ( p2 ) ;
assign n5841 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n5842 =  ( n5841 ) & (wr )  ;
assign n5843 =  ( n5842 ) ? ( n4906 ) : ( p2 ) ;
assign n5844 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n5845 =  ( n5844 ) & (wr )  ;
assign n5846 =  ( n5845 ) ? ( n5485 ) : ( p2 ) ;
assign n5847 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n5848 =  ( n5847 ) & (wr )  ;
assign n5849 =  ( n5848 ) ? ( n5512 ) : ( p2 ) ;
assign n5850 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n5851 =  ( n5850 ) & (wr )  ;
assign n5852 =  ( n5851 ) ? ( bv_8_0_n69 ) : ( p2 ) ;
assign n5853 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n5854 =  ( n5853 ) & (wr )  ;
assign n5855 =  ( n5854 ) ? ( n5071 ) : ( p2 ) ;
assign n5856 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n5857 =  ( n5856 ) & (wr )  ;
assign n5858 =  ( n5857 ) ? ( n5096 ) : ( p2 ) ;
assign n5859 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n5860 =  ( n5859 ) & (wr )  ;
assign n5861 =  ( n5860 ) ? ( n5123 ) : ( p2 ) ;
assign n5862 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n5863 =  ( n5862 ) & (wr )  ;
assign n5864 =  ( n5863 ) ? ( n5165 ) : ( p2 ) ;
assign n5865 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n5866 =  ( n5865 ) & (wr )  ;
assign n5867 =  ( n5866 ) ? ( n5204 ) : ( p2 ) ;
assign n5868 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n5869 =  ( n5868 ) & (wr )  ;
assign n5870 =  ( n5869 ) ? ( n5262 ) : ( p2 ) ;
assign n5871 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n5872 =  ( n5871 ) & (wr )  ;
assign n5873 =  ( n5872 ) ? ( n5298 ) : ( p2 ) ;
assign n5874 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n5875 =  ( n5874 ) & (wr )  ;
assign n5876 =  ( n5875 ) ? ( n5325 ) : ( p2 ) ;
assign n5877 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n5878 =  ( n5877 ) & (wr )  ;
assign n5879 =  ( n5878 ) ? ( n4782 ) : ( p3 ) ;
assign n5880 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n5881 =  ( n5880 ) & (wr )  ;
assign n5882 =  ( n5881 ) ? ( n4841 ) : ( p3 ) ;
assign n5883 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n5884 =  ( n5883 ) & (wr )  ;
assign n5885 =  ( n5884 ) ? ( n5449 ) : ( p3 ) ;
assign n5886 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n5887 =  ( n5886 ) & (wr )  ;
assign n5888 =  ( n5887 ) ? ( n4906 ) : ( p3 ) ;
assign n5889 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n5890 =  ( n5889 ) & (wr )  ;
assign n5891 =  ( n5890 ) ? ( n5485 ) : ( p3 ) ;
assign n5892 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n5893 =  ( n5892 ) & (wr )  ;
assign n5894 =  ( n5893 ) ? ( n5512 ) : ( p3 ) ;
assign n5895 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n5896 =  ( n5895 ) & (wr )  ;
assign n5897 =  ( n5896 ) ? ( bv_8_0_n69 ) : ( p3 ) ;
assign n5898 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n5899 =  ( n5898 ) & (wr )  ;
assign n5900 =  ( n5899 ) ? ( n5071 ) : ( p3 ) ;
assign n5901 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n5902 =  ( n5901 ) & (wr )  ;
assign n5903 =  ( n5902 ) ? ( n5096 ) : ( p3 ) ;
assign n5904 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n5905 =  ( n5904 ) & (wr )  ;
assign n5906 =  ( n5905 ) ? ( n5123 ) : ( p3 ) ;
assign n5907 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n5908 =  ( n5907 ) & (wr )  ;
assign n5909 =  ( n5908 ) ? ( n5165 ) : ( p3 ) ;
assign n5910 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n5911 =  ( n5910 ) & (wr )  ;
assign n5912 =  ( n5911 ) ? ( n5204 ) : ( p3 ) ;
assign n5913 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n5914 =  ( n5913 ) & (wr )  ;
assign n5915 =  ( n5914 ) ? ( n5262 ) : ( p3 ) ;
assign n5916 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n5917 =  ( n5916 ) & (wr )  ;
assign n5918 =  ( n5917 ) ? ( n5298 ) : ( p3 ) ;
assign n5919 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n5920 =  ( n5919 ) & (wr )  ;
assign n5921 =  ( n5920 ) ? ( n5325 ) : ( p3 ) ;
assign n5922 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n5923 =  ( n5922 ) & (wr )  ;
assign n5924 =  ( n5923 ) ? ( n4782 ) : ( tcon ) ;
assign n5925 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n5926 =  ( n5925 ) & (wr )  ;
assign n5927 =  ( n5926 ) ? ( n4841 ) : ( tcon ) ;
assign n5928 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n5929 =  ( n5928 ) & (wr )  ;
assign n5930 =  ( n5929 ) ? ( n4867 ) : ( tcon ) ;
assign n5931 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n5932 =  ( n5931 ) & (wr )  ;
assign n5933 =  ( n5932 ) ? ( n4937 ) : ( tcon ) ;
assign n5934 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n5935 =  ( n5934 ) & (wr )  ;
assign n5936 =  ( n5935 ) ? ( n4948 ) : ( tcon ) ;
assign n5937 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n5938 =  ( n5937 ) & (wr )  ;
assign n5939 =  ( n5938 ) ? ( n4959 ) : ( tcon ) ;
assign n5940 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n5941 =  ( n5940 ) & (wr )  ;
assign n5942 =  ( n5941 ) ? ( n5035 ) : ( tcon ) ;
assign n5943 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n5944 =  ( n5943 ) & (wr )  ;
assign n5945 =  ( n5944 ) ? ( n5071 ) : ( tcon ) ;
assign n5946 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n5947 =  ( n5946 ) & (wr )  ;
assign n5948 =  ( n5947 ) ? ( n5099 ) : ( tcon ) ;
assign n5949 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n5950 =  ( n5949 ) & (wr )  ;
assign n5951 =  ( n5950 ) ? ( n5140 ) : ( tcon ) ;
assign n5952 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n5953 =  ( n5952 ) & (wr )  ;
assign n5954 =  ( n5953 ) ? ( n5168 ) : ( tcon ) ;
assign n5955 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n5956 =  ( n5955 ) & (wr )  ;
assign n5957 =  ( n5956 ) ? ( n5206 ) : ( tcon ) ;
assign n5958 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n5959 =  ( n5958 ) & (wr )  ;
assign n5960 =  ( n5959 ) ? ( n5262 ) : ( tcon ) ;
assign n5961 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n5962 =  ( n5961 ) & (wr )  ;
assign n5963 =  ( n5962 ) ? ( n5298 ) : ( tcon ) ;
assign n5964 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n5965 =  ( n5964 ) & (wr )  ;
assign n5966 =  ( n5965 ) ? ( n5378 ) : ( tcon ) ;
assign n5967 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n5968 =  ( n5967 ) & (wr )  ;
assign n5969 =  ( n5968 ) ? ( n4782 ) : ( scon ) ;
assign n5970 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n5971 =  ( n5970 ) & (wr )  ;
assign n5972 =  ( n5971 ) ? ( n4841 ) : ( scon ) ;
assign n5973 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n5974 =  ( n5973 ) & (wr )  ;
assign n5975 =  ( n5974 ) ? ( n4867 ) : ( scon ) ;
assign n5976 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n5977 =  ( n5976 ) & (wr )  ;
assign n5978 =  ( n5977 ) ? ( n4937 ) : ( scon ) ;
assign n5979 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n5980 =  ( n5979 ) & (wr )  ;
assign n5981 =  ( n5980 ) ? ( n4948 ) : ( scon ) ;
assign n5982 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n5983 =  ( n5982 ) & (wr )  ;
assign n5984 =  ( n5983 ) ? ( n4959 ) : ( scon ) ;
assign n5985 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n5986 =  ( n5985 ) & (wr )  ;
assign n5987 =  ( n5986 ) ? ( n5035 ) : ( scon ) ;
assign n5988 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n5989 =  ( n5988 ) & (wr )  ;
assign n5990 =  ( n5989 ) ? ( n5071 ) : ( scon ) ;
assign n5991 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n5992 =  ( n5991 ) & (wr )  ;
assign n5993 =  ( n5992 ) ? ( n5099 ) : ( scon ) ;
assign n5994 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n5995 =  ( n5994 ) & (wr )  ;
assign n5996 =  ( n5995 ) ? ( n5140 ) : ( scon ) ;
assign n5997 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n5998 =  ( n5997 ) & (wr )  ;
assign n5999 =  ( n5998 ) ? ( n5168 ) : ( scon ) ;
assign n6000 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n6001 =  ( n6000 ) & (wr )  ;
assign n6002 =  ( n6001 ) ? ( n5206 ) : ( scon ) ;
assign n6003 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n6004 =  ( n6003 ) & (wr )  ;
assign n6005 =  ( n6004 ) ? ( n5262 ) : ( scon ) ;
assign n6006 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n6007 =  ( n6006 ) & (wr )  ;
assign n6008 =  ( n6007 ) ? ( n5298 ) : ( scon ) ;
assign n6009 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n6010 =  ( n6009 ) & (wr )  ;
assign n6011 =  ( n6010 ) ? ( n5378 ) : ( scon ) ;
assign n6012 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n6013 =  ( n6012 ) & (wr )  ;
assign n6014 =  ( n6013 ) ? ( n4782 ) : ( pcon ) ;
assign n6015 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n6016 =  ( n6015 ) & (wr )  ;
assign n6017 =  ( n6016 ) ? ( n4841 ) : ( pcon ) ;
assign n6018 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n6019 =  ( n6018 ) & (wr )  ;
assign n6020 =  ( n6019 ) ? ( n4867 ) : ( pcon ) ;
assign n6021 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n6022 =  ( n6021 ) & (wr )  ;
assign n6023 =  ( n6022 ) ? ( n4937 ) : ( pcon ) ;
assign n6024 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n6025 =  ( n6024 ) & (wr )  ;
assign n6026 =  ( n6025 ) ? ( n4948 ) : ( pcon ) ;
assign n6027 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n6028 =  ( n6027 ) & (wr )  ;
assign n6029 =  ( n6028 ) ? ( n4959 ) : ( pcon ) ;
assign n6030 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n6031 =  ( n6030 ) & (wr )  ;
assign n6032 =  ( n6031 ) ? ( n5035 ) : ( pcon ) ;
assign n6033 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n6034 =  ( n6033 ) & (wr )  ;
assign n6035 =  ( n6034 ) ? ( n5071 ) : ( pcon ) ;
assign n6036 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n6037 =  ( n6036 ) & (wr )  ;
assign n6038 =  ( n6037 ) ? ( n5099 ) : ( pcon ) ;
assign n6039 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n6040 =  ( n6039 ) & (wr )  ;
assign n6041 =  ( n6040 ) ? ( n5140 ) : ( pcon ) ;
assign n6042 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n6043 =  ( n6042 ) & (wr )  ;
assign n6044 =  ( n6043 ) ? ( n5168 ) : ( pcon ) ;
assign n6045 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n6046 =  ( n6045 ) & (wr )  ;
assign n6047 =  ( n6046 ) ? ( n5206 ) : ( pcon ) ;
assign n6048 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n6049 =  ( n6048 ) & (wr )  ;
assign n6050 =  ( n6049 ) ? ( n5262 ) : ( pcon ) ;
assign n6051 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n6052 =  ( n6051 ) & (wr )  ;
assign n6053 =  ( n6052 ) ? ( n5298 ) : ( pcon ) ;
assign n6054 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n6055 =  ( n6054 ) & (wr )  ;
assign n6056 =  ( n6055 ) ? ( n5378 ) : ( pcon ) ;
assign n6057 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n6058 =  ( n6057 ) & (wr )  ;
assign n6059 =  ( n6058 ) ? ( n4782 ) : ( sbuf ) ;
assign n6060 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n6061 =  ( n6060 ) & (wr )  ;
assign n6062 =  ( n6061 ) ? ( n4841 ) : ( sbuf ) ;
assign n6063 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n6064 =  ( n6063 ) & (wr )  ;
assign n6065 =  ( n6064 ) ? ( n4867 ) : ( sbuf ) ;
assign n6066 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n6067 =  ( n6066 ) & (wr )  ;
assign n6068 =  ( n6067 ) ? ( n4937 ) : ( sbuf ) ;
assign n6069 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n6070 =  ( n6069 ) & (wr )  ;
assign n6071 =  ( n6070 ) ? ( n4948 ) : ( sbuf ) ;
assign n6072 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n6073 =  ( n6072 ) & (wr )  ;
assign n6074 =  ( n6073 ) ? ( n4959 ) : ( sbuf ) ;
assign n6075 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n6076 =  ( n6075 ) & (wr )  ;
assign n6077 =  ( n6076 ) ? ( n5035 ) : ( sbuf ) ;
assign n6078 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n6079 =  ( n6078 ) & (wr )  ;
assign n6080 =  ( n6079 ) ? ( n5071 ) : ( sbuf ) ;
assign n6081 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n6082 =  ( n6081 ) & (wr )  ;
assign n6083 =  ( n6082 ) ? ( n5099 ) : ( sbuf ) ;
assign n6084 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n6085 =  ( n6084 ) & (wr )  ;
assign n6086 =  ( n6085 ) ? ( n5140 ) : ( sbuf ) ;
assign n6087 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n6088 =  ( n6087 ) & (wr )  ;
assign n6089 =  ( n6088 ) ? ( n5168 ) : ( sbuf ) ;
assign n6090 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n6091 =  ( n6090 ) & (wr )  ;
assign n6092 =  ( n6091 ) ? ( n5206 ) : ( sbuf ) ;
assign n6093 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n6094 =  ( n6093 ) & (wr )  ;
assign n6095 =  ( n6094 ) ? ( n5262 ) : ( sbuf ) ;
assign n6096 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n6097 =  ( n6096 ) & (wr )  ;
assign n6098 =  ( n6097 ) ? ( n5298 ) : ( sbuf ) ;
assign n6099 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n6100 =  ( n6099 ) & (wr )  ;
assign n6101 =  ( n6100 ) ? ( n5378 ) : ( sbuf ) ;
assign n6102 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n6103 =  ( n6102 ) & (wr )  ;
assign n6104 =  ( n6103 ) ? ( n4782 ) : ( th0 ) ;
assign n6105 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n6106 =  ( n6105 ) & (wr )  ;
assign n6107 =  ( n6106 ) ? ( n4841 ) : ( th0 ) ;
assign n6108 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n6109 =  ( n6108 ) & (wr )  ;
assign n6110 =  ( n6109 ) ? ( n4867 ) : ( th0 ) ;
assign n6111 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n6112 =  ( n6111 ) & (wr )  ;
assign n6113 =  ( n6112 ) ? ( n4937 ) : ( th0 ) ;
assign n6114 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n6115 =  ( n6114 ) & (wr )  ;
assign n6116 =  ( n6115 ) ? ( n4948 ) : ( th0 ) ;
assign n6117 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n6118 =  ( n6117 ) & (wr )  ;
assign n6119 =  ( n6118 ) ? ( n4959 ) : ( th0 ) ;
assign n6120 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n6121 =  ( n6120 ) & (wr )  ;
assign n6122 =  ( n6121 ) ? ( n5035 ) : ( th0 ) ;
assign n6123 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n6124 =  ( n6123 ) & (wr )  ;
assign n6125 =  ( n6124 ) ? ( n5071 ) : ( th0 ) ;
assign n6126 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n6127 =  ( n6126 ) & (wr )  ;
assign n6128 =  ( n6127 ) ? ( n5099 ) : ( th0 ) ;
assign n6129 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n6130 =  ( n6129 ) & (wr )  ;
assign n6131 =  ( n6130 ) ? ( n5140 ) : ( th0 ) ;
assign n6132 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n6133 =  ( n6132 ) & (wr )  ;
assign n6134 =  ( n6133 ) ? ( n5168 ) : ( th0 ) ;
assign n6135 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n6136 =  ( n6135 ) & (wr )  ;
assign n6137 =  ( n6136 ) ? ( n5206 ) : ( th0 ) ;
assign n6138 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n6139 =  ( n6138 ) & (wr )  ;
assign n6140 =  ( n6139 ) ? ( n5262 ) : ( th0 ) ;
assign n6141 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n6142 =  ( n6141 ) & (wr )  ;
assign n6143 =  ( n6142 ) ? ( n5298 ) : ( th0 ) ;
assign n6144 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n6145 =  ( n6144 ) & (wr )  ;
assign n6146 =  ( n6145 ) ? ( n5378 ) : ( th0 ) ;
assign n6147 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n6148 =  ( n6147 ) & (wr )  ;
assign n6149 =  ( n6148 ) ? ( n4782 ) : ( th1 ) ;
assign n6150 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n6151 =  ( n6150 ) & (wr )  ;
assign n6152 =  ( n6151 ) ? ( n4841 ) : ( th1 ) ;
assign n6153 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n6154 =  ( n6153 ) & (wr )  ;
assign n6155 =  ( n6154 ) ? ( n4867 ) : ( th1 ) ;
assign n6156 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n6157 =  ( n6156 ) & (wr )  ;
assign n6158 =  ( n6157 ) ? ( n4937 ) : ( th1 ) ;
assign n6159 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n6160 =  ( n6159 ) & (wr )  ;
assign n6161 =  ( n6160 ) ? ( n4948 ) : ( th1 ) ;
assign n6162 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n6163 =  ( n6162 ) & (wr )  ;
assign n6164 =  ( n6163 ) ? ( n4959 ) : ( th1 ) ;
assign n6165 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n6166 =  ( n6165 ) & (wr )  ;
assign n6167 =  ( n6166 ) ? ( n5035 ) : ( th1 ) ;
assign n6168 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n6169 =  ( n6168 ) & (wr )  ;
assign n6170 =  ( n6169 ) ? ( n5071 ) : ( th1 ) ;
assign n6171 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n6172 =  ( n6171 ) & (wr )  ;
assign n6173 =  ( n6172 ) ? ( n5099 ) : ( th1 ) ;
assign n6174 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n6175 =  ( n6174 ) & (wr )  ;
assign n6176 =  ( n6175 ) ? ( n5140 ) : ( th1 ) ;
assign n6177 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n6178 =  ( n6177 ) & (wr )  ;
assign n6179 =  ( n6178 ) ? ( n5168 ) : ( th1 ) ;
assign n6180 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n6181 =  ( n6180 ) & (wr )  ;
assign n6182 =  ( n6181 ) ? ( n5206 ) : ( th1 ) ;
assign n6183 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n6184 =  ( n6183 ) & (wr )  ;
assign n6185 =  ( n6184 ) ? ( n5262 ) : ( th1 ) ;
assign n6186 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n6187 =  ( n6186 ) & (wr )  ;
assign n6188 =  ( n6187 ) ? ( n5298 ) : ( th1 ) ;
assign n6189 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n6190 =  ( n6189 ) & (wr )  ;
assign n6191 =  ( n6190 ) ? ( n5378 ) : ( th1 ) ;
assign n6192 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n6193 =  ( n6192 ) & (wr )  ;
assign n6194 =  ( n6193 ) ? ( n4782 ) : ( tl0 ) ;
assign n6195 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n6196 =  ( n6195 ) & (wr )  ;
assign n6197 =  ( n6196 ) ? ( n4841 ) : ( tl0 ) ;
assign n6198 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n6199 =  ( n6198 ) & (wr )  ;
assign n6200 =  ( n6199 ) ? ( n4867 ) : ( tl0 ) ;
assign n6201 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n6202 =  ( n6201 ) & (wr )  ;
assign n6203 =  ( n6202 ) ? ( n4937 ) : ( tl0 ) ;
assign n6204 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n6205 =  ( n6204 ) & (wr )  ;
assign n6206 =  ( n6205 ) ? ( n4948 ) : ( tl0 ) ;
assign n6207 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n6208 =  ( n6207 ) & (wr )  ;
assign n6209 =  ( n6208 ) ? ( n4959 ) : ( tl0 ) ;
assign n6210 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n6211 =  ( n6210 ) & (wr )  ;
assign n6212 =  ( n6211 ) ? ( n5035 ) : ( tl0 ) ;
assign n6213 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n6214 =  ( n6213 ) & (wr )  ;
assign n6215 =  ( n6214 ) ? ( n5071 ) : ( tl0 ) ;
assign n6216 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n6217 =  ( n6216 ) & (wr )  ;
assign n6218 =  ( n6217 ) ? ( n5099 ) : ( tl0 ) ;
assign n6219 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n6220 =  ( n6219 ) & (wr )  ;
assign n6221 =  ( n6220 ) ? ( n5140 ) : ( tl0 ) ;
assign n6222 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n6223 =  ( n6222 ) & (wr )  ;
assign n6224 =  ( n6223 ) ? ( n5168 ) : ( tl0 ) ;
assign n6225 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n6226 =  ( n6225 ) & (wr )  ;
assign n6227 =  ( n6226 ) ? ( n5206 ) : ( tl0 ) ;
assign n6228 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n6229 =  ( n6228 ) & (wr )  ;
assign n6230 =  ( n6229 ) ? ( n5262 ) : ( tl0 ) ;
assign n6231 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n6232 =  ( n6231 ) & (wr )  ;
assign n6233 =  ( n6232 ) ? ( n5298 ) : ( tl0 ) ;
assign n6234 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n6235 =  ( n6234 ) & (wr )  ;
assign n6236 =  ( n6235 ) ? ( n5378 ) : ( tl0 ) ;
assign n6237 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n6238 =  ( n6237 ) & (wr )  ;
assign n6239 =  ( n6238 ) ? ( n4782 ) : ( tl1 ) ;
assign n6240 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n6241 =  ( n6240 ) & (wr )  ;
assign n6242 =  ( n6241 ) ? ( n4841 ) : ( tl1 ) ;
assign n6243 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n6244 =  ( n6243 ) & (wr )  ;
assign n6245 =  ( n6244 ) ? ( n4867 ) : ( tl1 ) ;
assign n6246 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n6247 =  ( n6246 ) & (wr )  ;
assign n6248 =  ( n6247 ) ? ( n4937 ) : ( tl1 ) ;
assign n6249 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n6250 =  ( n6249 ) & (wr )  ;
assign n6251 =  ( n6250 ) ? ( n4948 ) : ( tl1 ) ;
assign n6252 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n6253 =  ( n6252 ) & (wr )  ;
assign n6254 =  ( n6253 ) ? ( n4959 ) : ( tl1 ) ;
assign n6255 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n6256 =  ( n6255 ) & (wr )  ;
assign n6257 =  ( n6256 ) ? ( n5035 ) : ( tl1 ) ;
assign n6258 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n6259 =  ( n6258 ) & (wr )  ;
assign n6260 =  ( n6259 ) ? ( n5071 ) : ( tl1 ) ;
assign n6261 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n6262 =  ( n6261 ) & (wr )  ;
assign n6263 =  ( n6262 ) ? ( n5099 ) : ( tl1 ) ;
assign n6264 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n6265 =  ( n6264 ) & (wr )  ;
assign n6266 =  ( n6265 ) ? ( n5140 ) : ( tl1 ) ;
assign n6267 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n6268 =  ( n6267 ) & (wr )  ;
assign n6269 =  ( n6268 ) ? ( n5168 ) : ( tl1 ) ;
assign n6270 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n6271 =  ( n6270 ) & (wr )  ;
assign n6272 =  ( n6271 ) ? ( n5206 ) : ( tl1 ) ;
assign n6273 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n6274 =  ( n6273 ) & (wr )  ;
assign n6275 =  ( n6274 ) ? ( n5262 ) : ( tl1 ) ;
assign n6276 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n6277 =  ( n6276 ) & (wr )  ;
assign n6278 =  ( n6277 ) ? ( n5298 ) : ( tl1 ) ;
assign n6279 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n6280 =  ( n6279 ) & (wr )  ;
assign n6281 =  ( n6280 ) ? ( n5378 ) : ( tl1 ) ;
assign n6282 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n6283 =  ( n6282 ) & (wr )  ;
assign n6284 =  ( n6283 ) ? ( n4782 ) : ( tmod ) ;
assign n6285 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n6286 =  ( n6285 ) & (wr )  ;
assign n6287 =  ( n6286 ) ? ( n4841 ) : ( tmod ) ;
assign n6288 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n6289 =  ( n6288 ) & (wr )  ;
assign n6290 =  ( n6289 ) ? ( n4867 ) : ( tmod ) ;
assign n6291 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n6292 =  ( n6291 ) & (wr )  ;
assign n6293 =  ( n6292 ) ? ( n4937 ) : ( tmod ) ;
assign n6294 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n6295 =  ( n6294 ) & (wr )  ;
assign n6296 =  ( n6295 ) ? ( n4948 ) : ( tmod ) ;
assign n6297 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n6298 =  ( n6297 ) & (wr )  ;
assign n6299 =  ( n6298 ) ? ( n4959 ) : ( tmod ) ;
assign n6300 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n6301 =  ( n6300 ) & (wr )  ;
assign n6302 =  ( n6301 ) ? ( n5035 ) : ( tmod ) ;
assign n6303 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n6304 =  ( n6303 ) & (wr )  ;
assign n6305 =  ( n6304 ) ? ( n5071 ) : ( tmod ) ;
assign n6306 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n6307 =  ( n6306 ) & (wr )  ;
assign n6308 =  ( n6307 ) ? ( n5099 ) : ( tmod ) ;
assign n6309 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n6310 =  ( n6309 ) & (wr )  ;
assign n6311 =  ( n6310 ) ? ( n5140 ) : ( tmod ) ;
assign n6312 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n6313 =  ( n6312 ) & (wr )  ;
assign n6314 =  ( n6313 ) ? ( n5168 ) : ( tmod ) ;
assign n6315 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n6316 =  ( n6315 ) & (wr )  ;
assign n6317 =  ( n6316 ) ? ( n5206 ) : ( tmod ) ;
assign n6318 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n6319 =  ( n6318 ) & (wr )  ;
assign n6320 =  ( n6319 ) ? ( n5262 ) : ( tmod ) ;
assign n6321 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n6322 =  ( n6321 ) & (wr )  ;
assign n6323 =  ( n6322 ) ? ( n5298 ) : ( tmod ) ;
assign n6324 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n6325 =  ( n6324 ) & (wr )  ;
assign n6326 =  ( n6325 ) ? ( n5378 ) : ( tmod ) ;
assign n6327 = wr_addr[7:7] ;
assign n6328 =  ( n6327 ) == ( bv_1_0_n53 )  ;
assign n6329 =  ( wr_addr ) == ( bv_8_0_n69 )  ;
assign n6330 =  ( n6328 ) & (n6329 )  ;
assign n6331 =  ( n6330 ) & (wr )  ;
assign n6332 =  ( n6331 ) ? ( n4782 ) : ( iram_0 ) ;
assign n6333 = wr_addr[7:7] ;
assign n6334 =  ( n6333 ) == ( bv_1_0_n53 )  ;
assign n6335 =  ( wr_addr ) == ( bv_8_0_n69 )  ;
assign n6336 =  ( n6334 ) & (n6335 )  ;
assign n6337 =  ( n6336 ) & (wr )  ;
assign n6338 =  ( n6337 ) ? ( n4841 ) : ( iram_0 ) ;
assign n6339 = wr_addr[7:7] ;
assign n6340 =  ( n6339 ) == ( bv_1_0_n53 )  ;
assign n6341 =  ( wr_addr ) == ( bv_8_0_n69 )  ;
assign n6342 =  ( n6340 ) & (n6341 )  ;
assign n6343 =  ( n6342 ) & (wr )  ;
assign n6344 =  ( n6343 ) ? ( n5449 ) : ( iram_0 ) ;
assign n6345 = wr_addr[7:7] ;
assign n6346 =  ( n6345 ) == ( bv_1_0_n53 )  ;
assign n6347 =  ( wr_addr ) == ( bv_8_0_n69 )  ;
assign n6348 =  ( n6346 ) & (n6347 )  ;
assign n6349 =  ( n6348 ) & (wr )  ;
assign n6350 =  ( n6349 ) ? ( n4906 ) : ( iram_0 ) ;
assign n6351 = wr_addr[7:7] ;
assign n6352 =  ( n6351 ) == ( bv_1_0_n53 )  ;
assign n6353 =  ( wr_addr ) == ( bv_8_0_n69 )  ;
assign n6354 =  ( n6352 ) & (n6353 )  ;
assign n6355 =  ( n6354 ) & (wr )  ;
assign n6356 =  ( n6355 ) ? ( n5485 ) : ( iram_0 ) ;
assign n6357 = wr_addr[7:7] ;
assign n6358 =  ( n6357 ) == ( bv_1_0_n53 )  ;
assign n6359 =  ( wr_addr ) == ( bv_8_0_n69 )  ;
assign n6360 =  ( n6358 ) & (n6359 )  ;
assign n6361 =  ( n6360 ) & (wr )  ;
assign n6362 =  ( n6361 ) ? ( n5512 ) : ( iram_0 ) ;
assign n6363 = wr_addr[7:7] ;
assign n6364 =  ( n6363 ) == ( bv_1_0_n53 )  ;
assign n6365 =  ( wr_addr ) == ( bv_8_0_n69 )  ;
assign n6366 =  ( n6364 ) & (n6365 )  ;
assign n6367 =  ( n6366 ) & (wr )  ;
assign n6368 =  ( n6367 ) ? ( bv_8_0_n69 ) : ( iram_0 ) ;
assign n6369 = wr_addr[7:7] ;
assign n6370 =  ( n6369 ) == ( bv_1_0_n53 )  ;
assign n6371 =  ( wr_addr ) == ( bv_8_0_n69 )  ;
assign n6372 =  ( n6370 ) & (n6371 )  ;
assign n6373 =  ( n6372 ) & (wr )  ;
assign n6374 =  ( n6373 ) ? ( n5071 ) : ( iram_0 ) ;
assign n6375 = wr_addr[7:7] ;
assign n6376 =  ( n6375 ) == ( bv_1_0_n53 )  ;
assign n6377 =  ( wr_addr ) == ( bv_8_0_n69 )  ;
assign n6378 =  ( n6376 ) & (n6377 )  ;
assign n6379 =  ( n6378 ) & (wr )  ;
assign n6380 =  ( n6379 ) ? ( n5096 ) : ( iram_0 ) ;
assign n6381 = wr_addr[7:7] ;
assign n6382 =  ( n6381 ) == ( bv_1_0_n53 )  ;
assign n6383 =  ( wr_addr ) == ( bv_8_0_n69 )  ;
assign n6384 =  ( n6382 ) & (n6383 )  ;
assign n6385 =  ( n6384 ) & (wr )  ;
assign n6386 =  ( n6385 ) ? ( n5123 ) : ( iram_0 ) ;
assign n6387 = wr_addr[7:7] ;
assign n6388 =  ( n6387 ) == ( bv_1_0_n53 )  ;
assign n6389 =  ( wr_addr ) == ( bv_8_0_n69 )  ;
assign n6390 =  ( n6388 ) & (n6389 )  ;
assign n6391 =  ( n6390 ) & (wr )  ;
assign n6392 =  ( n6391 ) ? ( n5165 ) : ( iram_0 ) ;
assign n6393 = wr_addr[7:7] ;
assign n6394 =  ( n6393 ) == ( bv_1_0_n53 )  ;
assign n6395 =  ( wr_addr ) == ( bv_8_0_n69 )  ;
assign n6396 =  ( n6394 ) & (n6395 )  ;
assign n6397 =  ( n6396 ) & (wr )  ;
assign n6398 =  ( n6397 ) ? ( n5204 ) : ( iram_0 ) ;
assign n6399 = wr_addr[7:7] ;
assign n6400 =  ( n6399 ) == ( bv_1_0_n53 )  ;
assign n6401 =  ( wr_addr ) == ( bv_8_0_n69 )  ;
assign n6402 =  ( n6400 ) & (n6401 )  ;
assign n6403 =  ( n6402 ) & (wr )  ;
assign n6404 =  ( n6403 ) ? ( n5262 ) : ( iram_0 ) ;
assign n6405 = wr_addr[7:7] ;
assign n6406 =  ( n6405 ) == ( bv_1_0_n53 )  ;
assign n6407 =  ( wr_addr ) == ( bv_8_0_n69 )  ;
assign n6408 =  ( n6406 ) & (n6407 )  ;
assign n6409 =  ( n6408 ) & (wr )  ;
assign n6410 =  ( n6409 ) ? ( n5298 ) : ( iram_0 ) ;
assign n6411 = wr_addr[7:7] ;
assign n6412 =  ( n6411 ) == ( bv_1_0_n53 )  ;
assign n6413 =  ( wr_addr ) == ( bv_8_0_n69 )  ;
assign n6414 =  ( n6412 ) & (n6413 )  ;
assign n6415 =  ( n6414 ) & (wr )  ;
assign n6416 =  ( n6415 ) ? ( n5325 ) : ( iram_0 ) ;
assign n6417 = wr_addr[7:7] ;
assign n6418 =  ( n6417 ) == ( bv_1_0_n53 )  ;
assign n6419 =  ( wr_addr ) == ( bv_8_1_n71 )  ;
assign n6420 =  ( n6418 ) & (n6419 )  ;
assign n6421 =  ( n6420 ) & (wr )  ;
assign n6422 =  ( n6421 ) ? ( n4782 ) : ( iram_1 ) ;
assign n6423 = wr_addr[7:7] ;
assign n6424 =  ( n6423 ) == ( bv_1_0_n53 )  ;
assign n6425 =  ( wr_addr ) == ( bv_8_1_n71 )  ;
assign n6426 =  ( n6424 ) & (n6425 )  ;
assign n6427 =  ( n6426 ) & (wr )  ;
assign n6428 =  ( n6427 ) ? ( n4841 ) : ( iram_1 ) ;
assign n6429 = wr_addr[7:7] ;
assign n6430 =  ( n6429 ) == ( bv_1_0_n53 )  ;
assign n6431 =  ( wr_addr ) == ( bv_8_1_n71 )  ;
assign n6432 =  ( n6430 ) & (n6431 )  ;
assign n6433 =  ( n6432 ) & (wr )  ;
assign n6434 =  ( n6433 ) ? ( n5449 ) : ( iram_1 ) ;
assign n6435 = wr_addr[7:7] ;
assign n6436 =  ( n6435 ) == ( bv_1_0_n53 )  ;
assign n6437 =  ( wr_addr ) == ( bv_8_1_n71 )  ;
assign n6438 =  ( n6436 ) & (n6437 )  ;
assign n6439 =  ( n6438 ) & (wr )  ;
assign n6440 =  ( n6439 ) ? ( n4906 ) : ( iram_1 ) ;
assign n6441 = wr_addr[7:7] ;
assign n6442 =  ( n6441 ) == ( bv_1_0_n53 )  ;
assign n6443 =  ( wr_addr ) == ( bv_8_1_n71 )  ;
assign n6444 =  ( n6442 ) & (n6443 )  ;
assign n6445 =  ( n6444 ) & (wr )  ;
assign n6446 =  ( n6445 ) ? ( n5485 ) : ( iram_1 ) ;
assign n6447 = wr_addr[7:7] ;
assign n6448 =  ( n6447 ) == ( bv_1_0_n53 )  ;
assign n6449 =  ( wr_addr ) == ( bv_8_1_n71 )  ;
assign n6450 =  ( n6448 ) & (n6449 )  ;
assign n6451 =  ( n6450 ) & (wr )  ;
assign n6452 =  ( n6451 ) ? ( n5512 ) : ( iram_1 ) ;
assign n6453 = wr_addr[7:7] ;
assign n6454 =  ( n6453 ) == ( bv_1_0_n53 )  ;
assign n6455 =  ( wr_addr ) == ( bv_8_1_n71 )  ;
assign n6456 =  ( n6454 ) & (n6455 )  ;
assign n6457 =  ( n6456 ) & (wr )  ;
assign n6458 =  ( n6457 ) ? ( bv_8_0_n69 ) : ( iram_1 ) ;
assign n6459 = wr_addr[7:7] ;
assign n6460 =  ( n6459 ) == ( bv_1_0_n53 )  ;
assign n6461 =  ( wr_addr ) == ( bv_8_1_n71 )  ;
assign n6462 =  ( n6460 ) & (n6461 )  ;
assign n6463 =  ( n6462 ) & (wr )  ;
assign n6464 =  ( n6463 ) ? ( n5071 ) : ( iram_1 ) ;
assign n6465 = wr_addr[7:7] ;
assign n6466 =  ( n6465 ) == ( bv_1_0_n53 )  ;
assign n6467 =  ( wr_addr ) == ( bv_8_1_n71 )  ;
assign n6468 =  ( n6466 ) & (n6467 )  ;
assign n6469 =  ( n6468 ) & (wr )  ;
assign n6470 =  ( n6469 ) ? ( n5096 ) : ( iram_1 ) ;
assign n6471 = wr_addr[7:7] ;
assign n6472 =  ( n6471 ) == ( bv_1_0_n53 )  ;
assign n6473 =  ( wr_addr ) == ( bv_8_1_n71 )  ;
assign n6474 =  ( n6472 ) & (n6473 )  ;
assign n6475 =  ( n6474 ) & (wr )  ;
assign n6476 =  ( n6475 ) ? ( n5123 ) : ( iram_1 ) ;
assign n6477 = wr_addr[7:7] ;
assign n6478 =  ( n6477 ) == ( bv_1_0_n53 )  ;
assign n6479 =  ( wr_addr ) == ( bv_8_1_n71 )  ;
assign n6480 =  ( n6478 ) & (n6479 )  ;
assign n6481 =  ( n6480 ) & (wr )  ;
assign n6482 =  ( n6481 ) ? ( n5165 ) : ( iram_1 ) ;
assign n6483 = wr_addr[7:7] ;
assign n6484 =  ( n6483 ) == ( bv_1_0_n53 )  ;
assign n6485 =  ( wr_addr ) == ( bv_8_1_n71 )  ;
assign n6486 =  ( n6484 ) & (n6485 )  ;
assign n6487 =  ( n6486 ) & (wr )  ;
assign n6488 =  ( n6487 ) ? ( n5204 ) : ( iram_1 ) ;
assign n6489 = wr_addr[7:7] ;
assign n6490 =  ( n6489 ) == ( bv_1_0_n53 )  ;
assign n6491 =  ( wr_addr ) == ( bv_8_1_n71 )  ;
assign n6492 =  ( n6490 ) & (n6491 )  ;
assign n6493 =  ( n6492 ) & (wr )  ;
assign n6494 =  ( n6493 ) ? ( n5262 ) : ( iram_1 ) ;
assign n6495 = wr_addr[7:7] ;
assign n6496 =  ( n6495 ) == ( bv_1_0_n53 )  ;
assign n6497 =  ( wr_addr ) == ( bv_8_1_n71 )  ;
assign n6498 =  ( n6496 ) & (n6497 )  ;
assign n6499 =  ( n6498 ) & (wr )  ;
assign n6500 =  ( n6499 ) ? ( n5298 ) : ( iram_1 ) ;
assign n6501 = wr_addr[7:7] ;
assign n6502 =  ( n6501 ) == ( bv_1_0_n53 )  ;
assign n6503 =  ( wr_addr ) == ( bv_8_1_n71 )  ;
assign n6504 =  ( n6502 ) & (n6503 )  ;
assign n6505 =  ( n6504 ) & (wr )  ;
assign n6506 =  ( n6505 ) ? ( n5325 ) : ( iram_1 ) ;
assign n6507 = wr_addr[7:7] ;
assign n6508 =  ( n6507 ) == ( bv_1_0_n53 )  ;
assign n6509 =  ( wr_addr ) == ( bv_8_2_n73 )  ;
assign n6510 =  ( n6508 ) & (n6509 )  ;
assign n6511 =  ( n6510 ) & (wr )  ;
assign n6512 =  ( n6511 ) ? ( n4782 ) : ( iram_2 ) ;
assign n6513 = wr_addr[7:7] ;
assign n6514 =  ( n6513 ) == ( bv_1_0_n53 )  ;
assign n6515 =  ( wr_addr ) == ( bv_8_2_n73 )  ;
assign n6516 =  ( n6514 ) & (n6515 )  ;
assign n6517 =  ( n6516 ) & (wr )  ;
assign n6518 =  ( n6517 ) ? ( n4841 ) : ( iram_2 ) ;
assign n6519 = wr_addr[7:7] ;
assign n6520 =  ( n6519 ) == ( bv_1_0_n53 )  ;
assign n6521 =  ( wr_addr ) == ( bv_8_2_n73 )  ;
assign n6522 =  ( n6520 ) & (n6521 )  ;
assign n6523 =  ( n6522 ) & (wr )  ;
assign n6524 =  ( n6523 ) ? ( n5449 ) : ( iram_2 ) ;
assign n6525 = wr_addr[7:7] ;
assign n6526 =  ( n6525 ) == ( bv_1_0_n53 )  ;
assign n6527 =  ( wr_addr ) == ( bv_8_2_n73 )  ;
assign n6528 =  ( n6526 ) & (n6527 )  ;
assign n6529 =  ( n6528 ) & (wr )  ;
assign n6530 =  ( n6529 ) ? ( n4906 ) : ( iram_2 ) ;
assign n6531 = wr_addr[7:7] ;
assign n6532 =  ( n6531 ) == ( bv_1_0_n53 )  ;
assign n6533 =  ( wr_addr ) == ( bv_8_2_n73 )  ;
assign n6534 =  ( n6532 ) & (n6533 )  ;
assign n6535 =  ( n6534 ) & (wr )  ;
assign n6536 =  ( n6535 ) ? ( n5485 ) : ( iram_2 ) ;
assign n6537 = wr_addr[7:7] ;
assign n6538 =  ( n6537 ) == ( bv_1_0_n53 )  ;
assign n6539 =  ( wr_addr ) == ( bv_8_2_n73 )  ;
assign n6540 =  ( n6538 ) & (n6539 )  ;
assign n6541 =  ( n6540 ) & (wr )  ;
assign n6542 =  ( n6541 ) ? ( n5512 ) : ( iram_2 ) ;
assign n6543 = wr_addr[7:7] ;
assign n6544 =  ( n6543 ) == ( bv_1_0_n53 )  ;
assign n6545 =  ( wr_addr ) == ( bv_8_2_n73 )  ;
assign n6546 =  ( n6544 ) & (n6545 )  ;
assign n6547 =  ( n6546 ) & (wr )  ;
assign n6548 =  ( n6547 ) ? ( bv_8_0_n69 ) : ( iram_2 ) ;
assign n6549 = wr_addr[7:7] ;
assign n6550 =  ( n6549 ) == ( bv_1_0_n53 )  ;
assign n6551 =  ( wr_addr ) == ( bv_8_2_n73 )  ;
assign n6552 =  ( n6550 ) & (n6551 )  ;
assign n6553 =  ( n6552 ) & (wr )  ;
assign n6554 =  ( n6553 ) ? ( n5071 ) : ( iram_2 ) ;
assign n6555 = wr_addr[7:7] ;
assign n6556 =  ( n6555 ) == ( bv_1_0_n53 )  ;
assign n6557 =  ( wr_addr ) == ( bv_8_2_n73 )  ;
assign n6558 =  ( n6556 ) & (n6557 )  ;
assign n6559 =  ( n6558 ) & (wr )  ;
assign n6560 =  ( n6559 ) ? ( n5096 ) : ( iram_2 ) ;
assign n6561 = wr_addr[7:7] ;
assign n6562 =  ( n6561 ) == ( bv_1_0_n53 )  ;
assign n6563 =  ( wr_addr ) == ( bv_8_2_n73 )  ;
assign n6564 =  ( n6562 ) & (n6563 )  ;
assign n6565 =  ( n6564 ) & (wr )  ;
assign n6566 =  ( n6565 ) ? ( n5123 ) : ( iram_2 ) ;
assign n6567 = wr_addr[7:7] ;
assign n6568 =  ( n6567 ) == ( bv_1_0_n53 )  ;
assign n6569 =  ( wr_addr ) == ( bv_8_2_n73 )  ;
assign n6570 =  ( n6568 ) & (n6569 )  ;
assign n6571 =  ( n6570 ) & (wr )  ;
assign n6572 =  ( n6571 ) ? ( n5165 ) : ( iram_2 ) ;
assign n6573 = wr_addr[7:7] ;
assign n6574 =  ( n6573 ) == ( bv_1_0_n53 )  ;
assign n6575 =  ( wr_addr ) == ( bv_8_2_n73 )  ;
assign n6576 =  ( n6574 ) & (n6575 )  ;
assign n6577 =  ( n6576 ) & (wr )  ;
assign n6578 =  ( n6577 ) ? ( n5204 ) : ( iram_2 ) ;
assign n6579 = wr_addr[7:7] ;
assign n6580 =  ( n6579 ) == ( bv_1_0_n53 )  ;
assign n6581 =  ( wr_addr ) == ( bv_8_2_n73 )  ;
assign n6582 =  ( n6580 ) & (n6581 )  ;
assign n6583 =  ( n6582 ) & (wr )  ;
assign n6584 =  ( n6583 ) ? ( n5262 ) : ( iram_2 ) ;
assign n6585 = wr_addr[7:7] ;
assign n6586 =  ( n6585 ) == ( bv_1_0_n53 )  ;
assign n6587 =  ( wr_addr ) == ( bv_8_2_n73 )  ;
assign n6588 =  ( n6586 ) & (n6587 )  ;
assign n6589 =  ( n6588 ) & (wr )  ;
assign n6590 =  ( n6589 ) ? ( n5298 ) : ( iram_2 ) ;
assign n6591 = wr_addr[7:7] ;
assign n6592 =  ( n6591 ) == ( bv_1_0_n53 )  ;
assign n6593 =  ( wr_addr ) == ( bv_8_2_n73 )  ;
assign n6594 =  ( n6592 ) & (n6593 )  ;
assign n6595 =  ( n6594 ) & (wr )  ;
assign n6596 =  ( n6595 ) ? ( n5325 ) : ( iram_2 ) ;
assign n6597 = wr_addr[7:7] ;
assign n6598 =  ( n6597 ) == ( bv_1_0_n53 )  ;
assign n6599 =  ( wr_addr ) == ( bv_8_3_n75 )  ;
assign n6600 =  ( n6598 ) & (n6599 )  ;
assign n6601 =  ( n6600 ) & (wr )  ;
assign n6602 =  ( n6601 ) ? ( n4782 ) : ( iram_3 ) ;
assign n6603 = wr_addr[7:7] ;
assign n6604 =  ( n6603 ) == ( bv_1_0_n53 )  ;
assign n6605 =  ( wr_addr ) == ( bv_8_3_n75 )  ;
assign n6606 =  ( n6604 ) & (n6605 )  ;
assign n6607 =  ( n6606 ) & (wr )  ;
assign n6608 =  ( n6607 ) ? ( n4841 ) : ( iram_3 ) ;
assign n6609 = wr_addr[7:7] ;
assign n6610 =  ( n6609 ) == ( bv_1_0_n53 )  ;
assign n6611 =  ( wr_addr ) == ( bv_8_3_n75 )  ;
assign n6612 =  ( n6610 ) & (n6611 )  ;
assign n6613 =  ( n6612 ) & (wr )  ;
assign n6614 =  ( n6613 ) ? ( n5449 ) : ( iram_3 ) ;
assign n6615 = wr_addr[7:7] ;
assign n6616 =  ( n6615 ) == ( bv_1_0_n53 )  ;
assign n6617 =  ( wr_addr ) == ( bv_8_3_n75 )  ;
assign n6618 =  ( n6616 ) & (n6617 )  ;
assign n6619 =  ( n6618 ) & (wr )  ;
assign n6620 =  ( n6619 ) ? ( n4906 ) : ( iram_3 ) ;
assign n6621 = wr_addr[7:7] ;
assign n6622 =  ( n6621 ) == ( bv_1_0_n53 )  ;
assign n6623 =  ( wr_addr ) == ( bv_8_3_n75 )  ;
assign n6624 =  ( n6622 ) & (n6623 )  ;
assign n6625 =  ( n6624 ) & (wr )  ;
assign n6626 =  ( n6625 ) ? ( n5485 ) : ( iram_3 ) ;
assign n6627 = wr_addr[7:7] ;
assign n6628 =  ( n6627 ) == ( bv_1_0_n53 )  ;
assign n6629 =  ( wr_addr ) == ( bv_8_3_n75 )  ;
assign n6630 =  ( n6628 ) & (n6629 )  ;
assign n6631 =  ( n6630 ) & (wr )  ;
assign n6632 =  ( n6631 ) ? ( n5512 ) : ( iram_3 ) ;
assign n6633 = wr_addr[7:7] ;
assign n6634 =  ( n6633 ) == ( bv_1_0_n53 )  ;
assign n6635 =  ( wr_addr ) == ( bv_8_3_n75 )  ;
assign n6636 =  ( n6634 ) & (n6635 )  ;
assign n6637 =  ( n6636 ) & (wr )  ;
assign n6638 =  ( n6637 ) ? ( bv_8_0_n69 ) : ( iram_3 ) ;
assign n6639 = wr_addr[7:7] ;
assign n6640 =  ( n6639 ) == ( bv_1_0_n53 )  ;
assign n6641 =  ( wr_addr ) == ( bv_8_3_n75 )  ;
assign n6642 =  ( n6640 ) & (n6641 )  ;
assign n6643 =  ( n6642 ) & (wr )  ;
assign n6644 =  ( n6643 ) ? ( n5071 ) : ( iram_3 ) ;
assign n6645 = wr_addr[7:7] ;
assign n6646 =  ( n6645 ) == ( bv_1_0_n53 )  ;
assign n6647 =  ( wr_addr ) == ( bv_8_3_n75 )  ;
assign n6648 =  ( n6646 ) & (n6647 )  ;
assign n6649 =  ( n6648 ) & (wr )  ;
assign n6650 =  ( n6649 ) ? ( n5096 ) : ( iram_3 ) ;
assign n6651 = wr_addr[7:7] ;
assign n6652 =  ( n6651 ) == ( bv_1_0_n53 )  ;
assign n6653 =  ( wr_addr ) == ( bv_8_3_n75 )  ;
assign n6654 =  ( n6652 ) & (n6653 )  ;
assign n6655 =  ( n6654 ) & (wr )  ;
assign n6656 =  ( n6655 ) ? ( n5123 ) : ( iram_3 ) ;
assign n6657 = wr_addr[7:7] ;
assign n6658 =  ( n6657 ) == ( bv_1_0_n53 )  ;
assign n6659 =  ( wr_addr ) == ( bv_8_3_n75 )  ;
assign n6660 =  ( n6658 ) & (n6659 )  ;
assign n6661 =  ( n6660 ) & (wr )  ;
assign n6662 =  ( n6661 ) ? ( n5165 ) : ( iram_3 ) ;
assign n6663 = wr_addr[7:7] ;
assign n6664 =  ( n6663 ) == ( bv_1_0_n53 )  ;
assign n6665 =  ( wr_addr ) == ( bv_8_3_n75 )  ;
assign n6666 =  ( n6664 ) & (n6665 )  ;
assign n6667 =  ( n6666 ) & (wr )  ;
assign n6668 =  ( n6667 ) ? ( n5204 ) : ( iram_3 ) ;
assign n6669 = wr_addr[7:7] ;
assign n6670 =  ( n6669 ) == ( bv_1_0_n53 )  ;
assign n6671 =  ( wr_addr ) == ( bv_8_3_n75 )  ;
assign n6672 =  ( n6670 ) & (n6671 )  ;
assign n6673 =  ( n6672 ) & (wr )  ;
assign n6674 =  ( n6673 ) ? ( n5262 ) : ( iram_3 ) ;
assign n6675 = wr_addr[7:7] ;
assign n6676 =  ( n6675 ) == ( bv_1_0_n53 )  ;
assign n6677 =  ( wr_addr ) == ( bv_8_3_n75 )  ;
assign n6678 =  ( n6676 ) & (n6677 )  ;
assign n6679 =  ( n6678 ) & (wr )  ;
assign n6680 =  ( n6679 ) ? ( n5298 ) : ( iram_3 ) ;
assign n6681 = wr_addr[7:7] ;
assign n6682 =  ( n6681 ) == ( bv_1_0_n53 )  ;
assign n6683 =  ( wr_addr ) == ( bv_8_3_n75 )  ;
assign n6684 =  ( n6682 ) & (n6683 )  ;
assign n6685 =  ( n6684 ) & (wr )  ;
assign n6686 =  ( n6685 ) ? ( n5325 ) : ( iram_3 ) ;
assign n6687 = wr_addr[7:7] ;
assign n6688 =  ( n6687 ) == ( bv_1_0_n53 )  ;
assign n6689 =  ( wr_addr ) == ( bv_8_4_n77 )  ;
assign n6690 =  ( n6688 ) & (n6689 )  ;
assign n6691 =  ( n6690 ) & (wr )  ;
assign n6692 =  ( n6691 ) ? ( n4782 ) : ( iram_4 ) ;
assign n6693 = wr_addr[7:7] ;
assign n6694 =  ( n6693 ) == ( bv_1_0_n53 )  ;
assign n6695 =  ( wr_addr ) == ( bv_8_4_n77 )  ;
assign n6696 =  ( n6694 ) & (n6695 )  ;
assign n6697 =  ( n6696 ) & (wr )  ;
assign n6698 =  ( n6697 ) ? ( n4841 ) : ( iram_4 ) ;
assign n6699 = wr_addr[7:7] ;
assign n6700 =  ( n6699 ) == ( bv_1_0_n53 )  ;
assign n6701 =  ( wr_addr ) == ( bv_8_4_n77 )  ;
assign n6702 =  ( n6700 ) & (n6701 )  ;
assign n6703 =  ( n6702 ) & (wr )  ;
assign n6704 =  ( n6703 ) ? ( n5449 ) : ( iram_4 ) ;
assign n6705 = wr_addr[7:7] ;
assign n6706 =  ( n6705 ) == ( bv_1_0_n53 )  ;
assign n6707 =  ( wr_addr ) == ( bv_8_4_n77 )  ;
assign n6708 =  ( n6706 ) & (n6707 )  ;
assign n6709 =  ( n6708 ) & (wr )  ;
assign n6710 =  ( n6709 ) ? ( n4906 ) : ( iram_4 ) ;
assign n6711 = wr_addr[7:7] ;
assign n6712 =  ( n6711 ) == ( bv_1_0_n53 )  ;
assign n6713 =  ( wr_addr ) == ( bv_8_4_n77 )  ;
assign n6714 =  ( n6712 ) & (n6713 )  ;
assign n6715 =  ( n6714 ) & (wr )  ;
assign n6716 =  ( n6715 ) ? ( n5485 ) : ( iram_4 ) ;
assign n6717 = wr_addr[7:7] ;
assign n6718 =  ( n6717 ) == ( bv_1_0_n53 )  ;
assign n6719 =  ( wr_addr ) == ( bv_8_4_n77 )  ;
assign n6720 =  ( n6718 ) & (n6719 )  ;
assign n6721 =  ( n6720 ) & (wr )  ;
assign n6722 =  ( n6721 ) ? ( n5512 ) : ( iram_4 ) ;
assign n6723 = wr_addr[7:7] ;
assign n6724 =  ( n6723 ) == ( bv_1_0_n53 )  ;
assign n6725 =  ( wr_addr ) == ( bv_8_4_n77 )  ;
assign n6726 =  ( n6724 ) & (n6725 )  ;
assign n6727 =  ( n6726 ) & (wr )  ;
assign n6728 =  ( n6727 ) ? ( bv_8_0_n69 ) : ( iram_4 ) ;
assign n6729 = wr_addr[7:7] ;
assign n6730 =  ( n6729 ) == ( bv_1_0_n53 )  ;
assign n6731 =  ( wr_addr ) == ( bv_8_4_n77 )  ;
assign n6732 =  ( n6730 ) & (n6731 )  ;
assign n6733 =  ( n6732 ) & (wr )  ;
assign n6734 =  ( n6733 ) ? ( n5071 ) : ( iram_4 ) ;
assign n6735 = wr_addr[7:7] ;
assign n6736 =  ( n6735 ) == ( bv_1_0_n53 )  ;
assign n6737 =  ( wr_addr ) == ( bv_8_4_n77 )  ;
assign n6738 =  ( n6736 ) & (n6737 )  ;
assign n6739 =  ( n6738 ) & (wr )  ;
assign n6740 =  ( n6739 ) ? ( n5096 ) : ( iram_4 ) ;
assign n6741 = wr_addr[7:7] ;
assign n6742 =  ( n6741 ) == ( bv_1_0_n53 )  ;
assign n6743 =  ( wr_addr ) == ( bv_8_4_n77 )  ;
assign n6744 =  ( n6742 ) & (n6743 )  ;
assign n6745 =  ( n6744 ) & (wr )  ;
assign n6746 =  ( n6745 ) ? ( n5123 ) : ( iram_4 ) ;
assign n6747 = wr_addr[7:7] ;
assign n6748 =  ( n6747 ) == ( bv_1_0_n53 )  ;
assign n6749 =  ( wr_addr ) == ( bv_8_4_n77 )  ;
assign n6750 =  ( n6748 ) & (n6749 )  ;
assign n6751 =  ( n6750 ) & (wr )  ;
assign n6752 =  ( n6751 ) ? ( n5165 ) : ( iram_4 ) ;
assign n6753 = wr_addr[7:7] ;
assign n6754 =  ( n6753 ) == ( bv_1_0_n53 )  ;
assign n6755 =  ( wr_addr ) == ( bv_8_4_n77 )  ;
assign n6756 =  ( n6754 ) & (n6755 )  ;
assign n6757 =  ( n6756 ) & (wr )  ;
assign n6758 =  ( n6757 ) ? ( n5204 ) : ( iram_4 ) ;
assign n6759 = wr_addr[7:7] ;
assign n6760 =  ( n6759 ) == ( bv_1_0_n53 )  ;
assign n6761 =  ( wr_addr ) == ( bv_8_4_n77 )  ;
assign n6762 =  ( n6760 ) & (n6761 )  ;
assign n6763 =  ( n6762 ) & (wr )  ;
assign n6764 =  ( n6763 ) ? ( n5262 ) : ( iram_4 ) ;
assign n6765 = wr_addr[7:7] ;
assign n6766 =  ( n6765 ) == ( bv_1_0_n53 )  ;
assign n6767 =  ( wr_addr ) == ( bv_8_4_n77 )  ;
assign n6768 =  ( n6766 ) & (n6767 )  ;
assign n6769 =  ( n6768 ) & (wr )  ;
assign n6770 =  ( n6769 ) ? ( n5298 ) : ( iram_4 ) ;
assign n6771 = wr_addr[7:7] ;
assign n6772 =  ( n6771 ) == ( bv_1_0_n53 )  ;
assign n6773 =  ( wr_addr ) == ( bv_8_4_n77 )  ;
assign n6774 =  ( n6772 ) & (n6773 )  ;
assign n6775 =  ( n6774 ) & (wr )  ;
assign n6776 =  ( n6775 ) ? ( n5325 ) : ( iram_4 ) ;
assign n6777 = wr_addr[7:7] ;
assign n6778 =  ( n6777 ) == ( bv_1_0_n53 )  ;
assign n6779 =  ( wr_addr ) == ( bv_8_5_n79 )  ;
assign n6780 =  ( n6778 ) & (n6779 )  ;
assign n6781 =  ( n6780 ) & (wr )  ;
assign n6782 =  ( n6781 ) ? ( n4782 ) : ( iram_5 ) ;
assign n6783 = wr_addr[7:7] ;
assign n6784 =  ( n6783 ) == ( bv_1_0_n53 )  ;
assign n6785 =  ( wr_addr ) == ( bv_8_5_n79 )  ;
assign n6786 =  ( n6784 ) & (n6785 )  ;
assign n6787 =  ( n6786 ) & (wr )  ;
assign n6788 =  ( n6787 ) ? ( n4841 ) : ( iram_5 ) ;
assign n6789 = wr_addr[7:7] ;
assign n6790 =  ( n6789 ) == ( bv_1_0_n53 )  ;
assign n6791 =  ( wr_addr ) == ( bv_8_5_n79 )  ;
assign n6792 =  ( n6790 ) & (n6791 )  ;
assign n6793 =  ( n6792 ) & (wr )  ;
assign n6794 =  ( n6793 ) ? ( n5449 ) : ( iram_5 ) ;
assign n6795 = wr_addr[7:7] ;
assign n6796 =  ( n6795 ) == ( bv_1_0_n53 )  ;
assign n6797 =  ( wr_addr ) == ( bv_8_5_n79 )  ;
assign n6798 =  ( n6796 ) & (n6797 )  ;
assign n6799 =  ( n6798 ) & (wr )  ;
assign n6800 =  ( n6799 ) ? ( n4906 ) : ( iram_5 ) ;
assign n6801 = wr_addr[7:7] ;
assign n6802 =  ( n6801 ) == ( bv_1_0_n53 )  ;
assign n6803 =  ( wr_addr ) == ( bv_8_5_n79 )  ;
assign n6804 =  ( n6802 ) & (n6803 )  ;
assign n6805 =  ( n6804 ) & (wr )  ;
assign n6806 =  ( n6805 ) ? ( n5485 ) : ( iram_5 ) ;
assign n6807 = wr_addr[7:7] ;
assign n6808 =  ( n6807 ) == ( bv_1_0_n53 )  ;
assign n6809 =  ( wr_addr ) == ( bv_8_5_n79 )  ;
assign n6810 =  ( n6808 ) & (n6809 )  ;
assign n6811 =  ( n6810 ) & (wr )  ;
assign n6812 =  ( n6811 ) ? ( n5512 ) : ( iram_5 ) ;
assign n6813 = wr_addr[7:7] ;
assign n6814 =  ( n6813 ) == ( bv_1_0_n53 )  ;
assign n6815 =  ( wr_addr ) == ( bv_8_5_n79 )  ;
assign n6816 =  ( n6814 ) & (n6815 )  ;
assign n6817 =  ( n6816 ) & (wr )  ;
assign n6818 =  ( n6817 ) ? ( bv_8_0_n69 ) : ( iram_5 ) ;
assign n6819 = wr_addr[7:7] ;
assign n6820 =  ( n6819 ) == ( bv_1_0_n53 )  ;
assign n6821 =  ( wr_addr ) == ( bv_8_5_n79 )  ;
assign n6822 =  ( n6820 ) & (n6821 )  ;
assign n6823 =  ( n6822 ) & (wr )  ;
assign n6824 =  ( n6823 ) ? ( n5071 ) : ( iram_5 ) ;
assign n6825 = wr_addr[7:7] ;
assign n6826 =  ( n6825 ) == ( bv_1_0_n53 )  ;
assign n6827 =  ( wr_addr ) == ( bv_8_5_n79 )  ;
assign n6828 =  ( n6826 ) & (n6827 )  ;
assign n6829 =  ( n6828 ) & (wr )  ;
assign n6830 =  ( n6829 ) ? ( n5096 ) : ( iram_5 ) ;
assign n6831 = wr_addr[7:7] ;
assign n6832 =  ( n6831 ) == ( bv_1_0_n53 )  ;
assign n6833 =  ( wr_addr ) == ( bv_8_5_n79 )  ;
assign n6834 =  ( n6832 ) & (n6833 )  ;
assign n6835 =  ( n6834 ) & (wr )  ;
assign n6836 =  ( n6835 ) ? ( n5123 ) : ( iram_5 ) ;
assign n6837 = wr_addr[7:7] ;
assign n6838 =  ( n6837 ) == ( bv_1_0_n53 )  ;
assign n6839 =  ( wr_addr ) == ( bv_8_5_n79 )  ;
assign n6840 =  ( n6838 ) & (n6839 )  ;
assign n6841 =  ( n6840 ) & (wr )  ;
assign n6842 =  ( n6841 ) ? ( n5165 ) : ( iram_5 ) ;
assign n6843 = wr_addr[7:7] ;
assign n6844 =  ( n6843 ) == ( bv_1_0_n53 )  ;
assign n6845 =  ( wr_addr ) == ( bv_8_5_n79 )  ;
assign n6846 =  ( n6844 ) & (n6845 )  ;
assign n6847 =  ( n6846 ) & (wr )  ;
assign n6848 =  ( n6847 ) ? ( n5204 ) : ( iram_5 ) ;
assign n6849 = wr_addr[7:7] ;
assign n6850 =  ( n6849 ) == ( bv_1_0_n53 )  ;
assign n6851 =  ( wr_addr ) == ( bv_8_5_n79 )  ;
assign n6852 =  ( n6850 ) & (n6851 )  ;
assign n6853 =  ( n6852 ) & (wr )  ;
assign n6854 =  ( n6853 ) ? ( n5262 ) : ( iram_5 ) ;
assign n6855 = wr_addr[7:7] ;
assign n6856 =  ( n6855 ) == ( bv_1_0_n53 )  ;
assign n6857 =  ( wr_addr ) == ( bv_8_5_n79 )  ;
assign n6858 =  ( n6856 ) & (n6857 )  ;
assign n6859 =  ( n6858 ) & (wr )  ;
assign n6860 =  ( n6859 ) ? ( n5298 ) : ( iram_5 ) ;
assign n6861 = wr_addr[7:7] ;
assign n6862 =  ( n6861 ) == ( bv_1_0_n53 )  ;
assign n6863 =  ( wr_addr ) == ( bv_8_5_n79 )  ;
assign n6864 =  ( n6862 ) & (n6863 )  ;
assign n6865 =  ( n6864 ) & (wr )  ;
assign n6866 =  ( n6865 ) ? ( n5325 ) : ( iram_5 ) ;
assign n6867 = wr_addr[7:7] ;
assign n6868 =  ( n6867 ) == ( bv_1_0_n53 )  ;
assign n6869 =  ( wr_addr ) == ( bv_8_6_n81 )  ;
assign n6870 =  ( n6868 ) & (n6869 )  ;
assign n6871 =  ( n6870 ) & (wr )  ;
assign n6872 =  ( n6871 ) ? ( n4782 ) : ( iram_6 ) ;
assign n6873 = wr_addr[7:7] ;
assign n6874 =  ( n6873 ) == ( bv_1_0_n53 )  ;
assign n6875 =  ( wr_addr ) == ( bv_8_6_n81 )  ;
assign n6876 =  ( n6874 ) & (n6875 )  ;
assign n6877 =  ( n6876 ) & (wr )  ;
assign n6878 =  ( n6877 ) ? ( n4841 ) : ( iram_6 ) ;
assign n6879 = wr_addr[7:7] ;
assign n6880 =  ( n6879 ) == ( bv_1_0_n53 )  ;
assign n6881 =  ( wr_addr ) == ( bv_8_6_n81 )  ;
assign n6882 =  ( n6880 ) & (n6881 )  ;
assign n6883 =  ( n6882 ) & (wr )  ;
assign n6884 =  ( n6883 ) ? ( n5449 ) : ( iram_6 ) ;
assign n6885 = wr_addr[7:7] ;
assign n6886 =  ( n6885 ) == ( bv_1_0_n53 )  ;
assign n6887 =  ( wr_addr ) == ( bv_8_6_n81 )  ;
assign n6888 =  ( n6886 ) & (n6887 )  ;
assign n6889 =  ( n6888 ) & (wr )  ;
assign n6890 =  ( n6889 ) ? ( n4906 ) : ( iram_6 ) ;
assign n6891 = wr_addr[7:7] ;
assign n6892 =  ( n6891 ) == ( bv_1_0_n53 )  ;
assign n6893 =  ( wr_addr ) == ( bv_8_6_n81 )  ;
assign n6894 =  ( n6892 ) & (n6893 )  ;
assign n6895 =  ( n6894 ) & (wr )  ;
assign n6896 =  ( n6895 ) ? ( n5485 ) : ( iram_6 ) ;
assign n6897 = wr_addr[7:7] ;
assign n6898 =  ( n6897 ) == ( bv_1_0_n53 )  ;
assign n6899 =  ( wr_addr ) == ( bv_8_6_n81 )  ;
assign n6900 =  ( n6898 ) & (n6899 )  ;
assign n6901 =  ( n6900 ) & (wr )  ;
assign n6902 =  ( n6901 ) ? ( n5512 ) : ( iram_6 ) ;
assign n6903 = wr_addr[7:7] ;
assign n6904 =  ( n6903 ) == ( bv_1_0_n53 )  ;
assign n6905 =  ( wr_addr ) == ( bv_8_6_n81 )  ;
assign n6906 =  ( n6904 ) & (n6905 )  ;
assign n6907 =  ( n6906 ) & (wr )  ;
assign n6908 =  ( n6907 ) ? ( bv_8_0_n69 ) : ( iram_6 ) ;
assign n6909 = wr_addr[7:7] ;
assign n6910 =  ( n6909 ) == ( bv_1_0_n53 )  ;
assign n6911 =  ( wr_addr ) == ( bv_8_6_n81 )  ;
assign n6912 =  ( n6910 ) & (n6911 )  ;
assign n6913 =  ( n6912 ) & (wr )  ;
assign n6914 =  ( n6913 ) ? ( n5071 ) : ( iram_6 ) ;
assign n6915 = wr_addr[7:7] ;
assign n6916 =  ( n6915 ) == ( bv_1_0_n53 )  ;
assign n6917 =  ( wr_addr ) == ( bv_8_6_n81 )  ;
assign n6918 =  ( n6916 ) & (n6917 )  ;
assign n6919 =  ( n6918 ) & (wr )  ;
assign n6920 =  ( n6919 ) ? ( n5096 ) : ( iram_6 ) ;
assign n6921 = wr_addr[7:7] ;
assign n6922 =  ( n6921 ) == ( bv_1_0_n53 )  ;
assign n6923 =  ( wr_addr ) == ( bv_8_6_n81 )  ;
assign n6924 =  ( n6922 ) & (n6923 )  ;
assign n6925 =  ( n6924 ) & (wr )  ;
assign n6926 =  ( n6925 ) ? ( n5123 ) : ( iram_6 ) ;
assign n6927 = wr_addr[7:7] ;
assign n6928 =  ( n6927 ) == ( bv_1_0_n53 )  ;
assign n6929 =  ( wr_addr ) == ( bv_8_6_n81 )  ;
assign n6930 =  ( n6928 ) & (n6929 )  ;
assign n6931 =  ( n6930 ) & (wr )  ;
assign n6932 =  ( n6931 ) ? ( n5165 ) : ( iram_6 ) ;
assign n6933 = wr_addr[7:7] ;
assign n6934 =  ( n6933 ) == ( bv_1_0_n53 )  ;
assign n6935 =  ( wr_addr ) == ( bv_8_6_n81 )  ;
assign n6936 =  ( n6934 ) & (n6935 )  ;
assign n6937 =  ( n6936 ) & (wr )  ;
assign n6938 =  ( n6937 ) ? ( n5204 ) : ( iram_6 ) ;
assign n6939 = wr_addr[7:7] ;
assign n6940 =  ( n6939 ) == ( bv_1_0_n53 )  ;
assign n6941 =  ( wr_addr ) == ( bv_8_6_n81 )  ;
assign n6942 =  ( n6940 ) & (n6941 )  ;
assign n6943 =  ( n6942 ) & (wr )  ;
assign n6944 =  ( n6943 ) ? ( n5262 ) : ( iram_6 ) ;
assign n6945 = wr_addr[7:7] ;
assign n6946 =  ( n6945 ) == ( bv_1_0_n53 )  ;
assign n6947 =  ( wr_addr ) == ( bv_8_6_n81 )  ;
assign n6948 =  ( n6946 ) & (n6947 )  ;
assign n6949 =  ( n6948 ) & (wr )  ;
assign n6950 =  ( n6949 ) ? ( n5298 ) : ( iram_6 ) ;
assign n6951 = wr_addr[7:7] ;
assign n6952 =  ( n6951 ) == ( bv_1_0_n53 )  ;
assign n6953 =  ( wr_addr ) == ( bv_8_6_n81 )  ;
assign n6954 =  ( n6952 ) & (n6953 )  ;
assign n6955 =  ( n6954 ) & (wr )  ;
assign n6956 =  ( n6955 ) ? ( n5325 ) : ( iram_6 ) ;
assign n6957 = wr_addr[7:7] ;
assign n6958 =  ( n6957 ) == ( bv_1_0_n53 )  ;
assign n6959 =  ( wr_addr ) == ( bv_8_7_n83 )  ;
assign n6960 =  ( n6958 ) & (n6959 )  ;
assign n6961 =  ( n6960 ) & (wr )  ;
assign n6962 =  ( n6961 ) ? ( n4782 ) : ( iram_7 ) ;
assign n6963 = wr_addr[7:7] ;
assign n6964 =  ( n6963 ) == ( bv_1_0_n53 )  ;
assign n6965 =  ( wr_addr ) == ( bv_8_7_n83 )  ;
assign n6966 =  ( n6964 ) & (n6965 )  ;
assign n6967 =  ( n6966 ) & (wr )  ;
assign n6968 =  ( n6967 ) ? ( n4841 ) : ( iram_7 ) ;
assign n6969 = wr_addr[7:7] ;
assign n6970 =  ( n6969 ) == ( bv_1_0_n53 )  ;
assign n6971 =  ( wr_addr ) == ( bv_8_7_n83 )  ;
assign n6972 =  ( n6970 ) & (n6971 )  ;
assign n6973 =  ( n6972 ) & (wr )  ;
assign n6974 =  ( n6973 ) ? ( n5449 ) : ( iram_7 ) ;
assign n6975 = wr_addr[7:7] ;
assign n6976 =  ( n6975 ) == ( bv_1_0_n53 )  ;
assign n6977 =  ( wr_addr ) == ( bv_8_7_n83 )  ;
assign n6978 =  ( n6976 ) & (n6977 )  ;
assign n6979 =  ( n6978 ) & (wr )  ;
assign n6980 =  ( n6979 ) ? ( n4906 ) : ( iram_7 ) ;
assign n6981 = wr_addr[7:7] ;
assign n6982 =  ( n6981 ) == ( bv_1_0_n53 )  ;
assign n6983 =  ( wr_addr ) == ( bv_8_7_n83 )  ;
assign n6984 =  ( n6982 ) & (n6983 )  ;
assign n6985 =  ( n6984 ) & (wr )  ;
assign n6986 =  ( n6985 ) ? ( n5485 ) : ( iram_7 ) ;
assign n6987 = wr_addr[7:7] ;
assign n6988 =  ( n6987 ) == ( bv_1_0_n53 )  ;
assign n6989 =  ( wr_addr ) == ( bv_8_7_n83 )  ;
assign n6990 =  ( n6988 ) & (n6989 )  ;
assign n6991 =  ( n6990 ) & (wr )  ;
assign n6992 =  ( n6991 ) ? ( n5512 ) : ( iram_7 ) ;
assign n6993 = wr_addr[7:7] ;
assign n6994 =  ( n6993 ) == ( bv_1_0_n53 )  ;
assign n6995 =  ( wr_addr ) == ( bv_8_7_n83 )  ;
assign n6996 =  ( n6994 ) & (n6995 )  ;
assign n6997 =  ( n6996 ) & (wr )  ;
assign n6998 =  ( n6997 ) ? ( bv_8_0_n69 ) : ( iram_7 ) ;
assign n6999 = wr_addr[7:7] ;
assign n7000 =  ( n6999 ) == ( bv_1_0_n53 )  ;
assign n7001 =  ( wr_addr ) == ( bv_8_7_n83 )  ;
assign n7002 =  ( n7000 ) & (n7001 )  ;
assign n7003 =  ( n7002 ) & (wr )  ;
assign n7004 =  ( n7003 ) ? ( n5071 ) : ( iram_7 ) ;
assign n7005 = wr_addr[7:7] ;
assign n7006 =  ( n7005 ) == ( bv_1_0_n53 )  ;
assign n7007 =  ( wr_addr ) == ( bv_8_7_n83 )  ;
assign n7008 =  ( n7006 ) & (n7007 )  ;
assign n7009 =  ( n7008 ) & (wr )  ;
assign n7010 =  ( n7009 ) ? ( n5096 ) : ( iram_7 ) ;
assign n7011 = wr_addr[7:7] ;
assign n7012 =  ( n7011 ) == ( bv_1_0_n53 )  ;
assign n7013 =  ( wr_addr ) == ( bv_8_7_n83 )  ;
assign n7014 =  ( n7012 ) & (n7013 )  ;
assign n7015 =  ( n7014 ) & (wr )  ;
assign n7016 =  ( n7015 ) ? ( n5123 ) : ( iram_7 ) ;
assign n7017 = wr_addr[7:7] ;
assign n7018 =  ( n7017 ) == ( bv_1_0_n53 )  ;
assign n7019 =  ( wr_addr ) == ( bv_8_7_n83 )  ;
assign n7020 =  ( n7018 ) & (n7019 )  ;
assign n7021 =  ( n7020 ) & (wr )  ;
assign n7022 =  ( n7021 ) ? ( n5165 ) : ( iram_7 ) ;
assign n7023 = wr_addr[7:7] ;
assign n7024 =  ( n7023 ) == ( bv_1_0_n53 )  ;
assign n7025 =  ( wr_addr ) == ( bv_8_7_n83 )  ;
assign n7026 =  ( n7024 ) & (n7025 )  ;
assign n7027 =  ( n7026 ) & (wr )  ;
assign n7028 =  ( n7027 ) ? ( n5204 ) : ( iram_7 ) ;
assign n7029 = wr_addr[7:7] ;
assign n7030 =  ( n7029 ) == ( bv_1_0_n53 )  ;
assign n7031 =  ( wr_addr ) == ( bv_8_7_n83 )  ;
assign n7032 =  ( n7030 ) & (n7031 )  ;
assign n7033 =  ( n7032 ) & (wr )  ;
assign n7034 =  ( n7033 ) ? ( n5262 ) : ( iram_7 ) ;
assign n7035 = wr_addr[7:7] ;
assign n7036 =  ( n7035 ) == ( bv_1_0_n53 )  ;
assign n7037 =  ( wr_addr ) == ( bv_8_7_n83 )  ;
assign n7038 =  ( n7036 ) & (n7037 )  ;
assign n7039 =  ( n7038 ) & (wr )  ;
assign n7040 =  ( n7039 ) ? ( n5298 ) : ( iram_7 ) ;
assign n7041 = wr_addr[7:7] ;
assign n7042 =  ( n7041 ) == ( bv_1_0_n53 )  ;
assign n7043 =  ( wr_addr ) == ( bv_8_7_n83 )  ;
assign n7044 =  ( n7042 ) & (n7043 )  ;
assign n7045 =  ( n7044 ) & (wr )  ;
assign n7046 =  ( n7045 ) ? ( n5325 ) : ( iram_7 ) ;
assign n7047 = wr_addr[7:7] ;
assign n7048 =  ( n7047 ) == ( bv_1_0_n53 )  ;
assign n7049 =  ( wr_addr ) == ( bv_8_8_n85 )  ;
assign n7050 =  ( n7048 ) & (n7049 )  ;
assign n7051 =  ( n7050 ) & (wr )  ;
assign n7052 =  ( n7051 ) ? ( n4782 ) : ( iram_8 ) ;
assign n7053 = wr_addr[7:7] ;
assign n7054 =  ( n7053 ) == ( bv_1_0_n53 )  ;
assign n7055 =  ( wr_addr ) == ( bv_8_8_n85 )  ;
assign n7056 =  ( n7054 ) & (n7055 )  ;
assign n7057 =  ( n7056 ) & (wr )  ;
assign n7058 =  ( n7057 ) ? ( n4841 ) : ( iram_8 ) ;
assign n7059 = wr_addr[7:7] ;
assign n7060 =  ( n7059 ) == ( bv_1_0_n53 )  ;
assign n7061 =  ( wr_addr ) == ( bv_8_8_n85 )  ;
assign n7062 =  ( n7060 ) & (n7061 )  ;
assign n7063 =  ( n7062 ) & (wr )  ;
assign n7064 =  ( n7063 ) ? ( n5449 ) : ( iram_8 ) ;
assign n7065 = wr_addr[7:7] ;
assign n7066 =  ( n7065 ) == ( bv_1_0_n53 )  ;
assign n7067 =  ( wr_addr ) == ( bv_8_8_n85 )  ;
assign n7068 =  ( n7066 ) & (n7067 )  ;
assign n7069 =  ( n7068 ) & (wr )  ;
assign n7070 =  ( n7069 ) ? ( n4906 ) : ( iram_8 ) ;
assign n7071 = wr_addr[7:7] ;
assign n7072 =  ( n7071 ) == ( bv_1_0_n53 )  ;
assign n7073 =  ( wr_addr ) == ( bv_8_8_n85 )  ;
assign n7074 =  ( n7072 ) & (n7073 )  ;
assign n7075 =  ( n7074 ) & (wr )  ;
assign n7076 =  ( n7075 ) ? ( n5485 ) : ( iram_8 ) ;
assign n7077 = wr_addr[7:7] ;
assign n7078 =  ( n7077 ) == ( bv_1_0_n53 )  ;
assign n7079 =  ( wr_addr ) == ( bv_8_8_n85 )  ;
assign n7080 =  ( n7078 ) & (n7079 )  ;
assign n7081 =  ( n7080 ) & (wr )  ;
assign n7082 =  ( n7081 ) ? ( n5512 ) : ( iram_8 ) ;
assign n7083 = wr_addr[7:7] ;
assign n7084 =  ( n7083 ) == ( bv_1_0_n53 )  ;
assign n7085 =  ( wr_addr ) == ( bv_8_8_n85 )  ;
assign n7086 =  ( n7084 ) & (n7085 )  ;
assign n7087 =  ( n7086 ) & (wr )  ;
assign n7088 =  ( n7087 ) ? ( bv_8_0_n69 ) : ( iram_8 ) ;
assign n7089 = wr_addr[7:7] ;
assign n7090 =  ( n7089 ) == ( bv_1_0_n53 )  ;
assign n7091 =  ( wr_addr ) == ( bv_8_8_n85 )  ;
assign n7092 =  ( n7090 ) & (n7091 )  ;
assign n7093 =  ( n7092 ) & (wr )  ;
assign n7094 =  ( n7093 ) ? ( n5071 ) : ( iram_8 ) ;
assign n7095 = wr_addr[7:7] ;
assign n7096 =  ( n7095 ) == ( bv_1_0_n53 )  ;
assign n7097 =  ( wr_addr ) == ( bv_8_8_n85 )  ;
assign n7098 =  ( n7096 ) & (n7097 )  ;
assign n7099 =  ( n7098 ) & (wr )  ;
assign n7100 =  ( n7099 ) ? ( n5096 ) : ( iram_8 ) ;
assign n7101 = wr_addr[7:7] ;
assign n7102 =  ( n7101 ) == ( bv_1_0_n53 )  ;
assign n7103 =  ( wr_addr ) == ( bv_8_8_n85 )  ;
assign n7104 =  ( n7102 ) & (n7103 )  ;
assign n7105 =  ( n7104 ) & (wr )  ;
assign n7106 =  ( n7105 ) ? ( n5123 ) : ( iram_8 ) ;
assign n7107 = wr_addr[7:7] ;
assign n7108 =  ( n7107 ) == ( bv_1_0_n53 )  ;
assign n7109 =  ( wr_addr ) == ( bv_8_8_n85 )  ;
assign n7110 =  ( n7108 ) & (n7109 )  ;
assign n7111 =  ( n7110 ) & (wr )  ;
assign n7112 =  ( n7111 ) ? ( n5165 ) : ( iram_8 ) ;
assign n7113 = wr_addr[7:7] ;
assign n7114 =  ( n7113 ) == ( bv_1_0_n53 )  ;
assign n7115 =  ( wr_addr ) == ( bv_8_8_n85 )  ;
assign n7116 =  ( n7114 ) & (n7115 )  ;
assign n7117 =  ( n7116 ) & (wr )  ;
assign n7118 =  ( n7117 ) ? ( n5204 ) : ( iram_8 ) ;
assign n7119 = wr_addr[7:7] ;
assign n7120 =  ( n7119 ) == ( bv_1_0_n53 )  ;
assign n7121 =  ( wr_addr ) == ( bv_8_8_n85 )  ;
assign n7122 =  ( n7120 ) & (n7121 )  ;
assign n7123 =  ( n7122 ) & (wr )  ;
assign n7124 =  ( n7123 ) ? ( n5262 ) : ( iram_8 ) ;
assign n7125 = wr_addr[7:7] ;
assign n7126 =  ( n7125 ) == ( bv_1_0_n53 )  ;
assign n7127 =  ( wr_addr ) == ( bv_8_8_n85 )  ;
assign n7128 =  ( n7126 ) & (n7127 )  ;
assign n7129 =  ( n7128 ) & (wr )  ;
assign n7130 =  ( n7129 ) ? ( n5298 ) : ( iram_8 ) ;
assign n7131 = wr_addr[7:7] ;
assign n7132 =  ( n7131 ) == ( bv_1_0_n53 )  ;
assign n7133 =  ( wr_addr ) == ( bv_8_8_n85 )  ;
assign n7134 =  ( n7132 ) & (n7133 )  ;
assign n7135 =  ( n7134 ) & (wr )  ;
assign n7136 =  ( n7135 ) ? ( n5325 ) : ( iram_8 ) ;
assign n7137 = wr_addr[7:7] ;
assign n7138 =  ( n7137 ) == ( bv_1_0_n53 )  ;
assign n7139 =  ( wr_addr ) == ( bv_8_9_n87 )  ;
assign n7140 =  ( n7138 ) & (n7139 )  ;
assign n7141 =  ( n7140 ) & (wr )  ;
assign n7142 =  ( n7141 ) ? ( n4782 ) : ( iram_9 ) ;
assign n7143 = wr_addr[7:7] ;
assign n7144 =  ( n7143 ) == ( bv_1_0_n53 )  ;
assign n7145 =  ( wr_addr ) == ( bv_8_9_n87 )  ;
assign n7146 =  ( n7144 ) & (n7145 )  ;
assign n7147 =  ( n7146 ) & (wr )  ;
assign n7148 =  ( n7147 ) ? ( n4841 ) : ( iram_9 ) ;
assign n7149 = wr_addr[7:7] ;
assign n7150 =  ( n7149 ) == ( bv_1_0_n53 )  ;
assign n7151 =  ( wr_addr ) == ( bv_8_9_n87 )  ;
assign n7152 =  ( n7150 ) & (n7151 )  ;
assign n7153 =  ( n7152 ) & (wr )  ;
assign n7154 =  ( n7153 ) ? ( n5449 ) : ( iram_9 ) ;
assign n7155 = wr_addr[7:7] ;
assign n7156 =  ( n7155 ) == ( bv_1_0_n53 )  ;
assign n7157 =  ( wr_addr ) == ( bv_8_9_n87 )  ;
assign n7158 =  ( n7156 ) & (n7157 )  ;
assign n7159 =  ( n7158 ) & (wr )  ;
assign n7160 =  ( n7159 ) ? ( n4906 ) : ( iram_9 ) ;
assign n7161 = wr_addr[7:7] ;
assign n7162 =  ( n7161 ) == ( bv_1_0_n53 )  ;
assign n7163 =  ( wr_addr ) == ( bv_8_9_n87 )  ;
assign n7164 =  ( n7162 ) & (n7163 )  ;
assign n7165 =  ( n7164 ) & (wr )  ;
assign n7166 =  ( n7165 ) ? ( n5485 ) : ( iram_9 ) ;
assign n7167 = wr_addr[7:7] ;
assign n7168 =  ( n7167 ) == ( bv_1_0_n53 )  ;
assign n7169 =  ( wr_addr ) == ( bv_8_9_n87 )  ;
assign n7170 =  ( n7168 ) & (n7169 )  ;
assign n7171 =  ( n7170 ) & (wr )  ;
assign n7172 =  ( n7171 ) ? ( n5512 ) : ( iram_9 ) ;
assign n7173 = wr_addr[7:7] ;
assign n7174 =  ( n7173 ) == ( bv_1_0_n53 )  ;
assign n7175 =  ( wr_addr ) == ( bv_8_9_n87 )  ;
assign n7176 =  ( n7174 ) & (n7175 )  ;
assign n7177 =  ( n7176 ) & (wr )  ;
assign n7178 =  ( n7177 ) ? ( bv_8_0_n69 ) : ( iram_9 ) ;
assign n7179 = wr_addr[7:7] ;
assign n7180 =  ( n7179 ) == ( bv_1_0_n53 )  ;
assign n7181 =  ( wr_addr ) == ( bv_8_9_n87 )  ;
assign n7182 =  ( n7180 ) & (n7181 )  ;
assign n7183 =  ( n7182 ) & (wr )  ;
assign n7184 =  ( n7183 ) ? ( n5071 ) : ( iram_9 ) ;
assign n7185 = wr_addr[7:7] ;
assign n7186 =  ( n7185 ) == ( bv_1_0_n53 )  ;
assign n7187 =  ( wr_addr ) == ( bv_8_9_n87 )  ;
assign n7188 =  ( n7186 ) & (n7187 )  ;
assign n7189 =  ( n7188 ) & (wr )  ;
assign n7190 =  ( n7189 ) ? ( n5096 ) : ( iram_9 ) ;
assign n7191 = wr_addr[7:7] ;
assign n7192 =  ( n7191 ) == ( bv_1_0_n53 )  ;
assign n7193 =  ( wr_addr ) == ( bv_8_9_n87 )  ;
assign n7194 =  ( n7192 ) & (n7193 )  ;
assign n7195 =  ( n7194 ) & (wr )  ;
assign n7196 =  ( n7195 ) ? ( n5123 ) : ( iram_9 ) ;
assign n7197 = wr_addr[7:7] ;
assign n7198 =  ( n7197 ) == ( bv_1_0_n53 )  ;
assign n7199 =  ( wr_addr ) == ( bv_8_9_n87 )  ;
assign n7200 =  ( n7198 ) & (n7199 )  ;
assign n7201 =  ( n7200 ) & (wr )  ;
assign n7202 =  ( n7201 ) ? ( n5165 ) : ( iram_9 ) ;
assign n7203 = wr_addr[7:7] ;
assign n7204 =  ( n7203 ) == ( bv_1_0_n53 )  ;
assign n7205 =  ( wr_addr ) == ( bv_8_9_n87 )  ;
assign n7206 =  ( n7204 ) & (n7205 )  ;
assign n7207 =  ( n7206 ) & (wr )  ;
assign n7208 =  ( n7207 ) ? ( n5204 ) : ( iram_9 ) ;
assign n7209 = wr_addr[7:7] ;
assign n7210 =  ( n7209 ) == ( bv_1_0_n53 )  ;
assign n7211 =  ( wr_addr ) == ( bv_8_9_n87 )  ;
assign n7212 =  ( n7210 ) & (n7211 )  ;
assign n7213 =  ( n7212 ) & (wr )  ;
assign n7214 =  ( n7213 ) ? ( n5262 ) : ( iram_9 ) ;
assign n7215 = wr_addr[7:7] ;
assign n7216 =  ( n7215 ) == ( bv_1_0_n53 )  ;
assign n7217 =  ( wr_addr ) == ( bv_8_9_n87 )  ;
assign n7218 =  ( n7216 ) & (n7217 )  ;
assign n7219 =  ( n7218 ) & (wr )  ;
assign n7220 =  ( n7219 ) ? ( n5298 ) : ( iram_9 ) ;
assign n7221 = wr_addr[7:7] ;
assign n7222 =  ( n7221 ) == ( bv_1_0_n53 )  ;
assign n7223 =  ( wr_addr ) == ( bv_8_9_n87 )  ;
assign n7224 =  ( n7222 ) & (n7223 )  ;
assign n7225 =  ( n7224 ) & (wr )  ;
assign n7226 =  ( n7225 ) ? ( n5325 ) : ( iram_9 ) ;
assign n7227 = wr_addr[7:7] ;
assign n7228 =  ( n7227 ) == ( bv_1_0_n53 )  ;
assign n7229 =  ( wr_addr ) == ( bv_8_10_n89 )  ;
assign n7230 =  ( n7228 ) & (n7229 )  ;
assign n7231 =  ( n7230 ) & (wr )  ;
assign n7232 =  ( n7231 ) ? ( n4782 ) : ( iram_10 ) ;
assign n7233 = wr_addr[7:7] ;
assign n7234 =  ( n7233 ) == ( bv_1_0_n53 )  ;
assign n7235 =  ( wr_addr ) == ( bv_8_10_n89 )  ;
assign n7236 =  ( n7234 ) & (n7235 )  ;
assign n7237 =  ( n7236 ) & (wr )  ;
assign n7238 =  ( n7237 ) ? ( n4841 ) : ( iram_10 ) ;
assign n7239 = wr_addr[7:7] ;
assign n7240 =  ( n7239 ) == ( bv_1_0_n53 )  ;
assign n7241 =  ( wr_addr ) == ( bv_8_10_n89 )  ;
assign n7242 =  ( n7240 ) & (n7241 )  ;
assign n7243 =  ( n7242 ) & (wr )  ;
assign n7244 =  ( n7243 ) ? ( n5449 ) : ( iram_10 ) ;
assign n7245 = wr_addr[7:7] ;
assign n7246 =  ( n7245 ) == ( bv_1_0_n53 )  ;
assign n7247 =  ( wr_addr ) == ( bv_8_10_n89 )  ;
assign n7248 =  ( n7246 ) & (n7247 )  ;
assign n7249 =  ( n7248 ) & (wr )  ;
assign n7250 =  ( n7249 ) ? ( n4906 ) : ( iram_10 ) ;
assign n7251 = wr_addr[7:7] ;
assign n7252 =  ( n7251 ) == ( bv_1_0_n53 )  ;
assign n7253 =  ( wr_addr ) == ( bv_8_10_n89 )  ;
assign n7254 =  ( n7252 ) & (n7253 )  ;
assign n7255 =  ( n7254 ) & (wr )  ;
assign n7256 =  ( n7255 ) ? ( n5485 ) : ( iram_10 ) ;
assign n7257 = wr_addr[7:7] ;
assign n7258 =  ( n7257 ) == ( bv_1_0_n53 )  ;
assign n7259 =  ( wr_addr ) == ( bv_8_10_n89 )  ;
assign n7260 =  ( n7258 ) & (n7259 )  ;
assign n7261 =  ( n7260 ) & (wr )  ;
assign n7262 =  ( n7261 ) ? ( n5512 ) : ( iram_10 ) ;
assign n7263 = wr_addr[7:7] ;
assign n7264 =  ( n7263 ) == ( bv_1_0_n53 )  ;
assign n7265 =  ( wr_addr ) == ( bv_8_10_n89 )  ;
assign n7266 =  ( n7264 ) & (n7265 )  ;
assign n7267 =  ( n7266 ) & (wr )  ;
assign n7268 =  ( n7267 ) ? ( bv_8_0_n69 ) : ( iram_10 ) ;
assign n7269 = wr_addr[7:7] ;
assign n7270 =  ( n7269 ) == ( bv_1_0_n53 )  ;
assign n7271 =  ( wr_addr ) == ( bv_8_10_n89 )  ;
assign n7272 =  ( n7270 ) & (n7271 )  ;
assign n7273 =  ( n7272 ) & (wr )  ;
assign n7274 =  ( n7273 ) ? ( n5071 ) : ( iram_10 ) ;
assign n7275 = wr_addr[7:7] ;
assign n7276 =  ( n7275 ) == ( bv_1_0_n53 )  ;
assign n7277 =  ( wr_addr ) == ( bv_8_10_n89 )  ;
assign n7278 =  ( n7276 ) & (n7277 )  ;
assign n7279 =  ( n7278 ) & (wr )  ;
assign n7280 =  ( n7279 ) ? ( n5096 ) : ( iram_10 ) ;
assign n7281 = wr_addr[7:7] ;
assign n7282 =  ( n7281 ) == ( bv_1_0_n53 )  ;
assign n7283 =  ( wr_addr ) == ( bv_8_10_n89 )  ;
assign n7284 =  ( n7282 ) & (n7283 )  ;
assign n7285 =  ( n7284 ) & (wr )  ;
assign n7286 =  ( n7285 ) ? ( n5123 ) : ( iram_10 ) ;
assign n7287 = wr_addr[7:7] ;
assign n7288 =  ( n7287 ) == ( bv_1_0_n53 )  ;
assign n7289 =  ( wr_addr ) == ( bv_8_10_n89 )  ;
assign n7290 =  ( n7288 ) & (n7289 )  ;
assign n7291 =  ( n7290 ) & (wr )  ;
assign n7292 =  ( n7291 ) ? ( n5165 ) : ( iram_10 ) ;
assign n7293 = wr_addr[7:7] ;
assign n7294 =  ( n7293 ) == ( bv_1_0_n53 )  ;
assign n7295 =  ( wr_addr ) == ( bv_8_10_n89 )  ;
assign n7296 =  ( n7294 ) & (n7295 )  ;
assign n7297 =  ( n7296 ) & (wr )  ;
assign n7298 =  ( n7297 ) ? ( n5204 ) : ( iram_10 ) ;
assign n7299 = wr_addr[7:7] ;
assign n7300 =  ( n7299 ) == ( bv_1_0_n53 )  ;
assign n7301 =  ( wr_addr ) == ( bv_8_10_n89 )  ;
assign n7302 =  ( n7300 ) & (n7301 )  ;
assign n7303 =  ( n7302 ) & (wr )  ;
assign n7304 =  ( n7303 ) ? ( n5262 ) : ( iram_10 ) ;
assign n7305 = wr_addr[7:7] ;
assign n7306 =  ( n7305 ) == ( bv_1_0_n53 )  ;
assign n7307 =  ( wr_addr ) == ( bv_8_10_n89 )  ;
assign n7308 =  ( n7306 ) & (n7307 )  ;
assign n7309 =  ( n7308 ) & (wr )  ;
assign n7310 =  ( n7309 ) ? ( n5298 ) : ( iram_10 ) ;
assign n7311 = wr_addr[7:7] ;
assign n7312 =  ( n7311 ) == ( bv_1_0_n53 )  ;
assign n7313 =  ( wr_addr ) == ( bv_8_10_n89 )  ;
assign n7314 =  ( n7312 ) & (n7313 )  ;
assign n7315 =  ( n7314 ) & (wr )  ;
assign n7316 =  ( n7315 ) ? ( n5325 ) : ( iram_10 ) ;
assign n7317 = wr_addr[7:7] ;
assign n7318 =  ( n7317 ) == ( bv_1_0_n53 )  ;
assign n7319 =  ( wr_addr ) == ( bv_8_11_n91 )  ;
assign n7320 =  ( n7318 ) & (n7319 )  ;
assign n7321 =  ( n7320 ) & (wr )  ;
assign n7322 =  ( n7321 ) ? ( n4782 ) : ( iram_11 ) ;
assign n7323 = wr_addr[7:7] ;
assign n7324 =  ( n7323 ) == ( bv_1_0_n53 )  ;
assign n7325 =  ( wr_addr ) == ( bv_8_11_n91 )  ;
assign n7326 =  ( n7324 ) & (n7325 )  ;
assign n7327 =  ( n7326 ) & (wr )  ;
assign n7328 =  ( n7327 ) ? ( n4841 ) : ( iram_11 ) ;
assign n7329 = wr_addr[7:7] ;
assign n7330 =  ( n7329 ) == ( bv_1_0_n53 )  ;
assign n7331 =  ( wr_addr ) == ( bv_8_11_n91 )  ;
assign n7332 =  ( n7330 ) & (n7331 )  ;
assign n7333 =  ( n7332 ) & (wr )  ;
assign n7334 =  ( n7333 ) ? ( n5449 ) : ( iram_11 ) ;
assign n7335 = wr_addr[7:7] ;
assign n7336 =  ( n7335 ) == ( bv_1_0_n53 )  ;
assign n7337 =  ( wr_addr ) == ( bv_8_11_n91 )  ;
assign n7338 =  ( n7336 ) & (n7337 )  ;
assign n7339 =  ( n7338 ) & (wr )  ;
assign n7340 =  ( n7339 ) ? ( n4906 ) : ( iram_11 ) ;
assign n7341 = wr_addr[7:7] ;
assign n7342 =  ( n7341 ) == ( bv_1_0_n53 )  ;
assign n7343 =  ( wr_addr ) == ( bv_8_11_n91 )  ;
assign n7344 =  ( n7342 ) & (n7343 )  ;
assign n7345 =  ( n7344 ) & (wr )  ;
assign n7346 =  ( n7345 ) ? ( n5485 ) : ( iram_11 ) ;
assign n7347 = wr_addr[7:7] ;
assign n7348 =  ( n7347 ) == ( bv_1_0_n53 )  ;
assign n7349 =  ( wr_addr ) == ( bv_8_11_n91 )  ;
assign n7350 =  ( n7348 ) & (n7349 )  ;
assign n7351 =  ( n7350 ) & (wr )  ;
assign n7352 =  ( n7351 ) ? ( n5512 ) : ( iram_11 ) ;
assign n7353 = wr_addr[7:7] ;
assign n7354 =  ( n7353 ) == ( bv_1_0_n53 )  ;
assign n7355 =  ( wr_addr ) == ( bv_8_11_n91 )  ;
assign n7356 =  ( n7354 ) & (n7355 )  ;
assign n7357 =  ( n7356 ) & (wr )  ;
assign n7358 =  ( n7357 ) ? ( bv_8_0_n69 ) : ( iram_11 ) ;
assign n7359 = wr_addr[7:7] ;
assign n7360 =  ( n7359 ) == ( bv_1_0_n53 )  ;
assign n7361 =  ( wr_addr ) == ( bv_8_11_n91 )  ;
assign n7362 =  ( n7360 ) & (n7361 )  ;
assign n7363 =  ( n7362 ) & (wr )  ;
assign n7364 =  ( n7363 ) ? ( n5071 ) : ( iram_11 ) ;
assign n7365 = wr_addr[7:7] ;
assign n7366 =  ( n7365 ) == ( bv_1_0_n53 )  ;
assign n7367 =  ( wr_addr ) == ( bv_8_11_n91 )  ;
assign n7368 =  ( n7366 ) & (n7367 )  ;
assign n7369 =  ( n7368 ) & (wr )  ;
assign n7370 =  ( n7369 ) ? ( n5096 ) : ( iram_11 ) ;
assign n7371 = wr_addr[7:7] ;
assign n7372 =  ( n7371 ) == ( bv_1_0_n53 )  ;
assign n7373 =  ( wr_addr ) == ( bv_8_11_n91 )  ;
assign n7374 =  ( n7372 ) & (n7373 )  ;
assign n7375 =  ( n7374 ) & (wr )  ;
assign n7376 =  ( n7375 ) ? ( n5123 ) : ( iram_11 ) ;
assign n7377 = wr_addr[7:7] ;
assign n7378 =  ( n7377 ) == ( bv_1_0_n53 )  ;
assign n7379 =  ( wr_addr ) == ( bv_8_11_n91 )  ;
assign n7380 =  ( n7378 ) & (n7379 )  ;
assign n7381 =  ( n7380 ) & (wr )  ;
assign n7382 =  ( n7381 ) ? ( n5165 ) : ( iram_11 ) ;
assign n7383 = wr_addr[7:7] ;
assign n7384 =  ( n7383 ) == ( bv_1_0_n53 )  ;
assign n7385 =  ( wr_addr ) == ( bv_8_11_n91 )  ;
assign n7386 =  ( n7384 ) & (n7385 )  ;
assign n7387 =  ( n7386 ) & (wr )  ;
assign n7388 =  ( n7387 ) ? ( n5204 ) : ( iram_11 ) ;
assign n7389 = wr_addr[7:7] ;
assign n7390 =  ( n7389 ) == ( bv_1_0_n53 )  ;
assign n7391 =  ( wr_addr ) == ( bv_8_11_n91 )  ;
assign n7392 =  ( n7390 ) & (n7391 )  ;
assign n7393 =  ( n7392 ) & (wr )  ;
assign n7394 =  ( n7393 ) ? ( n5262 ) : ( iram_11 ) ;
assign n7395 = wr_addr[7:7] ;
assign n7396 =  ( n7395 ) == ( bv_1_0_n53 )  ;
assign n7397 =  ( wr_addr ) == ( bv_8_11_n91 )  ;
assign n7398 =  ( n7396 ) & (n7397 )  ;
assign n7399 =  ( n7398 ) & (wr )  ;
assign n7400 =  ( n7399 ) ? ( n5298 ) : ( iram_11 ) ;
assign n7401 = wr_addr[7:7] ;
assign n7402 =  ( n7401 ) == ( bv_1_0_n53 )  ;
assign n7403 =  ( wr_addr ) == ( bv_8_11_n91 )  ;
assign n7404 =  ( n7402 ) & (n7403 )  ;
assign n7405 =  ( n7404 ) & (wr )  ;
assign n7406 =  ( n7405 ) ? ( n5325 ) : ( iram_11 ) ;
assign n7407 = wr_addr[7:7] ;
assign n7408 =  ( n7407 ) == ( bv_1_0_n53 )  ;
assign n7409 =  ( wr_addr ) == ( bv_8_12_n93 )  ;
assign n7410 =  ( n7408 ) & (n7409 )  ;
assign n7411 =  ( n7410 ) & (wr )  ;
assign n7412 =  ( n7411 ) ? ( n4782 ) : ( iram_12 ) ;
assign n7413 = wr_addr[7:7] ;
assign n7414 =  ( n7413 ) == ( bv_1_0_n53 )  ;
assign n7415 =  ( wr_addr ) == ( bv_8_12_n93 )  ;
assign n7416 =  ( n7414 ) & (n7415 )  ;
assign n7417 =  ( n7416 ) & (wr )  ;
assign n7418 =  ( n7417 ) ? ( n4841 ) : ( iram_12 ) ;
assign n7419 = wr_addr[7:7] ;
assign n7420 =  ( n7419 ) == ( bv_1_0_n53 )  ;
assign n7421 =  ( wr_addr ) == ( bv_8_12_n93 )  ;
assign n7422 =  ( n7420 ) & (n7421 )  ;
assign n7423 =  ( n7422 ) & (wr )  ;
assign n7424 =  ( n7423 ) ? ( n5449 ) : ( iram_12 ) ;
assign n7425 = wr_addr[7:7] ;
assign n7426 =  ( n7425 ) == ( bv_1_0_n53 )  ;
assign n7427 =  ( wr_addr ) == ( bv_8_12_n93 )  ;
assign n7428 =  ( n7426 ) & (n7427 )  ;
assign n7429 =  ( n7428 ) & (wr )  ;
assign n7430 =  ( n7429 ) ? ( n4906 ) : ( iram_12 ) ;
assign n7431 = wr_addr[7:7] ;
assign n7432 =  ( n7431 ) == ( bv_1_0_n53 )  ;
assign n7433 =  ( wr_addr ) == ( bv_8_12_n93 )  ;
assign n7434 =  ( n7432 ) & (n7433 )  ;
assign n7435 =  ( n7434 ) & (wr )  ;
assign n7436 =  ( n7435 ) ? ( n5485 ) : ( iram_12 ) ;
assign n7437 = wr_addr[7:7] ;
assign n7438 =  ( n7437 ) == ( bv_1_0_n53 )  ;
assign n7439 =  ( wr_addr ) == ( bv_8_12_n93 )  ;
assign n7440 =  ( n7438 ) & (n7439 )  ;
assign n7441 =  ( n7440 ) & (wr )  ;
assign n7442 =  ( n7441 ) ? ( n5512 ) : ( iram_12 ) ;
assign n7443 = wr_addr[7:7] ;
assign n7444 =  ( n7443 ) == ( bv_1_0_n53 )  ;
assign n7445 =  ( wr_addr ) == ( bv_8_12_n93 )  ;
assign n7446 =  ( n7444 ) & (n7445 )  ;
assign n7447 =  ( n7446 ) & (wr )  ;
assign n7448 =  ( n7447 ) ? ( bv_8_0_n69 ) : ( iram_12 ) ;
assign n7449 = wr_addr[7:7] ;
assign n7450 =  ( n7449 ) == ( bv_1_0_n53 )  ;
assign n7451 =  ( wr_addr ) == ( bv_8_12_n93 )  ;
assign n7452 =  ( n7450 ) & (n7451 )  ;
assign n7453 =  ( n7452 ) & (wr )  ;
assign n7454 =  ( n7453 ) ? ( n5071 ) : ( iram_12 ) ;
assign n7455 = wr_addr[7:7] ;
assign n7456 =  ( n7455 ) == ( bv_1_0_n53 )  ;
assign n7457 =  ( wr_addr ) == ( bv_8_12_n93 )  ;
assign n7458 =  ( n7456 ) & (n7457 )  ;
assign n7459 =  ( n7458 ) & (wr )  ;
assign n7460 =  ( n7459 ) ? ( n5096 ) : ( iram_12 ) ;
assign n7461 = wr_addr[7:7] ;
assign n7462 =  ( n7461 ) == ( bv_1_0_n53 )  ;
assign n7463 =  ( wr_addr ) == ( bv_8_12_n93 )  ;
assign n7464 =  ( n7462 ) & (n7463 )  ;
assign n7465 =  ( n7464 ) & (wr )  ;
assign n7466 =  ( n7465 ) ? ( n5123 ) : ( iram_12 ) ;
assign n7467 = wr_addr[7:7] ;
assign n7468 =  ( n7467 ) == ( bv_1_0_n53 )  ;
assign n7469 =  ( wr_addr ) == ( bv_8_12_n93 )  ;
assign n7470 =  ( n7468 ) & (n7469 )  ;
assign n7471 =  ( n7470 ) & (wr )  ;
assign n7472 =  ( n7471 ) ? ( n5165 ) : ( iram_12 ) ;
assign n7473 = wr_addr[7:7] ;
assign n7474 =  ( n7473 ) == ( bv_1_0_n53 )  ;
assign n7475 =  ( wr_addr ) == ( bv_8_12_n93 )  ;
assign n7476 =  ( n7474 ) & (n7475 )  ;
assign n7477 =  ( n7476 ) & (wr )  ;
assign n7478 =  ( n7477 ) ? ( n5204 ) : ( iram_12 ) ;
assign n7479 = wr_addr[7:7] ;
assign n7480 =  ( n7479 ) == ( bv_1_0_n53 )  ;
assign n7481 =  ( wr_addr ) == ( bv_8_12_n93 )  ;
assign n7482 =  ( n7480 ) & (n7481 )  ;
assign n7483 =  ( n7482 ) & (wr )  ;
assign n7484 =  ( n7483 ) ? ( n5262 ) : ( iram_12 ) ;
assign n7485 = wr_addr[7:7] ;
assign n7486 =  ( n7485 ) == ( bv_1_0_n53 )  ;
assign n7487 =  ( wr_addr ) == ( bv_8_12_n93 )  ;
assign n7488 =  ( n7486 ) & (n7487 )  ;
assign n7489 =  ( n7488 ) & (wr )  ;
assign n7490 =  ( n7489 ) ? ( n5298 ) : ( iram_12 ) ;
assign n7491 = wr_addr[7:7] ;
assign n7492 =  ( n7491 ) == ( bv_1_0_n53 )  ;
assign n7493 =  ( wr_addr ) == ( bv_8_12_n93 )  ;
assign n7494 =  ( n7492 ) & (n7493 )  ;
assign n7495 =  ( n7494 ) & (wr )  ;
assign n7496 =  ( n7495 ) ? ( n5325 ) : ( iram_12 ) ;
assign n7497 = wr_addr[7:7] ;
assign n7498 =  ( n7497 ) == ( bv_1_0_n53 )  ;
assign n7499 =  ( wr_addr ) == ( bv_8_13_n95 )  ;
assign n7500 =  ( n7498 ) & (n7499 )  ;
assign n7501 =  ( n7500 ) & (wr )  ;
assign n7502 =  ( n7501 ) ? ( n4782 ) : ( iram_13 ) ;
assign n7503 = wr_addr[7:7] ;
assign n7504 =  ( n7503 ) == ( bv_1_0_n53 )  ;
assign n7505 =  ( wr_addr ) == ( bv_8_13_n95 )  ;
assign n7506 =  ( n7504 ) & (n7505 )  ;
assign n7507 =  ( n7506 ) & (wr )  ;
assign n7508 =  ( n7507 ) ? ( n4841 ) : ( iram_13 ) ;
assign n7509 = wr_addr[7:7] ;
assign n7510 =  ( n7509 ) == ( bv_1_0_n53 )  ;
assign n7511 =  ( wr_addr ) == ( bv_8_13_n95 )  ;
assign n7512 =  ( n7510 ) & (n7511 )  ;
assign n7513 =  ( n7512 ) & (wr )  ;
assign n7514 =  ( n7513 ) ? ( n5449 ) : ( iram_13 ) ;
assign n7515 = wr_addr[7:7] ;
assign n7516 =  ( n7515 ) == ( bv_1_0_n53 )  ;
assign n7517 =  ( wr_addr ) == ( bv_8_13_n95 )  ;
assign n7518 =  ( n7516 ) & (n7517 )  ;
assign n7519 =  ( n7518 ) & (wr )  ;
assign n7520 =  ( n7519 ) ? ( n4906 ) : ( iram_13 ) ;
assign n7521 = wr_addr[7:7] ;
assign n7522 =  ( n7521 ) == ( bv_1_0_n53 )  ;
assign n7523 =  ( wr_addr ) == ( bv_8_13_n95 )  ;
assign n7524 =  ( n7522 ) & (n7523 )  ;
assign n7525 =  ( n7524 ) & (wr )  ;
assign n7526 =  ( n7525 ) ? ( n5485 ) : ( iram_13 ) ;
assign n7527 = wr_addr[7:7] ;
assign n7528 =  ( n7527 ) == ( bv_1_0_n53 )  ;
assign n7529 =  ( wr_addr ) == ( bv_8_13_n95 )  ;
assign n7530 =  ( n7528 ) & (n7529 )  ;
assign n7531 =  ( n7530 ) & (wr )  ;
assign n7532 =  ( n7531 ) ? ( n5512 ) : ( iram_13 ) ;
assign n7533 = wr_addr[7:7] ;
assign n7534 =  ( n7533 ) == ( bv_1_0_n53 )  ;
assign n7535 =  ( wr_addr ) == ( bv_8_13_n95 )  ;
assign n7536 =  ( n7534 ) & (n7535 )  ;
assign n7537 =  ( n7536 ) & (wr )  ;
assign n7538 =  ( n7537 ) ? ( bv_8_0_n69 ) : ( iram_13 ) ;
assign n7539 = wr_addr[7:7] ;
assign n7540 =  ( n7539 ) == ( bv_1_0_n53 )  ;
assign n7541 =  ( wr_addr ) == ( bv_8_13_n95 )  ;
assign n7542 =  ( n7540 ) & (n7541 )  ;
assign n7543 =  ( n7542 ) & (wr )  ;
assign n7544 =  ( n7543 ) ? ( n5071 ) : ( iram_13 ) ;
assign n7545 = wr_addr[7:7] ;
assign n7546 =  ( n7545 ) == ( bv_1_0_n53 )  ;
assign n7547 =  ( wr_addr ) == ( bv_8_13_n95 )  ;
assign n7548 =  ( n7546 ) & (n7547 )  ;
assign n7549 =  ( n7548 ) & (wr )  ;
assign n7550 =  ( n7549 ) ? ( n5096 ) : ( iram_13 ) ;
assign n7551 = wr_addr[7:7] ;
assign n7552 =  ( n7551 ) == ( bv_1_0_n53 )  ;
assign n7553 =  ( wr_addr ) == ( bv_8_13_n95 )  ;
assign n7554 =  ( n7552 ) & (n7553 )  ;
assign n7555 =  ( n7554 ) & (wr )  ;
assign n7556 =  ( n7555 ) ? ( n5123 ) : ( iram_13 ) ;
assign n7557 = wr_addr[7:7] ;
assign n7558 =  ( n7557 ) == ( bv_1_0_n53 )  ;
assign n7559 =  ( wr_addr ) == ( bv_8_13_n95 )  ;
assign n7560 =  ( n7558 ) & (n7559 )  ;
assign n7561 =  ( n7560 ) & (wr )  ;
assign n7562 =  ( n7561 ) ? ( n5165 ) : ( iram_13 ) ;
assign n7563 = wr_addr[7:7] ;
assign n7564 =  ( n7563 ) == ( bv_1_0_n53 )  ;
assign n7565 =  ( wr_addr ) == ( bv_8_13_n95 )  ;
assign n7566 =  ( n7564 ) & (n7565 )  ;
assign n7567 =  ( n7566 ) & (wr )  ;
assign n7568 =  ( n7567 ) ? ( n5204 ) : ( iram_13 ) ;
assign n7569 = wr_addr[7:7] ;
assign n7570 =  ( n7569 ) == ( bv_1_0_n53 )  ;
assign n7571 =  ( wr_addr ) == ( bv_8_13_n95 )  ;
assign n7572 =  ( n7570 ) & (n7571 )  ;
assign n7573 =  ( n7572 ) & (wr )  ;
assign n7574 =  ( n7573 ) ? ( n5262 ) : ( iram_13 ) ;
assign n7575 = wr_addr[7:7] ;
assign n7576 =  ( n7575 ) == ( bv_1_0_n53 )  ;
assign n7577 =  ( wr_addr ) == ( bv_8_13_n95 )  ;
assign n7578 =  ( n7576 ) & (n7577 )  ;
assign n7579 =  ( n7578 ) & (wr )  ;
assign n7580 =  ( n7579 ) ? ( n5298 ) : ( iram_13 ) ;
assign n7581 = wr_addr[7:7] ;
assign n7582 =  ( n7581 ) == ( bv_1_0_n53 )  ;
assign n7583 =  ( wr_addr ) == ( bv_8_13_n95 )  ;
assign n7584 =  ( n7582 ) & (n7583 )  ;
assign n7585 =  ( n7584 ) & (wr )  ;
assign n7586 =  ( n7585 ) ? ( n5325 ) : ( iram_13 ) ;
assign n7587 = wr_addr[7:7] ;
assign n7588 =  ( n7587 ) == ( bv_1_0_n53 )  ;
assign n7589 =  ( wr_addr ) == ( bv_8_14_n97 )  ;
assign n7590 =  ( n7588 ) & (n7589 )  ;
assign n7591 =  ( n7590 ) & (wr )  ;
assign n7592 =  ( n7591 ) ? ( n4782 ) : ( iram_14 ) ;
assign n7593 = wr_addr[7:7] ;
assign n7594 =  ( n7593 ) == ( bv_1_0_n53 )  ;
assign n7595 =  ( wr_addr ) == ( bv_8_14_n97 )  ;
assign n7596 =  ( n7594 ) & (n7595 )  ;
assign n7597 =  ( n7596 ) & (wr )  ;
assign n7598 =  ( n7597 ) ? ( n4841 ) : ( iram_14 ) ;
assign n7599 = wr_addr[7:7] ;
assign n7600 =  ( n7599 ) == ( bv_1_0_n53 )  ;
assign n7601 =  ( wr_addr ) == ( bv_8_14_n97 )  ;
assign n7602 =  ( n7600 ) & (n7601 )  ;
assign n7603 =  ( n7602 ) & (wr )  ;
assign n7604 =  ( n7603 ) ? ( n5449 ) : ( iram_14 ) ;
assign n7605 = wr_addr[7:7] ;
assign n7606 =  ( n7605 ) == ( bv_1_0_n53 )  ;
assign n7607 =  ( wr_addr ) == ( bv_8_14_n97 )  ;
assign n7608 =  ( n7606 ) & (n7607 )  ;
assign n7609 =  ( n7608 ) & (wr )  ;
assign n7610 =  ( n7609 ) ? ( n4906 ) : ( iram_14 ) ;
assign n7611 = wr_addr[7:7] ;
assign n7612 =  ( n7611 ) == ( bv_1_0_n53 )  ;
assign n7613 =  ( wr_addr ) == ( bv_8_14_n97 )  ;
assign n7614 =  ( n7612 ) & (n7613 )  ;
assign n7615 =  ( n7614 ) & (wr )  ;
assign n7616 =  ( n7615 ) ? ( n5485 ) : ( iram_14 ) ;
assign n7617 = wr_addr[7:7] ;
assign n7618 =  ( n7617 ) == ( bv_1_0_n53 )  ;
assign n7619 =  ( wr_addr ) == ( bv_8_14_n97 )  ;
assign n7620 =  ( n7618 ) & (n7619 )  ;
assign n7621 =  ( n7620 ) & (wr )  ;
assign n7622 =  ( n7621 ) ? ( n5512 ) : ( iram_14 ) ;
assign n7623 = wr_addr[7:7] ;
assign n7624 =  ( n7623 ) == ( bv_1_0_n53 )  ;
assign n7625 =  ( wr_addr ) == ( bv_8_14_n97 )  ;
assign n7626 =  ( n7624 ) & (n7625 )  ;
assign n7627 =  ( n7626 ) & (wr )  ;
assign n7628 =  ( n7627 ) ? ( bv_8_0_n69 ) : ( iram_14 ) ;
assign n7629 = wr_addr[7:7] ;
assign n7630 =  ( n7629 ) == ( bv_1_0_n53 )  ;
assign n7631 =  ( wr_addr ) == ( bv_8_14_n97 )  ;
assign n7632 =  ( n7630 ) & (n7631 )  ;
assign n7633 =  ( n7632 ) & (wr )  ;
assign n7634 =  ( n7633 ) ? ( n5071 ) : ( iram_14 ) ;
assign n7635 = wr_addr[7:7] ;
assign n7636 =  ( n7635 ) == ( bv_1_0_n53 )  ;
assign n7637 =  ( wr_addr ) == ( bv_8_14_n97 )  ;
assign n7638 =  ( n7636 ) & (n7637 )  ;
assign n7639 =  ( n7638 ) & (wr )  ;
assign n7640 =  ( n7639 ) ? ( n5096 ) : ( iram_14 ) ;
assign n7641 = wr_addr[7:7] ;
assign n7642 =  ( n7641 ) == ( bv_1_0_n53 )  ;
assign n7643 =  ( wr_addr ) == ( bv_8_14_n97 )  ;
assign n7644 =  ( n7642 ) & (n7643 )  ;
assign n7645 =  ( n7644 ) & (wr )  ;
assign n7646 =  ( n7645 ) ? ( n5123 ) : ( iram_14 ) ;
assign n7647 = wr_addr[7:7] ;
assign n7648 =  ( n7647 ) == ( bv_1_0_n53 )  ;
assign n7649 =  ( wr_addr ) == ( bv_8_14_n97 )  ;
assign n7650 =  ( n7648 ) & (n7649 )  ;
assign n7651 =  ( n7650 ) & (wr )  ;
assign n7652 =  ( n7651 ) ? ( n5165 ) : ( iram_14 ) ;
assign n7653 = wr_addr[7:7] ;
assign n7654 =  ( n7653 ) == ( bv_1_0_n53 )  ;
assign n7655 =  ( wr_addr ) == ( bv_8_14_n97 )  ;
assign n7656 =  ( n7654 ) & (n7655 )  ;
assign n7657 =  ( n7656 ) & (wr )  ;
assign n7658 =  ( n7657 ) ? ( n5204 ) : ( iram_14 ) ;
assign n7659 = wr_addr[7:7] ;
assign n7660 =  ( n7659 ) == ( bv_1_0_n53 )  ;
assign n7661 =  ( wr_addr ) == ( bv_8_14_n97 )  ;
assign n7662 =  ( n7660 ) & (n7661 )  ;
assign n7663 =  ( n7662 ) & (wr )  ;
assign n7664 =  ( n7663 ) ? ( n5262 ) : ( iram_14 ) ;
assign n7665 = wr_addr[7:7] ;
assign n7666 =  ( n7665 ) == ( bv_1_0_n53 )  ;
assign n7667 =  ( wr_addr ) == ( bv_8_14_n97 )  ;
assign n7668 =  ( n7666 ) & (n7667 )  ;
assign n7669 =  ( n7668 ) & (wr )  ;
assign n7670 =  ( n7669 ) ? ( n5298 ) : ( iram_14 ) ;
assign n7671 = wr_addr[7:7] ;
assign n7672 =  ( n7671 ) == ( bv_1_0_n53 )  ;
assign n7673 =  ( wr_addr ) == ( bv_8_14_n97 )  ;
assign n7674 =  ( n7672 ) & (n7673 )  ;
assign n7675 =  ( n7674 ) & (wr )  ;
assign n7676 =  ( n7675 ) ? ( n5325 ) : ( iram_14 ) ;
assign n7677 = wr_addr[7:7] ;
assign n7678 =  ( n7677 ) == ( bv_1_0_n53 )  ;
assign n7679 =  ( wr_addr ) == ( bv_8_15_n99 )  ;
assign n7680 =  ( n7678 ) & (n7679 )  ;
assign n7681 =  ( n7680 ) & (wr )  ;
assign n7682 =  ( n7681 ) ? ( n4782 ) : ( iram_15 ) ;
assign n7683 = wr_addr[7:7] ;
assign n7684 =  ( n7683 ) == ( bv_1_0_n53 )  ;
assign n7685 =  ( wr_addr ) == ( bv_8_15_n99 )  ;
assign n7686 =  ( n7684 ) & (n7685 )  ;
assign n7687 =  ( n7686 ) & (wr )  ;
assign n7688 =  ( n7687 ) ? ( n4841 ) : ( iram_15 ) ;
assign n7689 = wr_addr[7:7] ;
assign n7690 =  ( n7689 ) == ( bv_1_0_n53 )  ;
assign n7691 =  ( wr_addr ) == ( bv_8_15_n99 )  ;
assign n7692 =  ( n7690 ) & (n7691 )  ;
assign n7693 =  ( n7692 ) & (wr )  ;
assign n7694 =  ( n7693 ) ? ( n5449 ) : ( iram_15 ) ;
assign n7695 = wr_addr[7:7] ;
assign n7696 =  ( n7695 ) == ( bv_1_0_n53 )  ;
assign n7697 =  ( wr_addr ) == ( bv_8_15_n99 )  ;
assign n7698 =  ( n7696 ) & (n7697 )  ;
assign n7699 =  ( n7698 ) & (wr )  ;
assign n7700 =  ( n7699 ) ? ( n4906 ) : ( iram_15 ) ;
assign n7701 = wr_addr[7:7] ;
assign n7702 =  ( n7701 ) == ( bv_1_0_n53 )  ;
assign n7703 =  ( wr_addr ) == ( bv_8_15_n99 )  ;
assign n7704 =  ( n7702 ) & (n7703 )  ;
assign n7705 =  ( n7704 ) & (wr )  ;
assign n7706 =  ( n7705 ) ? ( n5485 ) : ( iram_15 ) ;
assign n7707 = wr_addr[7:7] ;
assign n7708 =  ( n7707 ) == ( bv_1_0_n53 )  ;
assign n7709 =  ( wr_addr ) == ( bv_8_15_n99 )  ;
assign n7710 =  ( n7708 ) & (n7709 )  ;
assign n7711 =  ( n7710 ) & (wr )  ;
assign n7712 =  ( n7711 ) ? ( n5512 ) : ( iram_15 ) ;
assign n7713 = wr_addr[7:7] ;
assign n7714 =  ( n7713 ) == ( bv_1_0_n53 )  ;
assign n7715 =  ( wr_addr ) == ( bv_8_15_n99 )  ;
assign n7716 =  ( n7714 ) & (n7715 )  ;
assign n7717 =  ( n7716 ) & (wr )  ;
assign n7718 =  ( n7717 ) ? ( bv_8_0_n69 ) : ( iram_15 ) ;
assign n7719 = wr_addr[7:7] ;
assign n7720 =  ( n7719 ) == ( bv_1_0_n53 )  ;
assign n7721 =  ( wr_addr ) == ( bv_8_15_n99 )  ;
assign n7722 =  ( n7720 ) & (n7721 )  ;
assign n7723 =  ( n7722 ) & (wr )  ;
assign n7724 =  ( n7723 ) ? ( n5071 ) : ( iram_15 ) ;
assign n7725 = wr_addr[7:7] ;
assign n7726 =  ( n7725 ) == ( bv_1_0_n53 )  ;
assign n7727 =  ( wr_addr ) == ( bv_8_15_n99 )  ;
assign n7728 =  ( n7726 ) & (n7727 )  ;
assign n7729 =  ( n7728 ) & (wr )  ;
assign n7730 =  ( n7729 ) ? ( n5096 ) : ( iram_15 ) ;
assign n7731 = wr_addr[7:7] ;
assign n7732 =  ( n7731 ) == ( bv_1_0_n53 )  ;
assign n7733 =  ( wr_addr ) == ( bv_8_15_n99 )  ;
assign n7734 =  ( n7732 ) & (n7733 )  ;
assign n7735 =  ( n7734 ) & (wr )  ;
assign n7736 =  ( n7735 ) ? ( n5123 ) : ( iram_15 ) ;
assign n7737 = wr_addr[7:7] ;
assign n7738 =  ( n7737 ) == ( bv_1_0_n53 )  ;
assign n7739 =  ( wr_addr ) == ( bv_8_15_n99 )  ;
assign n7740 =  ( n7738 ) & (n7739 )  ;
assign n7741 =  ( n7740 ) & (wr )  ;
assign n7742 =  ( n7741 ) ? ( n5165 ) : ( iram_15 ) ;
assign n7743 = wr_addr[7:7] ;
assign n7744 =  ( n7743 ) == ( bv_1_0_n53 )  ;
assign n7745 =  ( wr_addr ) == ( bv_8_15_n99 )  ;
assign n7746 =  ( n7744 ) & (n7745 )  ;
assign n7747 =  ( n7746 ) & (wr )  ;
assign n7748 =  ( n7747 ) ? ( n5204 ) : ( iram_15 ) ;
assign n7749 = wr_addr[7:7] ;
assign n7750 =  ( n7749 ) == ( bv_1_0_n53 )  ;
assign n7751 =  ( wr_addr ) == ( bv_8_15_n99 )  ;
assign n7752 =  ( n7750 ) & (n7751 )  ;
assign n7753 =  ( n7752 ) & (wr )  ;
assign n7754 =  ( n7753 ) ? ( n5262 ) : ( iram_15 ) ;
assign n7755 = wr_addr[7:7] ;
assign n7756 =  ( n7755 ) == ( bv_1_0_n53 )  ;
assign n7757 =  ( wr_addr ) == ( bv_8_15_n99 )  ;
assign n7758 =  ( n7756 ) & (n7757 )  ;
assign n7759 =  ( n7758 ) & (wr )  ;
assign n7760 =  ( n7759 ) ? ( n5298 ) : ( iram_15 ) ;
assign n7761 = wr_addr[7:7] ;
assign n7762 =  ( n7761 ) == ( bv_1_0_n53 )  ;
assign n7763 =  ( wr_addr ) == ( bv_8_15_n99 )  ;
assign n7764 =  ( n7762 ) & (n7763 )  ;
assign n7765 =  ( n7764 ) & (wr )  ;
assign n7766 =  ( n7765 ) ? ( n5325 ) : ( iram_15 ) ;
assign n7767 = wr_addr[7:7] ;
assign n7768 =  ( n7767 ) == ( bv_1_0_n53 )  ;
assign n7769 =  ( wr_addr ) == ( bv_8_16_n101 )  ;
assign n7770 =  ( n7768 ) & (n7769 )  ;
assign n7771 =  ( n7770 ) & (wr )  ;
assign n7772 =  ( n7771 ) ? ( n4782 ) : ( iram_16 ) ;
assign n7773 = wr_addr[7:7] ;
assign n7774 =  ( n7773 ) == ( bv_1_0_n53 )  ;
assign n7775 =  ( wr_addr ) == ( bv_8_16_n101 )  ;
assign n7776 =  ( n7774 ) & (n7775 )  ;
assign n7777 =  ( n7776 ) & (wr )  ;
assign n7778 =  ( n7777 ) ? ( n4841 ) : ( iram_16 ) ;
assign n7779 = wr_addr[7:7] ;
assign n7780 =  ( n7779 ) == ( bv_1_0_n53 )  ;
assign n7781 =  ( wr_addr ) == ( bv_8_16_n101 )  ;
assign n7782 =  ( n7780 ) & (n7781 )  ;
assign n7783 =  ( n7782 ) & (wr )  ;
assign n7784 =  ( n7783 ) ? ( n5449 ) : ( iram_16 ) ;
assign n7785 = wr_addr[7:7] ;
assign n7786 =  ( n7785 ) == ( bv_1_0_n53 )  ;
assign n7787 =  ( wr_addr ) == ( bv_8_16_n101 )  ;
assign n7788 =  ( n7786 ) & (n7787 )  ;
assign n7789 =  ( n7788 ) & (wr )  ;
assign n7790 =  ( n7789 ) ? ( n4906 ) : ( iram_16 ) ;
assign n7791 = wr_addr[7:7] ;
assign n7792 =  ( n7791 ) == ( bv_1_0_n53 )  ;
assign n7793 =  ( wr_addr ) == ( bv_8_16_n101 )  ;
assign n7794 =  ( n7792 ) & (n7793 )  ;
assign n7795 =  ( n7794 ) & (wr )  ;
assign n7796 =  ( n7795 ) ? ( n5485 ) : ( iram_16 ) ;
assign n7797 = wr_addr[7:7] ;
assign n7798 =  ( n7797 ) == ( bv_1_0_n53 )  ;
assign n7799 =  ( wr_addr ) == ( bv_8_16_n101 )  ;
assign n7800 =  ( n7798 ) & (n7799 )  ;
assign n7801 =  ( n7800 ) & (wr )  ;
assign n7802 =  ( n7801 ) ? ( n5512 ) : ( iram_16 ) ;
assign n7803 = wr_addr[7:7] ;
assign n7804 =  ( n7803 ) == ( bv_1_0_n53 )  ;
assign n7805 =  ( wr_addr ) == ( bv_8_16_n101 )  ;
assign n7806 =  ( n7804 ) & (n7805 )  ;
assign n7807 =  ( n7806 ) & (wr )  ;
assign n7808 =  ( n7807 ) ? ( bv_8_0_n69 ) : ( iram_16 ) ;
assign n7809 = wr_addr[7:7] ;
assign n7810 =  ( n7809 ) == ( bv_1_0_n53 )  ;
assign n7811 =  ( wr_addr ) == ( bv_8_16_n101 )  ;
assign n7812 =  ( n7810 ) & (n7811 )  ;
assign n7813 =  ( n7812 ) & (wr )  ;
assign n7814 =  ( n7813 ) ? ( n5071 ) : ( iram_16 ) ;
assign n7815 = wr_addr[7:7] ;
assign n7816 =  ( n7815 ) == ( bv_1_0_n53 )  ;
assign n7817 =  ( wr_addr ) == ( bv_8_16_n101 )  ;
assign n7818 =  ( n7816 ) & (n7817 )  ;
assign n7819 =  ( n7818 ) & (wr )  ;
assign n7820 =  ( n7819 ) ? ( n5096 ) : ( iram_16 ) ;
assign n7821 = wr_addr[7:7] ;
assign n7822 =  ( n7821 ) == ( bv_1_0_n53 )  ;
assign n7823 =  ( wr_addr ) == ( bv_8_16_n101 )  ;
assign n7824 =  ( n7822 ) & (n7823 )  ;
assign n7825 =  ( n7824 ) & (wr )  ;
assign n7826 =  ( n7825 ) ? ( n5123 ) : ( iram_16 ) ;
assign n7827 = wr_addr[7:7] ;
assign n7828 =  ( n7827 ) == ( bv_1_0_n53 )  ;
assign n7829 =  ( wr_addr ) == ( bv_8_16_n101 )  ;
assign n7830 =  ( n7828 ) & (n7829 )  ;
assign n7831 =  ( n7830 ) & (wr )  ;
assign n7832 =  ( n7831 ) ? ( n5165 ) : ( iram_16 ) ;
assign n7833 = wr_addr[7:7] ;
assign n7834 =  ( n7833 ) == ( bv_1_0_n53 )  ;
assign n7835 =  ( wr_addr ) == ( bv_8_16_n101 )  ;
assign n7836 =  ( n7834 ) & (n7835 )  ;
assign n7837 =  ( n7836 ) & (wr )  ;
assign n7838 =  ( n7837 ) ? ( n5204 ) : ( iram_16 ) ;
assign n7839 = wr_addr[7:7] ;
assign n7840 =  ( n7839 ) == ( bv_1_0_n53 )  ;
assign n7841 =  ( wr_addr ) == ( bv_8_16_n101 )  ;
assign n7842 =  ( n7840 ) & (n7841 )  ;
assign n7843 =  ( n7842 ) & (wr )  ;
assign n7844 =  ( n7843 ) ? ( n5262 ) : ( iram_16 ) ;
assign n7845 = wr_addr[7:7] ;
assign n7846 =  ( n7845 ) == ( bv_1_0_n53 )  ;
assign n7847 =  ( wr_addr ) == ( bv_8_16_n101 )  ;
assign n7848 =  ( n7846 ) & (n7847 )  ;
assign n7849 =  ( n7848 ) & (wr )  ;
assign n7850 =  ( n7849 ) ? ( n5298 ) : ( iram_16 ) ;
assign n7851 = wr_addr[7:7] ;
assign n7852 =  ( n7851 ) == ( bv_1_0_n53 )  ;
assign n7853 =  ( wr_addr ) == ( bv_8_16_n101 )  ;
assign n7854 =  ( n7852 ) & (n7853 )  ;
assign n7855 =  ( n7854 ) & (wr )  ;
assign n7856 =  ( n7855 ) ? ( n5325 ) : ( iram_16 ) ;
assign n7857 = wr_addr[7:7] ;
assign n7858 =  ( n7857 ) == ( bv_1_0_n53 )  ;
assign n7859 =  ( wr_addr ) == ( bv_8_17_n103 )  ;
assign n7860 =  ( n7858 ) & (n7859 )  ;
assign n7861 =  ( n7860 ) & (wr )  ;
assign n7862 =  ( n7861 ) ? ( n4782 ) : ( iram_17 ) ;
assign n7863 = wr_addr[7:7] ;
assign n7864 =  ( n7863 ) == ( bv_1_0_n53 )  ;
assign n7865 =  ( wr_addr ) == ( bv_8_17_n103 )  ;
assign n7866 =  ( n7864 ) & (n7865 )  ;
assign n7867 =  ( n7866 ) & (wr )  ;
assign n7868 =  ( n7867 ) ? ( n4841 ) : ( iram_17 ) ;
assign n7869 = wr_addr[7:7] ;
assign n7870 =  ( n7869 ) == ( bv_1_0_n53 )  ;
assign n7871 =  ( wr_addr ) == ( bv_8_17_n103 )  ;
assign n7872 =  ( n7870 ) & (n7871 )  ;
assign n7873 =  ( n7872 ) & (wr )  ;
assign n7874 =  ( n7873 ) ? ( n5449 ) : ( iram_17 ) ;
assign n7875 = wr_addr[7:7] ;
assign n7876 =  ( n7875 ) == ( bv_1_0_n53 )  ;
assign n7877 =  ( wr_addr ) == ( bv_8_17_n103 )  ;
assign n7878 =  ( n7876 ) & (n7877 )  ;
assign n7879 =  ( n7878 ) & (wr )  ;
assign n7880 =  ( n7879 ) ? ( n4906 ) : ( iram_17 ) ;
assign n7881 = wr_addr[7:7] ;
assign n7882 =  ( n7881 ) == ( bv_1_0_n53 )  ;
assign n7883 =  ( wr_addr ) == ( bv_8_17_n103 )  ;
assign n7884 =  ( n7882 ) & (n7883 )  ;
assign n7885 =  ( n7884 ) & (wr )  ;
assign n7886 =  ( n7885 ) ? ( n5485 ) : ( iram_17 ) ;
assign n7887 = wr_addr[7:7] ;
assign n7888 =  ( n7887 ) == ( bv_1_0_n53 )  ;
assign n7889 =  ( wr_addr ) == ( bv_8_17_n103 )  ;
assign n7890 =  ( n7888 ) & (n7889 )  ;
assign n7891 =  ( n7890 ) & (wr )  ;
assign n7892 =  ( n7891 ) ? ( n5512 ) : ( iram_17 ) ;
assign n7893 = wr_addr[7:7] ;
assign n7894 =  ( n7893 ) == ( bv_1_0_n53 )  ;
assign n7895 =  ( wr_addr ) == ( bv_8_17_n103 )  ;
assign n7896 =  ( n7894 ) & (n7895 )  ;
assign n7897 =  ( n7896 ) & (wr )  ;
assign n7898 =  ( n7897 ) ? ( bv_8_0_n69 ) : ( iram_17 ) ;
assign n7899 = wr_addr[7:7] ;
assign n7900 =  ( n7899 ) == ( bv_1_0_n53 )  ;
assign n7901 =  ( wr_addr ) == ( bv_8_17_n103 )  ;
assign n7902 =  ( n7900 ) & (n7901 )  ;
assign n7903 =  ( n7902 ) & (wr )  ;
assign n7904 =  ( n7903 ) ? ( n5071 ) : ( iram_17 ) ;
assign n7905 = wr_addr[7:7] ;
assign n7906 =  ( n7905 ) == ( bv_1_0_n53 )  ;
assign n7907 =  ( wr_addr ) == ( bv_8_17_n103 )  ;
assign n7908 =  ( n7906 ) & (n7907 )  ;
assign n7909 =  ( n7908 ) & (wr )  ;
assign n7910 =  ( n7909 ) ? ( n5096 ) : ( iram_17 ) ;
assign n7911 = wr_addr[7:7] ;
assign n7912 =  ( n7911 ) == ( bv_1_0_n53 )  ;
assign n7913 =  ( wr_addr ) == ( bv_8_17_n103 )  ;
assign n7914 =  ( n7912 ) & (n7913 )  ;
assign n7915 =  ( n7914 ) & (wr )  ;
assign n7916 =  ( n7915 ) ? ( n5123 ) : ( iram_17 ) ;
assign n7917 = wr_addr[7:7] ;
assign n7918 =  ( n7917 ) == ( bv_1_0_n53 )  ;
assign n7919 =  ( wr_addr ) == ( bv_8_17_n103 )  ;
assign n7920 =  ( n7918 ) & (n7919 )  ;
assign n7921 =  ( n7920 ) & (wr )  ;
assign n7922 =  ( n7921 ) ? ( n5165 ) : ( iram_17 ) ;
assign n7923 = wr_addr[7:7] ;
assign n7924 =  ( n7923 ) == ( bv_1_0_n53 )  ;
assign n7925 =  ( wr_addr ) == ( bv_8_17_n103 )  ;
assign n7926 =  ( n7924 ) & (n7925 )  ;
assign n7927 =  ( n7926 ) & (wr )  ;
assign n7928 =  ( n7927 ) ? ( n5204 ) : ( iram_17 ) ;
assign n7929 = wr_addr[7:7] ;
assign n7930 =  ( n7929 ) == ( bv_1_0_n53 )  ;
assign n7931 =  ( wr_addr ) == ( bv_8_17_n103 )  ;
assign n7932 =  ( n7930 ) & (n7931 )  ;
assign n7933 =  ( n7932 ) & (wr )  ;
assign n7934 =  ( n7933 ) ? ( n5262 ) : ( iram_17 ) ;
assign n7935 = wr_addr[7:7] ;
assign n7936 =  ( n7935 ) == ( bv_1_0_n53 )  ;
assign n7937 =  ( wr_addr ) == ( bv_8_17_n103 )  ;
assign n7938 =  ( n7936 ) & (n7937 )  ;
assign n7939 =  ( n7938 ) & (wr )  ;
assign n7940 =  ( n7939 ) ? ( n5298 ) : ( iram_17 ) ;
assign n7941 = wr_addr[7:7] ;
assign n7942 =  ( n7941 ) == ( bv_1_0_n53 )  ;
assign n7943 =  ( wr_addr ) == ( bv_8_17_n103 )  ;
assign n7944 =  ( n7942 ) & (n7943 )  ;
assign n7945 =  ( n7944 ) & (wr )  ;
assign n7946 =  ( n7945 ) ? ( n5325 ) : ( iram_17 ) ;
assign n7947 = wr_addr[7:7] ;
assign n7948 =  ( n7947 ) == ( bv_1_0_n53 )  ;
assign n7949 =  ( wr_addr ) == ( bv_8_18_n105 )  ;
assign n7950 =  ( n7948 ) & (n7949 )  ;
assign n7951 =  ( n7950 ) & (wr )  ;
assign n7952 =  ( n7951 ) ? ( n4782 ) : ( iram_18 ) ;
assign n7953 = wr_addr[7:7] ;
assign n7954 =  ( n7953 ) == ( bv_1_0_n53 )  ;
assign n7955 =  ( wr_addr ) == ( bv_8_18_n105 )  ;
assign n7956 =  ( n7954 ) & (n7955 )  ;
assign n7957 =  ( n7956 ) & (wr )  ;
assign n7958 =  ( n7957 ) ? ( n4841 ) : ( iram_18 ) ;
assign n7959 = wr_addr[7:7] ;
assign n7960 =  ( n7959 ) == ( bv_1_0_n53 )  ;
assign n7961 =  ( wr_addr ) == ( bv_8_18_n105 )  ;
assign n7962 =  ( n7960 ) & (n7961 )  ;
assign n7963 =  ( n7962 ) & (wr )  ;
assign n7964 =  ( n7963 ) ? ( n5449 ) : ( iram_18 ) ;
assign n7965 = wr_addr[7:7] ;
assign n7966 =  ( n7965 ) == ( bv_1_0_n53 )  ;
assign n7967 =  ( wr_addr ) == ( bv_8_18_n105 )  ;
assign n7968 =  ( n7966 ) & (n7967 )  ;
assign n7969 =  ( n7968 ) & (wr )  ;
assign n7970 =  ( n7969 ) ? ( n4906 ) : ( iram_18 ) ;
assign n7971 = wr_addr[7:7] ;
assign n7972 =  ( n7971 ) == ( bv_1_0_n53 )  ;
assign n7973 =  ( wr_addr ) == ( bv_8_18_n105 )  ;
assign n7974 =  ( n7972 ) & (n7973 )  ;
assign n7975 =  ( n7974 ) & (wr )  ;
assign n7976 =  ( n7975 ) ? ( n5485 ) : ( iram_18 ) ;
assign n7977 = wr_addr[7:7] ;
assign n7978 =  ( n7977 ) == ( bv_1_0_n53 )  ;
assign n7979 =  ( wr_addr ) == ( bv_8_18_n105 )  ;
assign n7980 =  ( n7978 ) & (n7979 )  ;
assign n7981 =  ( n7980 ) & (wr )  ;
assign n7982 =  ( n7981 ) ? ( n5512 ) : ( iram_18 ) ;
assign n7983 = wr_addr[7:7] ;
assign n7984 =  ( n7983 ) == ( bv_1_0_n53 )  ;
assign n7985 =  ( wr_addr ) == ( bv_8_18_n105 )  ;
assign n7986 =  ( n7984 ) & (n7985 )  ;
assign n7987 =  ( n7986 ) & (wr )  ;
assign n7988 =  ( n7987 ) ? ( bv_8_0_n69 ) : ( iram_18 ) ;
assign n7989 = wr_addr[7:7] ;
assign n7990 =  ( n7989 ) == ( bv_1_0_n53 )  ;
assign n7991 =  ( wr_addr ) == ( bv_8_18_n105 )  ;
assign n7992 =  ( n7990 ) & (n7991 )  ;
assign n7993 =  ( n7992 ) & (wr )  ;
assign n7994 =  ( n7993 ) ? ( n5071 ) : ( iram_18 ) ;
assign n7995 = wr_addr[7:7] ;
assign n7996 =  ( n7995 ) == ( bv_1_0_n53 )  ;
assign n7997 =  ( wr_addr ) == ( bv_8_18_n105 )  ;
assign n7998 =  ( n7996 ) & (n7997 )  ;
assign n7999 =  ( n7998 ) & (wr )  ;
assign n8000 =  ( n7999 ) ? ( n5096 ) : ( iram_18 ) ;
assign n8001 = wr_addr[7:7] ;
assign n8002 =  ( n8001 ) == ( bv_1_0_n53 )  ;
assign n8003 =  ( wr_addr ) == ( bv_8_18_n105 )  ;
assign n8004 =  ( n8002 ) & (n8003 )  ;
assign n8005 =  ( n8004 ) & (wr )  ;
assign n8006 =  ( n8005 ) ? ( n5123 ) : ( iram_18 ) ;
assign n8007 = wr_addr[7:7] ;
assign n8008 =  ( n8007 ) == ( bv_1_0_n53 )  ;
assign n8009 =  ( wr_addr ) == ( bv_8_18_n105 )  ;
assign n8010 =  ( n8008 ) & (n8009 )  ;
assign n8011 =  ( n8010 ) & (wr )  ;
assign n8012 =  ( n8011 ) ? ( n5165 ) : ( iram_18 ) ;
assign n8013 = wr_addr[7:7] ;
assign n8014 =  ( n8013 ) == ( bv_1_0_n53 )  ;
assign n8015 =  ( wr_addr ) == ( bv_8_18_n105 )  ;
assign n8016 =  ( n8014 ) & (n8015 )  ;
assign n8017 =  ( n8016 ) & (wr )  ;
assign n8018 =  ( n8017 ) ? ( n5204 ) : ( iram_18 ) ;
assign n8019 = wr_addr[7:7] ;
assign n8020 =  ( n8019 ) == ( bv_1_0_n53 )  ;
assign n8021 =  ( wr_addr ) == ( bv_8_18_n105 )  ;
assign n8022 =  ( n8020 ) & (n8021 )  ;
assign n8023 =  ( n8022 ) & (wr )  ;
assign n8024 =  ( n8023 ) ? ( n5262 ) : ( iram_18 ) ;
assign n8025 = wr_addr[7:7] ;
assign n8026 =  ( n8025 ) == ( bv_1_0_n53 )  ;
assign n8027 =  ( wr_addr ) == ( bv_8_18_n105 )  ;
assign n8028 =  ( n8026 ) & (n8027 )  ;
assign n8029 =  ( n8028 ) & (wr )  ;
assign n8030 =  ( n8029 ) ? ( n5298 ) : ( iram_18 ) ;
assign n8031 = wr_addr[7:7] ;
assign n8032 =  ( n8031 ) == ( bv_1_0_n53 )  ;
assign n8033 =  ( wr_addr ) == ( bv_8_18_n105 )  ;
assign n8034 =  ( n8032 ) & (n8033 )  ;
assign n8035 =  ( n8034 ) & (wr )  ;
assign n8036 =  ( n8035 ) ? ( n5325 ) : ( iram_18 ) ;
assign n8037 = wr_addr[7:7] ;
assign n8038 =  ( n8037 ) == ( bv_1_0_n53 )  ;
assign n8039 =  ( wr_addr ) == ( bv_8_19_n107 )  ;
assign n8040 =  ( n8038 ) & (n8039 )  ;
assign n8041 =  ( n8040 ) & (wr )  ;
assign n8042 =  ( n8041 ) ? ( n4782 ) : ( iram_19 ) ;
assign n8043 = wr_addr[7:7] ;
assign n8044 =  ( n8043 ) == ( bv_1_0_n53 )  ;
assign n8045 =  ( wr_addr ) == ( bv_8_19_n107 )  ;
assign n8046 =  ( n8044 ) & (n8045 )  ;
assign n8047 =  ( n8046 ) & (wr )  ;
assign n8048 =  ( n8047 ) ? ( n4841 ) : ( iram_19 ) ;
assign n8049 = wr_addr[7:7] ;
assign n8050 =  ( n8049 ) == ( bv_1_0_n53 )  ;
assign n8051 =  ( wr_addr ) == ( bv_8_19_n107 )  ;
assign n8052 =  ( n8050 ) & (n8051 )  ;
assign n8053 =  ( n8052 ) & (wr )  ;
assign n8054 =  ( n8053 ) ? ( n5449 ) : ( iram_19 ) ;
assign n8055 = wr_addr[7:7] ;
assign n8056 =  ( n8055 ) == ( bv_1_0_n53 )  ;
assign n8057 =  ( wr_addr ) == ( bv_8_19_n107 )  ;
assign n8058 =  ( n8056 ) & (n8057 )  ;
assign n8059 =  ( n8058 ) & (wr )  ;
assign n8060 =  ( n8059 ) ? ( n4906 ) : ( iram_19 ) ;
assign n8061 = wr_addr[7:7] ;
assign n8062 =  ( n8061 ) == ( bv_1_0_n53 )  ;
assign n8063 =  ( wr_addr ) == ( bv_8_19_n107 )  ;
assign n8064 =  ( n8062 ) & (n8063 )  ;
assign n8065 =  ( n8064 ) & (wr )  ;
assign n8066 =  ( n8065 ) ? ( n5485 ) : ( iram_19 ) ;
assign n8067 = wr_addr[7:7] ;
assign n8068 =  ( n8067 ) == ( bv_1_0_n53 )  ;
assign n8069 =  ( wr_addr ) == ( bv_8_19_n107 )  ;
assign n8070 =  ( n8068 ) & (n8069 )  ;
assign n8071 =  ( n8070 ) & (wr )  ;
assign n8072 =  ( n8071 ) ? ( n5512 ) : ( iram_19 ) ;
assign n8073 = wr_addr[7:7] ;
assign n8074 =  ( n8073 ) == ( bv_1_0_n53 )  ;
assign n8075 =  ( wr_addr ) == ( bv_8_19_n107 )  ;
assign n8076 =  ( n8074 ) & (n8075 )  ;
assign n8077 =  ( n8076 ) & (wr )  ;
assign n8078 =  ( n8077 ) ? ( bv_8_0_n69 ) : ( iram_19 ) ;
assign n8079 = wr_addr[7:7] ;
assign n8080 =  ( n8079 ) == ( bv_1_0_n53 )  ;
assign n8081 =  ( wr_addr ) == ( bv_8_19_n107 )  ;
assign n8082 =  ( n8080 ) & (n8081 )  ;
assign n8083 =  ( n8082 ) & (wr )  ;
assign n8084 =  ( n8083 ) ? ( n5071 ) : ( iram_19 ) ;
assign n8085 = wr_addr[7:7] ;
assign n8086 =  ( n8085 ) == ( bv_1_0_n53 )  ;
assign n8087 =  ( wr_addr ) == ( bv_8_19_n107 )  ;
assign n8088 =  ( n8086 ) & (n8087 )  ;
assign n8089 =  ( n8088 ) & (wr )  ;
assign n8090 =  ( n8089 ) ? ( n5096 ) : ( iram_19 ) ;
assign n8091 = wr_addr[7:7] ;
assign n8092 =  ( n8091 ) == ( bv_1_0_n53 )  ;
assign n8093 =  ( wr_addr ) == ( bv_8_19_n107 )  ;
assign n8094 =  ( n8092 ) & (n8093 )  ;
assign n8095 =  ( n8094 ) & (wr )  ;
assign n8096 =  ( n8095 ) ? ( n5123 ) : ( iram_19 ) ;
assign n8097 = wr_addr[7:7] ;
assign n8098 =  ( n8097 ) == ( bv_1_0_n53 )  ;
assign n8099 =  ( wr_addr ) == ( bv_8_19_n107 )  ;
assign n8100 =  ( n8098 ) & (n8099 )  ;
assign n8101 =  ( n8100 ) & (wr )  ;
assign n8102 =  ( n8101 ) ? ( n5165 ) : ( iram_19 ) ;
assign n8103 = wr_addr[7:7] ;
assign n8104 =  ( n8103 ) == ( bv_1_0_n53 )  ;
assign n8105 =  ( wr_addr ) == ( bv_8_19_n107 )  ;
assign n8106 =  ( n8104 ) & (n8105 )  ;
assign n8107 =  ( n8106 ) & (wr )  ;
assign n8108 =  ( n8107 ) ? ( n5204 ) : ( iram_19 ) ;
assign n8109 = wr_addr[7:7] ;
assign n8110 =  ( n8109 ) == ( bv_1_0_n53 )  ;
assign n8111 =  ( wr_addr ) == ( bv_8_19_n107 )  ;
assign n8112 =  ( n8110 ) & (n8111 )  ;
assign n8113 =  ( n8112 ) & (wr )  ;
assign n8114 =  ( n8113 ) ? ( n5262 ) : ( iram_19 ) ;
assign n8115 = wr_addr[7:7] ;
assign n8116 =  ( n8115 ) == ( bv_1_0_n53 )  ;
assign n8117 =  ( wr_addr ) == ( bv_8_19_n107 )  ;
assign n8118 =  ( n8116 ) & (n8117 )  ;
assign n8119 =  ( n8118 ) & (wr )  ;
assign n8120 =  ( n8119 ) ? ( n5298 ) : ( iram_19 ) ;
assign n8121 = wr_addr[7:7] ;
assign n8122 =  ( n8121 ) == ( bv_1_0_n53 )  ;
assign n8123 =  ( wr_addr ) == ( bv_8_19_n107 )  ;
assign n8124 =  ( n8122 ) & (n8123 )  ;
assign n8125 =  ( n8124 ) & (wr )  ;
assign n8126 =  ( n8125 ) ? ( n5325 ) : ( iram_19 ) ;
assign n8127 = wr_addr[7:7] ;
assign n8128 =  ( n8127 ) == ( bv_1_0_n53 )  ;
assign n8129 =  ( wr_addr ) == ( bv_8_20_n109 )  ;
assign n8130 =  ( n8128 ) & (n8129 )  ;
assign n8131 =  ( n8130 ) & (wr )  ;
assign n8132 =  ( n8131 ) ? ( n4782 ) : ( iram_20 ) ;
assign n8133 = wr_addr[7:7] ;
assign n8134 =  ( n8133 ) == ( bv_1_0_n53 )  ;
assign n8135 =  ( wr_addr ) == ( bv_8_20_n109 )  ;
assign n8136 =  ( n8134 ) & (n8135 )  ;
assign n8137 =  ( n8136 ) & (wr )  ;
assign n8138 =  ( n8137 ) ? ( n4841 ) : ( iram_20 ) ;
assign n8139 = wr_addr[7:7] ;
assign n8140 =  ( n8139 ) == ( bv_1_0_n53 )  ;
assign n8141 =  ( wr_addr ) == ( bv_8_20_n109 )  ;
assign n8142 =  ( n8140 ) & (n8141 )  ;
assign n8143 =  ( n8142 ) & (wr )  ;
assign n8144 =  ( n8143 ) ? ( n5449 ) : ( iram_20 ) ;
assign n8145 = wr_addr[7:7] ;
assign n8146 =  ( n8145 ) == ( bv_1_0_n53 )  ;
assign n8147 =  ( wr_addr ) == ( bv_8_20_n109 )  ;
assign n8148 =  ( n8146 ) & (n8147 )  ;
assign n8149 =  ( n8148 ) & (wr )  ;
assign n8150 =  ( n8149 ) ? ( n4906 ) : ( iram_20 ) ;
assign n8151 = wr_addr[7:7] ;
assign n8152 =  ( n8151 ) == ( bv_1_0_n53 )  ;
assign n8153 =  ( wr_addr ) == ( bv_8_20_n109 )  ;
assign n8154 =  ( n8152 ) & (n8153 )  ;
assign n8155 =  ( n8154 ) & (wr )  ;
assign n8156 =  ( n8155 ) ? ( n5485 ) : ( iram_20 ) ;
assign n8157 = wr_addr[7:7] ;
assign n8158 =  ( n8157 ) == ( bv_1_0_n53 )  ;
assign n8159 =  ( wr_addr ) == ( bv_8_20_n109 )  ;
assign n8160 =  ( n8158 ) & (n8159 )  ;
assign n8161 =  ( n8160 ) & (wr )  ;
assign n8162 =  ( n8161 ) ? ( n5512 ) : ( iram_20 ) ;
assign n8163 = wr_addr[7:7] ;
assign n8164 =  ( n8163 ) == ( bv_1_0_n53 )  ;
assign n8165 =  ( wr_addr ) == ( bv_8_20_n109 )  ;
assign n8166 =  ( n8164 ) & (n8165 )  ;
assign n8167 =  ( n8166 ) & (wr )  ;
assign n8168 =  ( n8167 ) ? ( bv_8_0_n69 ) : ( iram_20 ) ;
assign n8169 = wr_addr[7:7] ;
assign n8170 =  ( n8169 ) == ( bv_1_0_n53 )  ;
assign n8171 =  ( wr_addr ) == ( bv_8_20_n109 )  ;
assign n8172 =  ( n8170 ) & (n8171 )  ;
assign n8173 =  ( n8172 ) & (wr )  ;
assign n8174 =  ( n8173 ) ? ( n5071 ) : ( iram_20 ) ;
assign n8175 = wr_addr[7:7] ;
assign n8176 =  ( n8175 ) == ( bv_1_0_n53 )  ;
assign n8177 =  ( wr_addr ) == ( bv_8_20_n109 )  ;
assign n8178 =  ( n8176 ) & (n8177 )  ;
assign n8179 =  ( n8178 ) & (wr )  ;
assign n8180 =  ( n8179 ) ? ( n5096 ) : ( iram_20 ) ;
assign n8181 = wr_addr[7:7] ;
assign n8182 =  ( n8181 ) == ( bv_1_0_n53 )  ;
assign n8183 =  ( wr_addr ) == ( bv_8_20_n109 )  ;
assign n8184 =  ( n8182 ) & (n8183 )  ;
assign n8185 =  ( n8184 ) & (wr )  ;
assign n8186 =  ( n8185 ) ? ( n5123 ) : ( iram_20 ) ;
assign n8187 = wr_addr[7:7] ;
assign n8188 =  ( n8187 ) == ( bv_1_0_n53 )  ;
assign n8189 =  ( wr_addr ) == ( bv_8_20_n109 )  ;
assign n8190 =  ( n8188 ) & (n8189 )  ;
assign n8191 =  ( n8190 ) & (wr )  ;
assign n8192 =  ( n8191 ) ? ( n5165 ) : ( iram_20 ) ;
assign n8193 = wr_addr[7:7] ;
assign n8194 =  ( n8193 ) == ( bv_1_0_n53 )  ;
assign n8195 =  ( wr_addr ) == ( bv_8_20_n109 )  ;
assign n8196 =  ( n8194 ) & (n8195 )  ;
assign n8197 =  ( n8196 ) & (wr )  ;
assign n8198 =  ( n8197 ) ? ( n5204 ) : ( iram_20 ) ;
assign n8199 = wr_addr[7:7] ;
assign n8200 =  ( n8199 ) == ( bv_1_0_n53 )  ;
assign n8201 =  ( wr_addr ) == ( bv_8_20_n109 )  ;
assign n8202 =  ( n8200 ) & (n8201 )  ;
assign n8203 =  ( n8202 ) & (wr )  ;
assign n8204 =  ( n8203 ) ? ( n5262 ) : ( iram_20 ) ;
assign n8205 = wr_addr[7:7] ;
assign n8206 =  ( n8205 ) == ( bv_1_0_n53 )  ;
assign n8207 =  ( wr_addr ) == ( bv_8_20_n109 )  ;
assign n8208 =  ( n8206 ) & (n8207 )  ;
assign n8209 =  ( n8208 ) & (wr )  ;
assign n8210 =  ( n8209 ) ? ( n5298 ) : ( iram_20 ) ;
assign n8211 = wr_addr[7:7] ;
assign n8212 =  ( n8211 ) == ( bv_1_0_n53 )  ;
assign n8213 =  ( wr_addr ) == ( bv_8_20_n109 )  ;
assign n8214 =  ( n8212 ) & (n8213 )  ;
assign n8215 =  ( n8214 ) & (wr )  ;
assign n8216 =  ( n8215 ) ? ( n5325 ) : ( iram_20 ) ;
assign n8217 = wr_addr[7:7] ;
assign n8218 =  ( n8217 ) == ( bv_1_0_n53 )  ;
assign n8219 =  ( wr_addr ) == ( bv_8_21_n111 )  ;
assign n8220 =  ( n8218 ) & (n8219 )  ;
assign n8221 =  ( n8220 ) & (wr )  ;
assign n8222 =  ( n8221 ) ? ( n4782 ) : ( iram_21 ) ;
assign n8223 = wr_addr[7:7] ;
assign n8224 =  ( n8223 ) == ( bv_1_0_n53 )  ;
assign n8225 =  ( wr_addr ) == ( bv_8_21_n111 )  ;
assign n8226 =  ( n8224 ) & (n8225 )  ;
assign n8227 =  ( n8226 ) & (wr )  ;
assign n8228 =  ( n8227 ) ? ( n4841 ) : ( iram_21 ) ;
assign n8229 = wr_addr[7:7] ;
assign n8230 =  ( n8229 ) == ( bv_1_0_n53 )  ;
assign n8231 =  ( wr_addr ) == ( bv_8_21_n111 )  ;
assign n8232 =  ( n8230 ) & (n8231 )  ;
assign n8233 =  ( n8232 ) & (wr )  ;
assign n8234 =  ( n8233 ) ? ( n5449 ) : ( iram_21 ) ;
assign n8235 = wr_addr[7:7] ;
assign n8236 =  ( n8235 ) == ( bv_1_0_n53 )  ;
assign n8237 =  ( wr_addr ) == ( bv_8_21_n111 )  ;
assign n8238 =  ( n8236 ) & (n8237 )  ;
assign n8239 =  ( n8238 ) & (wr )  ;
assign n8240 =  ( n8239 ) ? ( n4906 ) : ( iram_21 ) ;
assign n8241 = wr_addr[7:7] ;
assign n8242 =  ( n8241 ) == ( bv_1_0_n53 )  ;
assign n8243 =  ( wr_addr ) == ( bv_8_21_n111 )  ;
assign n8244 =  ( n8242 ) & (n8243 )  ;
assign n8245 =  ( n8244 ) & (wr )  ;
assign n8246 =  ( n8245 ) ? ( n5485 ) : ( iram_21 ) ;
assign n8247 = wr_addr[7:7] ;
assign n8248 =  ( n8247 ) == ( bv_1_0_n53 )  ;
assign n8249 =  ( wr_addr ) == ( bv_8_21_n111 )  ;
assign n8250 =  ( n8248 ) & (n8249 )  ;
assign n8251 =  ( n8250 ) & (wr )  ;
assign n8252 =  ( n8251 ) ? ( n5512 ) : ( iram_21 ) ;
assign n8253 = wr_addr[7:7] ;
assign n8254 =  ( n8253 ) == ( bv_1_0_n53 )  ;
assign n8255 =  ( wr_addr ) == ( bv_8_21_n111 )  ;
assign n8256 =  ( n8254 ) & (n8255 )  ;
assign n8257 =  ( n8256 ) & (wr )  ;
assign n8258 =  ( n8257 ) ? ( bv_8_0_n69 ) : ( iram_21 ) ;
assign n8259 = wr_addr[7:7] ;
assign n8260 =  ( n8259 ) == ( bv_1_0_n53 )  ;
assign n8261 =  ( wr_addr ) == ( bv_8_21_n111 )  ;
assign n8262 =  ( n8260 ) & (n8261 )  ;
assign n8263 =  ( n8262 ) & (wr )  ;
assign n8264 =  ( n8263 ) ? ( n5071 ) : ( iram_21 ) ;
assign n8265 = wr_addr[7:7] ;
assign n8266 =  ( n8265 ) == ( bv_1_0_n53 )  ;
assign n8267 =  ( wr_addr ) == ( bv_8_21_n111 )  ;
assign n8268 =  ( n8266 ) & (n8267 )  ;
assign n8269 =  ( n8268 ) & (wr )  ;
assign n8270 =  ( n8269 ) ? ( n5096 ) : ( iram_21 ) ;
assign n8271 = wr_addr[7:7] ;
assign n8272 =  ( n8271 ) == ( bv_1_0_n53 )  ;
assign n8273 =  ( wr_addr ) == ( bv_8_21_n111 )  ;
assign n8274 =  ( n8272 ) & (n8273 )  ;
assign n8275 =  ( n8274 ) & (wr )  ;
assign n8276 =  ( n8275 ) ? ( n5123 ) : ( iram_21 ) ;
assign n8277 = wr_addr[7:7] ;
assign n8278 =  ( n8277 ) == ( bv_1_0_n53 )  ;
assign n8279 =  ( wr_addr ) == ( bv_8_21_n111 )  ;
assign n8280 =  ( n8278 ) & (n8279 )  ;
assign n8281 =  ( n8280 ) & (wr )  ;
assign n8282 =  ( n8281 ) ? ( n5165 ) : ( iram_21 ) ;
assign n8283 = wr_addr[7:7] ;
assign n8284 =  ( n8283 ) == ( bv_1_0_n53 )  ;
assign n8285 =  ( wr_addr ) == ( bv_8_21_n111 )  ;
assign n8286 =  ( n8284 ) & (n8285 )  ;
assign n8287 =  ( n8286 ) & (wr )  ;
assign n8288 =  ( n8287 ) ? ( n5204 ) : ( iram_21 ) ;
assign n8289 = wr_addr[7:7] ;
assign n8290 =  ( n8289 ) == ( bv_1_0_n53 )  ;
assign n8291 =  ( wr_addr ) == ( bv_8_21_n111 )  ;
assign n8292 =  ( n8290 ) & (n8291 )  ;
assign n8293 =  ( n8292 ) & (wr )  ;
assign n8294 =  ( n8293 ) ? ( n5262 ) : ( iram_21 ) ;
assign n8295 = wr_addr[7:7] ;
assign n8296 =  ( n8295 ) == ( bv_1_0_n53 )  ;
assign n8297 =  ( wr_addr ) == ( bv_8_21_n111 )  ;
assign n8298 =  ( n8296 ) & (n8297 )  ;
assign n8299 =  ( n8298 ) & (wr )  ;
assign n8300 =  ( n8299 ) ? ( n5298 ) : ( iram_21 ) ;
assign n8301 = wr_addr[7:7] ;
assign n8302 =  ( n8301 ) == ( bv_1_0_n53 )  ;
assign n8303 =  ( wr_addr ) == ( bv_8_21_n111 )  ;
assign n8304 =  ( n8302 ) & (n8303 )  ;
assign n8305 =  ( n8304 ) & (wr )  ;
assign n8306 =  ( n8305 ) ? ( n5325 ) : ( iram_21 ) ;
assign n8307 = wr_addr[7:7] ;
assign n8308 =  ( n8307 ) == ( bv_1_0_n53 )  ;
assign n8309 =  ( wr_addr ) == ( bv_8_22_n113 )  ;
assign n8310 =  ( n8308 ) & (n8309 )  ;
assign n8311 =  ( n8310 ) & (wr )  ;
assign n8312 =  ( n8311 ) ? ( n4782 ) : ( iram_22 ) ;
assign n8313 = wr_addr[7:7] ;
assign n8314 =  ( n8313 ) == ( bv_1_0_n53 )  ;
assign n8315 =  ( wr_addr ) == ( bv_8_22_n113 )  ;
assign n8316 =  ( n8314 ) & (n8315 )  ;
assign n8317 =  ( n8316 ) & (wr )  ;
assign n8318 =  ( n8317 ) ? ( n4841 ) : ( iram_22 ) ;
assign n8319 = wr_addr[7:7] ;
assign n8320 =  ( n8319 ) == ( bv_1_0_n53 )  ;
assign n8321 =  ( wr_addr ) == ( bv_8_22_n113 )  ;
assign n8322 =  ( n8320 ) & (n8321 )  ;
assign n8323 =  ( n8322 ) & (wr )  ;
assign n8324 =  ( n8323 ) ? ( n5449 ) : ( iram_22 ) ;
assign n8325 = wr_addr[7:7] ;
assign n8326 =  ( n8325 ) == ( bv_1_0_n53 )  ;
assign n8327 =  ( wr_addr ) == ( bv_8_22_n113 )  ;
assign n8328 =  ( n8326 ) & (n8327 )  ;
assign n8329 =  ( n8328 ) & (wr )  ;
assign n8330 =  ( n8329 ) ? ( n4906 ) : ( iram_22 ) ;
assign n8331 = wr_addr[7:7] ;
assign n8332 =  ( n8331 ) == ( bv_1_0_n53 )  ;
assign n8333 =  ( wr_addr ) == ( bv_8_22_n113 )  ;
assign n8334 =  ( n8332 ) & (n8333 )  ;
assign n8335 =  ( n8334 ) & (wr )  ;
assign n8336 =  ( n8335 ) ? ( n5485 ) : ( iram_22 ) ;
assign n8337 = wr_addr[7:7] ;
assign n8338 =  ( n8337 ) == ( bv_1_0_n53 )  ;
assign n8339 =  ( wr_addr ) == ( bv_8_22_n113 )  ;
assign n8340 =  ( n8338 ) & (n8339 )  ;
assign n8341 =  ( n8340 ) & (wr )  ;
assign n8342 =  ( n8341 ) ? ( n5512 ) : ( iram_22 ) ;
assign n8343 = wr_addr[7:7] ;
assign n8344 =  ( n8343 ) == ( bv_1_0_n53 )  ;
assign n8345 =  ( wr_addr ) == ( bv_8_22_n113 )  ;
assign n8346 =  ( n8344 ) & (n8345 )  ;
assign n8347 =  ( n8346 ) & (wr )  ;
assign n8348 =  ( n8347 ) ? ( bv_8_0_n69 ) : ( iram_22 ) ;
assign n8349 = wr_addr[7:7] ;
assign n8350 =  ( n8349 ) == ( bv_1_0_n53 )  ;
assign n8351 =  ( wr_addr ) == ( bv_8_22_n113 )  ;
assign n8352 =  ( n8350 ) & (n8351 )  ;
assign n8353 =  ( n8352 ) & (wr )  ;
assign n8354 =  ( n8353 ) ? ( n5071 ) : ( iram_22 ) ;
assign n8355 = wr_addr[7:7] ;
assign n8356 =  ( n8355 ) == ( bv_1_0_n53 )  ;
assign n8357 =  ( wr_addr ) == ( bv_8_22_n113 )  ;
assign n8358 =  ( n8356 ) & (n8357 )  ;
assign n8359 =  ( n8358 ) & (wr )  ;
assign n8360 =  ( n8359 ) ? ( n5096 ) : ( iram_22 ) ;
assign n8361 = wr_addr[7:7] ;
assign n8362 =  ( n8361 ) == ( bv_1_0_n53 )  ;
assign n8363 =  ( wr_addr ) == ( bv_8_22_n113 )  ;
assign n8364 =  ( n8362 ) & (n8363 )  ;
assign n8365 =  ( n8364 ) & (wr )  ;
assign n8366 =  ( n8365 ) ? ( n5123 ) : ( iram_22 ) ;
assign n8367 = wr_addr[7:7] ;
assign n8368 =  ( n8367 ) == ( bv_1_0_n53 )  ;
assign n8369 =  ( wr_addr ) == ( bv_8_22_n113 )  ;
assign n8370 =  ( n8368 ) & (n8369 )  ;
assign n8371 =  ( n8370 ) & (wr )  ;
assign n8372 =  ( n8371 ) ? ( n5165 ) : ( iram_22 ) ;
assign n8373 = wr_addr[7:7] ;
assign n8374 =  ( n8373 ) == ( bv_1_0_n53 )  ;
assign n8375 =  ( wr_addr ) == ( bv_8_22_n113 )  ;
assign n8376 =  ( n8374 ) & (n8375 )  ;
assign n8377 =  ( n8376 ) & (wr )  ;
assign n8378 =  ( n8377 ) ? ( n5204 ) : ( iram_22 ) ;
assign n8379 = wr_addr[7:7] ;
assign n8380 =  ( n8379 ) == ( bv_1_0_n53 )  ;
assign n8381 =  ( wr_addr ) == ( bv_8_22_n113 )  ;
assign n8382 =  ( n8380 ) & (n8381 )  ;
assign n8383 =  ( n8382 ) & (wr )  ;
assign n8384 =  ( n8383 ) ? ( n5262 ) : ( iram_22 ) ;
assign n8385 = wr_addr[7:7] ;
assign n8386 =  ( n8385 ) == ( bv_1_0_n53 )  ;
assign n8387 =  ( wr_addr ) == ( bv_8_22_n113 )  ;
assign n8388 =  ( n8386 ) & (n8387 )  ;
assign n8389 =  ( n8388 ) & (wr )  ;
assign n8390 =  ( n8389 ) ? ( n5298 ) : ( iram_22 ) ;
assign n8391 = wr_addr[7:7] ;
assign n8392 =  ( n8391 ) == ( bv_1_0_n53 )  ;
assign n8393 =  ( wr_addr ) == ( bv_8_22_n113 )  ;
assign n8394 =  ( n8392 ) & (n8393 )  ;
assign n8395 =  ( n8394 ) & (wr )  ;
assign n8396 =  ( n8395 ) ? ( n5325 ) : ( iram_22 ) ;
assign n8397 = wr_addr[7:7] ;
assign n8398 =  ( n8397 ) == ( bv_1_0_n53 )  ;
assign n8399 =  ( wr_addr ) == ( bv_8_23_n115 )  ;
assign n8400 =  ( n8398 ) & (n8399 )  ;
assign n8401 =  ( n8400 ) & (wr )  ;
assign n8402 =  ( n8401 ) ? ( n4782 ) : ( iram_23 ) ;
assign n8403 = wr_addr[7:7] ;
assign n8404 =  ( n8403 ) == ( bv_1_0_n53 )  ;
assign n8405 =  ( wr_addr ) == ( bv_8_23_n115 )  ;
assign n8406 =  ( n8404 ) & (n8405 )  ;
assign n8407 =  ( n8406 ) & (wr )  ;
assign n8408 =  ( n8407 ) ? ( n4841 ) : ( iram_23 ) ;
assign n8409 = wr_addr[7:7] ;
assign n8410 =  ( n8409 ) == ( bv_1_0_n53 )  ;
assign n8411 =  ( wr_addr ) == ( bv_8_23_n115 )  ;
assign n8412 =  ( n8410 ) & (n8411 )  ;
assign n8413 =  ( n8412 ) & (wr )  ;
assign n8414 =  ( n8413 ) ? ( n5449 ) : ( iram_23 ) ;
assign n8415 = wr_addr[7:7] ;
assign n8416 =  ( n8415 ) == ( bv_1_0_n53 )  ;
assign n8417 =  ( wr_addr ) == ( bv_8_23_n115 )  ;
assign n8418 =  ( n8416 ) & (n8417 )  ;
assign n8419 =  ( n8418 ) & (wr )  ;
assign n8420 =  ( n8419 ) ? ( n4906 ) : ( iram_23 ) ;
assign n8421 = wr_addr[7:7] ;
assign n8422 =  ( n8421 ) == ( bv_1_0_n53 )  ;
assign n8423 =  ( wr_addr ) == ( bv_8_23_n115 )  ;
assign n8424 =  ( n8422 ) & (n8423 )  ;
assign n8425 =  ( n8424 ) & (wr )  ;
assign n8426 =  ( n8425 ) ? ( n5485 ) : ( iram_23 ) ;
assign n8427 = wr_addr[7:7] ;
assign n8428 =  ( n8427 ) == ( bv_1_0_n53 )  ;
assign n8429 =  ( wr_addr ) == ( bv_8_23_n115 )  ;
assign n8430 =  ( n8428 ) & (n8429 )  ;
assign n8431 =  ( n8430 ) & (wr )  ;
assign n8432 =  ( n8431 ) ? ( n5512 ) : ( iram_23 ) ;
assign n8433 = wr_addr[7:7] ;
assign n8434 =  ( n8433 ) == ( bv_1_0_n53 )  ;
assign n8435 =  ( wr_addr ) == ( bv_8_23_n115 )  ;
assign n8436 =  ( n8434 ) & (n8435 )  ;
assign n8437 =  ( n8436 ) & (wr )  ;
assign n8438 =  ( n8437 ) ? ( bv_8_0_n69 ) : ( iram_23 ) ;
assign n8439 = wr_addr[7:7] ;
assign n8440 =  ( n8439 ) == ( bv_1_0_n53 )  ;
assign n8441 =  ( wr_addr ) == ( bv_8_23_n115 )  ;
assign n8442 =  ( n8440 ) & (n8441 )  ;
assign n8443 =  ( n8442 ) & (wr )  ;
assign n8444 =  ( n8443 ) ? ( n5071 ) : ( iram_23 ) ;
assign n8445 = wr_addr[7:7] ;
assign n8446 =  ( n8445 ) == ( bv_1_0_n53 )  ;
assign n8447 =  ( wr_addr ) == ( bv_8_23_n115 )  ;
assign n8448 =  ( n8446 ) & (n8447 )  ;
assign n8449 =  ( n8448 ) & (wr )  ;
assign n8450 =  ( n8449 ) ? ( n5096 ) : ( iram_23 ) ;
assign n8451 = wr_addr[7:7] ;
assign n8452 =  ( n8451 ) == ( bv_1_0_n53 )  ;
assign n8453 =  ( wr_addr ) == ( bv_8_23_n115 )  ;
assign n8454 =  ( n8452 ) & (n8453 )  ;
assign n8455 =  ( n8454 ) & (wr )  ;
assign n8456 =  ( n8455 ) ? ( n5123 ) : ( iram_23 ) ;
assign n8457 = wr_addr[7:7] ;
assign n8458 =  ( n8457 ) == ( bv_1_0_n53 )  ;
assign n8459 =  ( wr_addr ) == ( bv_8_23_n115 )  ;
assign n8460 =  ( n8458 ) & (n8459 )  ;
assign n8461 =  ( n8460 ) & (wr )  ;
assign n8462 =  ( n8461 ) ? ( n5165 ) : ( iram_23 ) ;
assign n8463 = wr_addr[7:7] ;
assign n8464 =  ( n8463 ) == ( bv_1_0_n53 )  ;
assign n8465 =  ( wr_addr ) == ( bv_8_23_n115 )  ;
assign n8466 =  ( n8464 ) & (n8465 )  ;
assign n8467 =  ( n8466 ) & (wr )  ;
assign n8468 =  ( n8467 ) ? ( n5204 ) : ( iram_23 ) ;
assign n8469 = wr_addr[7:7] ;
assign n8470 =  ( n8469 ) == ( bv_1_0_n53 )  ;
assign n8471 =  ( wr_addr ) == ( bv_8_23_n115 )  ;
assign n8472 =  ( n8470 ) & (n8471 )  ;
assign n8473 =  ( n8472 ) & (wr )  ;
assign n8474 =  ( n8473 ) ? ( n5262 ) : ( iram_23 ) ;
assign n8475 = wr_addr[7:7] ;
assign n8476 =  ( n8475 ) == ( bv_1_0_n53 )  ;
assign n8477 =  ( wr_addr ) == ( bv_8_23_n115 )  ;
assign n8478 =  ( n8476 ) & (n8477 )  ;
assign n8479 =  ( n8478 ) & (wr )  ;
assign n8480 =  ( n8479 ) ? ( n5298 ) : ( iram_23 ) ;
assign n8481 = wr_addr[7:7] ;
assign n8482 =  ( n8481 ) == ( bv_1_0_n53 )  ;
assign n8483 =  ( wr_addr ) == ( bv_8_23_n115 )  ;
assign n8484 =  ( n8482 ) & (n8483 )  ;
assign n8485 =  ( n8484 ) & (wr )  ;
assign n8486 =  ( n8485 ) ? ( n5325 ) : ( iram_23 ) ;
assign n8487 = wr_addr[7:7] ;
assign n8488 =  ( n8487 ) == ( bv_1_0_n53 )  ;
assign n8489 =  ( wr_addr ) == ( bv_8_24_n117 )  ;
assign n8490 =  ( n8488 ) & (n8489 )  ;
assign n8491 =  ( n8490 ) & (wr )  ;
assign n8492 =  ( n8491 ) ? ( n4782 ) : ( iram_24 ) ;
assign n8493 = wr_addr[7:7] ;
assign n8494 =  ( n8493 ) == ( bv_1_0_n53 )  ;
assign n8495 =  ( wr_addr ) == ( bv_8_24_n117 )  ;
assign n8496 =  ( n8494 ) & (n8495 )  ;
assign n8497 =  ( n8496 ) & (wr )  ;
assign n8498 =  ( n8497 ) ? ( n4841 ) : ( iram_24 ) ;
assign n8499 = wr_addr[7:7] ;
assign n8500 =  ( n8499 ) == ( bv_1_0_n53 )  ;
assign n8501 =  ( wr_addr ) == ( bv_8_24_n117 )  ;
assign n8502 =  ( n8500 ) & (n8501 )  ;
assign n8503 =  ( n8502 ) & (wr )  ;
assign n8504 =  ( n8503 ) ? ( n5449 ) : ( iram_24 ) ;
assign n8505 = wr_addr[7:7] ;
assign n8506 =  ( n8505 ) == ( bv_1_0_n53 )  ;
assign n8507 =  ( wr_addr ) == ( bv_8_24_n117 )  ;
assign n8508 =  ( n8506 ) & (n8507 )  ;
assign n8509 =  ( n8508 ) & (wr )  ;
assign n8510 =  ( n8509 ) ? ( n4906 ) : ( iram_24 ) ;
assign n8511 = wr_addr[7:7] ;
assign n8512 =  ( n8511 ) == ( bv_1_0_n53 )  ;
assign n8513 =  ( wr_addr ) == ( bv_8_24_n117 )  ;
assign n8514 =  ( n8512 ) & (n8513 )  ;
assign n8515 =  ( n8514 ) & (wr )  ;
assign n8516 =  ( n8515 ) ? ( n5485 ) : ( iram_24 ) ;
assign n8517 = wr_addr[7:7] ;
assign n8518 =  ( n8517 ) == ( bv_1_0_n53 )  ;
assign n8519 =  ( wr_addr ) == ( bv_8_24_n117 )  ;
assign n8520 =  ( n8518 ) & (n8519 )  ;
assign n8521 =  ( n8520 ) & (wr )  ;
assign n8522 =  ( n8521 ) ? ( n5512 ) : ( iram_24 ) ;
assign n8523 = wr_addr[7:7] ;
assign n8524 =  ( n8523 ) == ( bv_1_0_n53 )  ;
assign n8525 =  ( wr_addr ) == ( bv_8_24_n117 )  ;
assign n8526 =  ( n8524 ) & (n8525 )  ;
assign n8527 =  ( n8526 ) & (wr )  ;
assign n8528 =  ( n8527 ) ? ( bv_8_0_n69 ) : ( iram_24 ) ;
assign n8529 = wr_addr[7:7] ;
assign n8530 =  ( n8529 ) == ( bv_1_0_n53 )  ;
assign n8531 =  ( wr_addr ) == ( bv_8_24_n117 )  ;
assign n8532 =  ( n8530 ) & (n8531 )  ;
assign n8533 =  ( n8532 ) & (wr )  ;
assign n8534 =  ( n8533 ) ? ( n5071 ) : ( iram_24 ) ;
assign n8535 = wr_addr[7:7] ;
assign n8536 =  ( n8535 ) == ( bv_1_0_n53 )  ;
assign n8537 =  ( wr_addr ) == ( bv_8_24_n117 )  ;
assign n8538 =  ( n8536 ) & (n8537 )  ;
assign n8539 =  ( n8538 ) & (wr )  ;
assign n8540 =  ( n8539 ) ? ( n5096 ) : ( iram_24 ) ;
assign n8541 = wr_addr[7:7] ;
assign n8542 =  ( n8541 ) == ( bv_1_0_n53 )  ;
assign n8543 =  ( wr_addr ) == ( bv_8_24_n117 )  ;
assign n8544 =  ( n8542 ) & (n8543 )  ;
assign n8545 =  ( n8544 ) & (wr )  ;
assign n8546 =  ( n8545 ) ? ( n5123 ) : ( iram_24 ) ;
assign n8547 = wr_addr[7:7] ;
assign n8548 =  ( n8547 ) == ( bv_1_0_n53 )  ;
assign n8549 =  ( wr_addr ) == ( bv_8_24_n117 )  ;
assign n8550 =  ( n8548 ) & (n8549 )  ;
assign n8551 =  ( n8550 ) & (wr )  ;
assign n8552 =  ( n8551 ) ? ( n5165 ) : ( iram_24 ) ;
assign n8553 = wr_addr[7:7] ;
assign n8554 =  ( n8553 ) == ( bv_1_0_n53 )  ;
assign n8555 =  ( wr_addr ) == ( bv_8_24_n117 )  ;
assign n8556 =  ( n8554 ) & (n8555 )  ;
assign n8557 =  ( n8556 ) & (wr )  ;
assign n8558 =  ( n8557 ) ? ( n5204 ) : ( iram_24 ) ;
assign n8559 = wr_addr[7:7] ;
assign n8560 =  ( n8559 ) == ( bv_1_0_n53 )  ;
assign n8561 =  ( wr_addr ) == ( bv_8_24_n117 )  ;
assign n8562 =  ( n8560 ) & (n8561 )  ;
assign n8563 =  ( n8562 ) & (wr )  ;
assign n8564 =  ( n8563 ) ? ( n5262 ) : ( iram_24 ) ;
assign n8565 = wr_addr[7:7] ;
assign n8566 =  ( n8565 ) == ( bv_1_0_n53 )  ;
assign n8567 =  ( wr_addr ) == ( bv_8_24_n117 )  ;
assign n8568 =  ( n8566 ) & (n8567 )  ;
assign n8569 =  ( n8568 ) & (wr )  ;
assign n8570 =  ( n8569 ) ? ( n5298 ) : ( iram_24 ) ;
assign n8571 = wr_addr[7:7] ;
assign n8572 =  ( n8571 ) == ( bv_1_0_n53 )  ;
assign n8573 =  ( wr_addr ) == ( bv_8_24_n117 )  ;
assign n8574 =  ( n8572 ) & (n8573 )  ;
assign n8575 =  ( n8574 ) & (wr )  ;
assign n8576 =  ( n8575 ) ? ( n5325 ) : ( iram_24 ) ;
assign n8577 = wr_addr[7:7] ;
assign n8578 =  ( n8577 ) == ( bv_1_0_n53 )  ;
assign n8579 =  ( wr_addr ) == ( bv_8_25_n119 )  ;
assign n8580 =  ( n8578 ) & (n8579 )  ;
assign n8581 =  ( n8580 ) & (wr )  ;
assign n8582 =  ( n8581 ) ? ( n4782 ) : ( iram_25 ) ;
assign n8583 = wr_addr[7:7] ;
assign n8584 =  ( n8583 ) == ( bv_1_0_n53 )  ;
assign n8585 =  ( wr_addr ) == ( bv_8_25_n119 )  ;
assign n8586 =  ( n8584 ) & (n8585 )  ;
assign n8587 =  ( n8586 ) & (wr )  ;
assign n8588 =  ( n8587 ) ? ( n4841 ) : ( iram_25 ) ;
assign n8589 = wr_addr[7:7] ;
assign n8590 =  ( n8589 ) == ( bv_1_0_n53 )  ;
assign n8591 =  ( wr_addr ) == ( bv_8_25_n119 )  ;
assign n8592 =  ( n8590 ) & (n8591 )  ;
assign n8593 =  ( n8592 ) & (wr )  ;
assign n8594 =  ( n8593 ) ? ( n5449 ) : ( iram_25 ) ;
assign n8595 = wr_addr[7:7] ;
assign n8596 =  ( n8595 ) == ( bv_1_0_n53 )  ;
assign n8597 =  ( wr_addr ) == ( bv_8_25_n119 )  ;
assign n8598 =  ( n8596 ) & (n8597 )  ;
assign n8599 =  ( n8598 ) & (wr )  ;
assign n8600 =  ( n8599 ) ? ( n4906 ) : ( iram_25 ) ;
assign n8601 = wr_addr[7:7] ;
assign n8602 =  ( n8601 ) == ( bv_1_0_n53 )  ;
assign n8603 =  ( wr_addr ) == ( bv_8_25_n119 )  ;
assign n8604 =  ( n8602 ) & (n8603 )  ;
assign n8605 =  ( n8604 ) & (wr )  ;
assign n8606 =  ( n8605 ) ? ( n5485 ) : ( iram_25 ) ;
assign n8607 = wr_addr[7:7] ;
assign n8608 =  ( n8607 ) == ( bv_1_0_n53 )  ;
assign n8609 =  ( wr_addr ) == ( bv_8_25_n119 )  ;
assign n8610 =  ( n8608 ) & (n8609 )  ;
assign n8611 =  ( n8610 ) & (wr )  ;
assign n8612 =  ( n8611 ) ? ( n5512 ) : ( iram_25 ) ;
assign n8613 = wr_addr[7:7] ;
assign n8614 =  ( n8613 ) == ( bv_1_0_n53 )  ;
assign n8615 =  ( wr_addr ) == ( bv_8_25_n119 )  ;
assign n8616 =  ( n8614 ) & (n8615 )  ;
assign n8617 =  ( n8616 ) & (wr )  ;
assign n8618 =  ( n8617 ) ? ( bv_8_0_n69 ) : ( iram_25 ) ;
assign n8619 = wr_addr[7:7] ;
assign n8620 =  ( n8619 ) == ( bv_1_0_n53 )  ;
assign n8621 =  ( wr_addr ) == ( bv_8_25_n119 )  ;
assign n8622 =  ( n8620 ) & (n8621 )  ;
assign n8623 =  ( n8622 ) & (wr )  ;
assign n8624 =  ( n8623 ) ? ( n5071 ) : ( iram_25 ) ;
assign n8625 = wr_addr[7:7] ;
assign n8626 =  ( n8625 ) == ( bv_1_0_n53 )  ;
assign n8627 =  ( wr_addr ) == ( bv_8_25_n119 )  ;
assign n8628 =  ( n8626 ) & (n8627 )  ;
assign n8629 =  ( n8628 ) & (wr )  ;
assign n8630 =  ( n8629 ) ? ( n5096 ) : ( iram_25 ) ;
assign n8631 = wr_addr[7:7] ;
assign n8632 =  ( n8631 ) == ( bv_1_0_n53 )  ;
assign n8633 =  ( wr_addr ) == ( bv_8_25_n119 )  ;
assign n8634 =  ( n8632 ) & (n8633 )  ;
assign n8635 =  ( n8634 ) & (wr )  ;
assign n8636 =  ( n8635 ) ? ( n5123 ) : ( iram_25 ) ;
assign n8637 = wr_addr[7:7] ;
assign n8638 =  ( n8637 ) == ( bv_1_0_n53 )  ;
assign n8639 =  ( wr_addr ) == ( bv_8_25_n119 )  ;
assign n8640 =  ( n8638 ) & (n8639 )  ;
assign n8641 =  ( n8640 ) & (wr )  ;
assign n8642 =  ( n8641 ) ? ( n5165 ) : ( iram_25 ) ;
assign n8643 = wr_addr[7:7] ;
assign n8644 =  ( n8643 ) == ( bv_1_0_n53 )  ;
assign n8645 =  ( wr_addr ) == ( bv_8_25_n119 )  ;
assign n8646 =  ( n8644 ) & (n8645 )  ;
assign n8647 =  ( n8646 ) & (wr )  ;
assign n8648 =  ( n8647 ) ? ( n5204 ) : ( iram_25 ) ;
assign n8649 = wr_addr[7:7] ;
assign n8650 =  ( n8649 ) == ( bv_1_0_n53 )  ;
assign n8651 =  ( wr_addr ) == ( bv_8_25_n119 )  ;
assign n8652 =  ( n8650 ) & (n8651 )  ;
assign n8653 =  ( n8652 ) & (wr )  ;
assign n8654 =  ( n8653 ) ? ( n5262 ) : ( iram_25 ) ;
assign n8655 = wr_addr[7:7] ;
assign n8656 =  ( n8655 ) == ( bv_1_0_n53 )  ;
assign n8657 =  ( wr_addr ) == ( bv_8_25_n119 )  ;
assign n8658 =  ( n8656 ) & (n8657 )  ;
assign n8659 =  ( n8658 ) & (wr )  ;
assign n8660 =  ( n8659 ) ? ( n5298 ) : ( iram_25 ) ;
assign n8661 = wr_addr[7:7] ;
assign n8662 =  ( n8661 ) == ( bv_1_0_n53 )  ;
assign n8663 =  ( wr_addr ) == ( bv_8_25_n119 )  ;
assign n8664 =  ( n8662 ) & (n8663 )  ;
assign n8665 =  ( n8664 ) & (wr )  ;
assign n8666 =  ( n8665 ) ? ( n5325 ) : ( iram_25 ) ;
assign n8667 = wr_addr[7:7] ;
assign n8668 =  ( n8667 ) == ( bv_1_0_n53 )  ;
assign n8669 =  ( wr_addr ) == ( bv_8_26_n121 )  ;
assign n8670 =  ( n8668 ) & (n8669 )  ;
assign n8671 =  ( n8670 ) & (wr )  ;
assign n8672 =  ( n8671 ) ? ( n4782 ) : ( iram_26 ) ;
assign n8673 = wr_addr[7:7] ;
assign n8674 =  ( n8673 ) == ( bv_1_0_n53 )  ;
assign n8675 =  ( wr_addr ) == ( bv_8_26_n121 )  ;
assign n8676 =  ( n8674 ) & (n8675 )  ;
assign n8677 =  ( n8676 ) & (wr )  ;
assign n8678 =  ( n8677 ) ? ( n4841 ) : ( iram_26 ) ;
assign n8679 = wr_addr[7:7] ;
assign n8680 =  ( n8679 ) == ( bv_1_0_n53 )  ;
assign n8681 =  ( wr_addr ) == ( bv_8_26_n121 )  ;
assign n8682 =  ( n8680 ) & (n8681 )  ;
assign n8683 =  ( n8682 ) & (wr )  ;
assign n8684 =  ( n8683 ) ? ( n5449 ) : ( iram_26 ) ;
assign n8685 = wr_addr[7:7] ;
assign n8686 =  ( n8685 ) == ( bv_1_0_n53 )  ;
assign n8687 =  ( wr_addr ) == ( bv_8_26_n121 )  ;
assign n8688 =  ( n8686 ) & (n8687 )  ;
assign n8689 =  ( n8688 ) & (wr )  ;
assign n8690 =  ( n8689 ) ? ( n4906 ) : ( iram_26 ) ;
assign n8691 = wr_addr[7:7] ;
assign n8692 =  ( n8691 ) == ( bv_1_0_n53 )  ;
assign n8693 =  ( wr_addr ) == ( bv_8_26_n121 )  ;
assign n8694 =  ( n8692 ) & (n8693 )  ;
assign n8695 =  ( n8694 ) & (wr )  ;
assign n8696 =  ( n8695 ) ? ( n5485 ) : ( iram_26 ) ;
assign n8697 = wr_addr[7:7] ;
assign n8698 =  ( n8697 ) == ( bv_1_0_n53 )  ;
assign n8699 =  ( wr_addr ) == ( bv_8_26_n121 )  ;
assign n8700 =  ( n8698 ) & (n8699 )  ;
assign n8701 =  ( n8700 ) & (wr )  ;
assign n8702 =  ( n8701 ) ? ( n5512 ) : ( iram_26 ) ;
assign n8703 = wr_addr[7:7] ;
assign n8704 =  ( n8703 ) == ( bv_1_0_n53 )  ;
assign n8705 =  ( wr_addr ) == ( bv_8_26_n121 )  ;
assign n8706 =  ( n8704 ) & (n8705 )  ;
assign n8707 =  ( n8706 ) & (wr )  ;
assign n8708 =  ( n8707 ) ? ( bv_8_0_n69 ) : ( iram_26 ) ;
assign n8709 = wr_addr[7:7] ;
assign n8710 =  ( n8709 ) == ( bv_1_0_n53 )  ;
assign n8711 =  ( wr_addr ) == ( bv_8_26_n121 )  ;
assign n8712 =  ( n8710 ) & (n8711 )  ;
assign n8713 =  ( n8712 ) & (wr )  ;
assign n8714 =  ( n8713 ) ? ( n5071 ) : ( iram_26 ) ;
assign n8715 = wr_addr[7:7] ;
assign n8716 =  ( n8715 ) == ( bv_1_0_n53 )  ;
assign n8717 =  ( wr_addr ) == ( bv_8_26_n121 )  ;
assign n8718 =  ( n8716 ) & (n8717 )  ;
assign n8719 =  ( n8718 ) & (wr )  ;
assign n8720 =  ( n8719 ) ? ( n5096 ) : ( iram_26 ) ;
assign n8721 = wr_addr[7:7] ;
assign n8722 =  ( n8721 ) == ( bv_1_0_n53 )  ;
assign n8723 =  ( wr_addr ) == ( bv_8_26_n121 )  ;
assign n8724 =  ( n8722 ) & (n8723 )  ;
assign n8725 =  ( n8724 ) & (wr )  ;
assign n8726 =  ( n8725 ) ? ( n5123 ) : ( iram_26 ) ;
assign n8727 = wr_addr[7:7] ;
assign n8728 =  ( n8727 ) == ( bv_1_0_n53 )  ;
assign n8729 =  ( wr_addr ) == ( bv_8_26_n121 )  ;
assign n8730 =  ( n8728 ) & (n8729 )  ;
assign n8731 =  ( n8730 ) & (wr )  ;
assign n8732 =  ( n8731 ) ? ( n5165 ) : ( iram_26 ) ;
assign n8733 = wr_addr[7:7] ;
assign n8734 =  ( n8733 ) == ( bv_1_0_n53 )  ;
assign n8735 =  ( wr_addr ) == ( bv_8_26_n121 )  ;
assign n8736 =  ( n8734 ) & (n8735 )  ;
assign n8737 =  ( n8736 ) & (wr )  ;
assign n8738 =  ( n8737 ) ? ( n5204 ) : ( iram_26 ) ;
assign n8739 = wr_addr[7:7] ;
assign n8740 =  ( n8739 ) == ( bv_1_0_n53 )  ;
assign n8741 =  ( wr_addr ) == ( bv_8_26_n121 )  ;
assign n8742 =  ( n8740 ) & (n8741 )  ;
assign n8743 =  ( n8742 ) & (wr )  ;
assign n8744 =  ( n8743 ) ? ( n5262 ) : ( iram_26 ) ;
assign n8745 = wr_addr[7:7] ;
assign n8746 =  ( n8745 ) == ( bv_1_0_n53 )  ;
assign n8747 =  ( wr_addr ) == ( bv_8_26_n121 )  ;
assign n8748 =  ( n8746 ) & (n8747 )  ;
assign n8749 =  ( n8748 ) & (wr )  ;
assign n8750 =  ( n8749 ) ? ( n5298 ) : ( iram_26 ) ;
assign n8751 = wr_addr[7:7] ;
assign n8752 =  ( n8751 ) == ( bv_1_0_n53 )  ;
assign n8753 =  ( wr_addr ) == ( bv_8_26_n121 )  ;
assign n8754 =  ( n8752 ) & (n8753 )  ;
assign n8755 =  ( n8754 ) & (wr )  ;
assign n8756 =  ( n8755 ) ? ( n5325 ) : ( iram_26 ) ;
assign n8757 = wr_addr[7:7] ;
assign n8758 =  ( n8757 ) == ( bv_1_0_n53 )  ;
assign n8759 =  ( wr_addr ) == ( bv_8_27_n123 )  ;
assign n8760 =  ( n8758 ) & (n8759 )  ;
assign n8761 =  ( n8760 ) & (wr )  ;
assign n8762 =  ( n8761 ) ? ( n4782 ) : ( iram_27 ) ;
assign n8763 = wr_addr[7:7] ;
assign n8764 =  ( n8763 ) == ( bv_1_0_n53 )  ;
assign n8765 =  ( wr_addr ) == ( bv_8_27_n123 )  ;
assign n8766 =  ( n8764 ) & (n8765 )  ;
assign n8767 =  ( n8766 ) & (wr )  ;
assign n8768 =  ( n8767 ) ? ( n4841 ) : ( iram_27 ) ;
assign n8769 = wr_addr[7:7] ;
assign n8770 =  ( n8769 ) == ( bv_1_0_n53 )  ;
assign n8771 =  ( wr_addr ) == ( bv_8_27_n123 )  ;
assign n8772 =  ( n8770 ) & (n8771 )  ;
assign n8773 =  ( n8772 ) & (wr )  ;
assign n8774 =  ( n8773 ) ? ( n5449 ) : ( iram_27 ) ;
assign n8775 = wr_addr[7:7] ;
assign n8776 =  ( n8775 ) == ( bv_1_0_n53 )  ;
assign n8777 =  ( wr_addr ) == ( bv_8_27_n123 )  ;
assign n8778 =  ( n8776 ) & (n8777 )  ;
assign n8779 =  ( n8778 ) & (wr )  ;
assign n8780 =  ( n8779 ) ? ( n4906 ) : ( iram_27 ) ;
assign n8781 = wr_addr[7:7] ;
assign n8782 =  ( n8781 ) == ( bv_1_0_n53 )  ;
assign n8783 =  ( wr_addr ) == ( bv_8_27_n123 )  ;
assign n8784 =  ( n8782 ) & (n8783 )  ;
assign n8785 =  ( n8784 ) & (wr )  ;
assign n8786 =  ( n8785 ) ? ( n5485 ) : ( iram_27 ) ;
assign n8787 = wr_addr[7:7] ;
assign n8788 =  ( n8787 ) == ( bv_1_0_n53 )  ;
assign n8789 =  ( wr_addr ) == ( bv_8_27_n123 )  ;
assign n8790 =  ( n8788 ) & (n8789 )  ;
assign n8791 =  ( n8790 ) & (wr )  ;
assign n8792 =  ( n8791 ) ? ( n5512 ) : ( iram_27 ) ;
assign n8793 = wr_addr[7:7] ;
assign n8794 =  ( n8793 ) == ( bv_1_0_n53 )  ;
assign n8795 =  ( wr_addr ) == ( bv_8_27_n123 )  ;
assign n8796 =  ( n8794 ) & (n8795 )  ;
assign n8797 =  ( n8796 ) & (wr )  ;
assign n8798 =  ( n8797 ) ? ( bv_8_0_n69 ) : ( iram_27 ) ;
assign n8799 = wr_addr[7:7] ;
assign n8800 =  ( n8799 ) == ( bv_1_0_n53 )  ;
assign n8801 =  ( wr_addr ) == ( bv_8_27_n123 )  ;
assign n8802 =  ( n8800 ) & (n8801 )  ;
assign n8803 =  ( n8802 ) & (wr )  ;
assign n8804 =  ( n8803 ) ? ( n5071 ) : ( iram_27 ) ;
assign n8805 = wr_addr[7:7] ;
assign n8806 =  ( n8805 ) == ( bv_1_0_n53 )  ;
assign n8807 =  ( wr_addr ) == ( bv_8_27_n123 )  ;
assign n8808 =  ( n8806 ) & (n8807 )  ;
assign n8809 =  ( n8808 ) & (wr )  ;
assign n8810 =  ( n8809 ) ? ( n5096 ) : ( iram_27 ) ;
assign n8811 = wr_addr[7:7] ;
assign n8812 =  ( n8811 ) == ( bv_1_0_n53 )  ;
assign n8813 =  ( wr_addr ) == ( bv_8_27_n123 )  ;
assign n8814 =  ( n8812 ) & (n8813 )  ;
assign n8815 =  ( n8814 ) & (wr )  ;
assign n8816 =  ( n8815 ) ? ( n5123 ) : ( iram_27 ) ;
assign n8817 = wr_addr[7:7] ;
assign n8818 =  ( n8817 ) == ( bv_1_0_n53 )  ;
assign n8819 =  ( wr_addr ) == ( bv_8_27_n123 )  ;
assign n8820 =  ( n8818 ) & (n8819 )  ;
assign n8821 =  ( n8820 ) & (wr )  ;
assign n8822 =  ( n8821 ) ? ( n5165 ) : ( iram_27 ) ;
assign n8823 = wr_addr[7:7] ;
assign n8824 =  ( n8823 ) == ( bv_1_0_n53 )  ;
assign n8825 =  ( wr_addr ) == ( bv_8_27_n123 )  ;
assign n8826 =  ( n8824 ) & (n8825 )  ;
assign n8827 =  ( n8826 ) & (wr )  ;
assign n8828 =  ( n8827 ) ? ( n5204 ) : ( iram_27 ) ;
assign n8829 = wr_addr[7:7] ;
assign n8830 =  ( n8829 ) == ( bv_1_0_n53 )  ;
assign n8831 =  ( wr_addr ) == ( bv_8_27_n123 )  ;
assign n8832 =  ( n8830 ) & (n8831 )  ;
assign n8833 =  ( n8832 ) & (wr )  ;
assign n8834 =  ( n8833 ) ? ( n5262 ) : ( iram_27 ) ;
assign n8835 = wr_addr[7:7] ;
assign n8836 =  ( n8835 ) == ( bv_1_0_n53 )  ;
assign n8837 =  ( wr_addr ) == ( bv_8_27_n123 )  ;
assign n8838 =  ( n8836 ) & (n8837 )  ;
assign n8839 =  ( n8838 ) & (wr )  ;
assign n8840 =  ( n8839 ) ? ( n5298 ) : ( iram_27 ) ;
assign n8841 = wr_addr[7:7] ;
assign n8842 =  ( n8841 ) == ( bv_1_0_n53 )  ;
assign n8843 =  ( wr_addr ) == ( bv_8_27_n123 )  ;
assign n8844 =  ( n8842 ) & (n8843 )  ;
assign n8845 =  ( n8844 ) & (wr )  ;
assign n8846 =  ( n8845 ) ? ( n5325 ) : ( iram_27 ) ;
assign n8847 = wr_addr[7:7] ;
assign n8848 =  ( n8847 ) == ( bv_1_0_n53 )  ;
assign n8849 =  ( wr_addr ) == ( bv_8_28_n125 )  ;
assign n8850 =  ( n8848 ) & (n8849 )  ;
assign n8851 =  ( n8850 ) & (wr )  ;
assign n8852 =  ( n8851 ) ? ( n4782 ) : ( iram_28 ) ;
assign n8853 = wr_addr[7:7] ;
assign n8854 =  ( n8853 ) == ( bv_1_0_n53 )  ;
assign n8855 =  ( wr_addr ) == ( bv_8_28_n125 )  ;
assign n8856 =  ( n8854 ) & (n8855 )  ;
assign n8857 =  ( n8856 ) & (wr )  ;
assign n8858 =  ( n8857 ) ? ( n4841 ) : ( iram_28 ) ;
assign n8859 = wr_addr[7:7] ;
assign n8860 =  ( n8859 ) == ( bv_1_0_n53 )  ;
assign n8861 =  ( wr_addr ) == ( bv_8_28_n125 )  ;
assign n8862 =  ( n8860 ) & (n8861 )  ;
assign n8863 =  ( n8862 ) & (wr )  ;
assign n8864 =  ( n8863 ) ? ( n5449 ) : ( iram_28 ) ;
assign n8865 = wr_addr[7:7] ;
assign n8866 =  ( n8865 ) == ( bv_1_0_n53 )  ;
assign n8867 =  ( wr_addr ) == ( bv_8_28_n125 )  ;
assign n8868 =  ( n8866 ) & (n8867 )  ;
assign n8869 =  ( n8868 ) & (wr )  ;
assign n8870 =  ( n8869 ) ? ( n4906 ) : ( iram_28 ) ;
assign n8871 = wr_addr[7:7] ;
assign n8872 =  ( n8871 ) == ( bv_1_0_n53 )  ;
assign n8873 =  ( wr_addr ) == ( bv_8_28_n125 )  ;
assign n8874 =  ( n8872 ) & (n8873 )  ;
assign n8875 =  ( n8874 ) & (wr )  ;
assign n8876 =  ( n8875 ) ? ( n5485 ) : ( iram_28 ) ;
assign n8877 = wr_addr[7:7] ;
assign n8878 =  ( n8877 ) == ( bv_1_0_n53 )  ;
assign n8879 =  ( wr_addr ) == ( bv_8_28_n125 )  ;
assign n8880 =  ( n8878 ) & (n8879 )  ;
assign n8881 =  ( n8880 ) & (wr )  ;
assign n8882 =  ( n8881 ) ? ( n5512 ) : ( iram_28 ) ;
assign n8883 = wr_addr[7:7] ;
assign n8884 =  ( n8883 ) == ( bv_1_0_n53 )  ;
assign n8885 =  ( wr_addr ) == ( bv_8_28_n125 )  ;
assign n8886 =  ( n8884 ) & (n8885 )  ;
assign n8887 =  ( n8886 ) & (wr )  ;
assign n8888 =  ( n8887 ) ? ( bv_8_0_n69 ) : ( iram_28 ) ;
assign n8889 = wr_addr[7:7] ;
assign n8890 =  ( n8889 ) == ( bv_1_0_n53 )  ;
assign n8891 =  ( wr_addr ) == ( bv_8_28_n125 )  ;
assign n8892 =  ( n8890 ) & (n8891 )  ;
assign n8893 =  ( n8892 ) & (wr )  ;
assign n8894 =  ( n8893 ) ? ( n5071 ) : ( iram_28 ) ;
assign n8895 = wr_addr[7:7] ;
assign n8896 =  ( n8895 ) == ( bv_1_0_n53 )  ;
assign n8897 =  ( wr_addr ) == ( bv_8_28_n125 )  ;
assign n8898 =  ( n8896 ) & (n8897 )  ;
assign n8899 =  ( n8898 ) & (wr )  ;
assign n8900 =  ( n8899 ) ? ( n5096 ) : ( iram_28 ) ;
assign n8901 = wr_addr[7:7] ;
assign n8902 =  ( n8901 ) == ( bv_1_0_n53 )  ;
assign n8903 =  ( wr_addr ) == ( bv_8_28_n125 )  ;
assign n8904 =  ( n8902 ) & (n8903 )  ;
assign n8905 =  ( n8904 ) & (wr )  ;
assign n8906 =  ( n8905 ) ? ( n5123 ) : ( iram_28 ) ;
assign n8907 = wr_addr[7:7] ;
assign n8908 =  ( n8907 ) == ( bv_1_0_n53 )  ;
assign n8909 =  ( wr_addr ) == ( bv_8_28_n125 )  ;
assign n8910 =  ( n8908 ) & (n8909 )  ;
assign n8911 =  ( n8910 ) & (wr )  ;
assign n8912 =  ( n8911 ) ? ( n5165 ) : ( iram_28 ) ;
assign n8913 = wr_addr[7:7] ;
assign n8914 =  ( n8913 ) == ( bv_1_0_n53 )  ;
assign n8915 =  ( wr_addr ) == ( bv_8_28_n125 )  ;
assign n8916 =  ( n8914 ) & (n8915 )  ;
assign n8917 =  ( n8916 ) & (wr )  ;
assign n8918 =  ( n8917 ) ? ( n5204 ) : ( iram_28 ) ;
assign n8919 = wr_addr[7:7] ;
assign n8920 =  ( n8919 ) == ( bv_1_0_n53 )  ;
assign n8921 =  ( wr_addr ) == ( bv_8_28_n125 )  ;
assign n8922 =  ( n8920 ) & (n8921 )  ;
assign n8923 =  ( n8922 ) & (wr )  ;
assign n8924 =  ( n8923 ) ? ( n5262 ) : ( iram_28 ) ;
assign n8925 = wr_addr[7:7] ;
assign n8926 =  ( n8925 ) == ( bv_1_0_n53 )  ;
assign n8927 =  ( wr_addr ) == ( bv_8_28_n125 )  ;
assign n8928 =  ( n8926 ) & (n8927 )  ;
assign n8929 =  ( n8928 ) & (wr )  ;
assign n8930 =  ( n8929 ) ? ( n5298 ) : ( iram_28 ) ;
assign n8931 = wr_addr[7:7] ;
assign n8932 =  ( n8931 ) == ( bv_1_0_n53 )  ;
assign n8933 =  ( wr_addr ) == ( bv_8_28_n125 )  ;
assign n8934 =  ( n8932 ) & (n8933 )  ;
assign n8935 =  ( n8934 ) & (wr )  ;
assign n8936 =  ( n8935 ) ? ( n5325 ) : ( iram_28 ) ;
assign n8937 = wr_addr[7:7] ;
assign n8938 =  ( n8937 ) == ( bv_1_0_n53 )  ;
assign n8939 =  ( wr_addr ) == ( bv_8_29_n127 )  ;
assign n8940 =  ( n8938 ) & (n8939 )  ;
assign n8941 =  ( n8940 ) & (wr )  ;
assign n8942 =  ( n8941 ) ? ( n4782 ) : ( iram_29 ) ;
assign n8943 = wr_addr[7:7] ;
assign n8944 =  ( n8943 ) == ( bv_1_0_n53 )  ;
assign n8945 =  ( wr_addr ) == ( bv_8_29_n127 )  ;
assign n8946 =  ( n8944 ) & (n8945 )  ;
assign n8947 =  ( n8946 ) & (wr )  ;
assign n8948 =  ( n8947 ) ? ( n4841 ) : ( iram_29 ) ;
assign n8949 = wr_addr[7:7] ;
assign n8950 =  ( n8949 ) == ( bv_1_0_n53 )  ;
assign n8951 =  ( wr_addr ) == ( bv_8_29_n127 )  ;
assign n8952 =  ( n8950 ) & (n8951 )  ;
assign n8953 =  ( n8952 ) & (wr )  ;
assign n8954 =  ( n8953 ) ? ( n5449 ) : ( iram_29 ) ;
assign n8955 = wr_addr[7:7] ;
assign n8956 =  ( n8955 ) == ( bv_1_0_n53 )  ;
assign n8957 =  ( wr_addr ) == ( bv_8_29_n127 )  ;
assign n8958 =  ( n8956 ) & (n8957 )  ;
assign n8959 =  ( n8958 ) & (wr )  ;
assign n8960 =  ( n8959 ) ? ( n4906 ) : ( iram_29 ) ;
assign n8961 = wr_addr[7:7] ;
assign n8962 =  ( n8961 ) == ( bv_1_0_n53 )  ;
assign n8963 =  ( wr_addr ) == ( bv_8_29_n127 )  ;
assign n8964 =  ( n8962 ) & (n8963 )  ;
assign n8965 =  ( n8964 ) & (wr )  ;
assign n8966 =  ( n8965 ) ? ( n5485 ) : ( iram_29 ) ;
assign n8967 = wr_addr[7:7] ;
assign n8968 =  ( n8967 ) == ( bv_1_0_n53 )  ;
assign n8969 =  ( wr_addr ) == ( bv_8_29_n127 )  ;
assign n8970 =  ( n8968 ) & (n8969 )  ;
assign n8971 =  ( n8970 ) & (wr )  ;
assign n8972 =  ( n8971 ) ? ( n5512 ) : ( iram_29 ) ;
assign n8973 = wr_addr[7:7] ;
assign n8974 =  ( n8973 ) == ( bv_1_0_n53 )  ;
assign n8975 =  ( wr_addr ) == ( bv_8_29_n127 )  ;
assign n8976 =  ( n8974 ) & (n8975 )  ;
assign n8977 =  ( n8976 ) & (wr )  ;
assign n8978 =  ( n8977 ) ? ( bv_8_0_n69 ) : ( iram_29 ) ;
assign n8979 = wr_addr[7:7] ;
assign n8980 =  ( n8979 ) == ( bv_1_0_n53 )  ;
assign n8981 =  ( wr_addr ) == ( bv_8_29_n127 )  ;
assign n8982 =  ( n8980 ) & (n8981 )  ;
assign n8983 =  ( n8982 ) & (wr )  ;
assign n8984 =  ( n8983 ) ? ( n5071 ) : ( iram_29 ) ;
assign n8985 = wr_addr[7:7] ;
assign n8986 =  ( n8985 ) == ( bv_1_0_n53 )  ;
assign n8987 =  ( wr_addr ) == ( bv_8_29_n127 )  ;
assign n8988 =  ( n8986 ) & (n8987 )  ;
assign n8989 =  ( n8988 ) & (wr )  ;
assign n8990 =  ( n8989 ) ? ( n5096 ) : ( iram_29 ) ;
assign n8991 = wr_addr[7:7] ;
assign n8992 =  ( n8991 ) == ( bv_1_0_n53 )  ;
assign n8993 =  ( wr_addr ) == ( bv_8_29_n127 )  ;
assign n8994 =  ( n8992 ) & (n8993 )  ;
assign n8995 =  ( n8994 ) & (wr )  ;
assign n8996 =  ( n8995 ) ? ( n5123 ) : ( iram_29 ) ;
assign n8997 = wr_addr[7:7] ;
assign n8998 =  ( n8997 ) == ( bv_1_0_n53 )  ;
assign n8999 =  ( wr_addr ) == ( bv_8_29_n127 )  ;
assign n9000 =  ( n8998 ) & (n8999 )  ;
assign n9001 =  ( n9000 ) & (wr )  ;
assign n9002 =  ( n9001 ) ? ( n5165 ) : ( iram_29 ) ;
assign n9003 = wr_addr[7:7] ;
assign n9004 =  ( n9003 ) == ( bv_1_0_n53 )  ;
assign n9005 =  ( wr_addr ) == ( bv_8_29_n127 )  ;
assign n9006 =  ( n9004 ) & (n9005 )  ;
assign n9007 =  ( n9006 ) & (wr )  ;
assign n9008 =  ( n9007 ) ? ( n5204 ) : ( iram_29 ) ;
assign n9009 = wr_addr[7:7] ;
assign n9010 =  ( n9009 ) == ( bv_1_0_n53 )  ;
assign n9011 =  ( wr_addr ) == ( bv_8_29_n127 )  ;
assign n9012 =  ( n9010 ) & (n9011 )  ;
assign n9013 =  ( n9012 ) & (wr )  ;
assign n9014 =  ( n9013 ) ? ( n5262 ) : ( iram_29 ) ;
assign n9015 = wr_addr[7:7] ;
assign n9016 =  ( n9015 ) == ( bv_1_0_n53 )  ;
assign n9017 =  ( wr_addr ) == ( bv_8_29_n127 )  ;
assign n9018 =  ( n9016 ) & (n9017 )  ;
assign n9019 =  ( n9018 ) & (wr )  ;
assign n9020 =  ( n9019 ) ? ( n5298 ) : ( iram_29 ) ;
assign n9021 = wr_addr[7:7] ;
assign n9022 =  ( n9021 ) == ( bv_1_0_n53 )  ;
assign n9023 =  ( wr_addr ) == ( bv_8_29_n127 )  ;
assign n9024 =  ( n9022 ) & (n9023 )  ;
assign n9025 =  ( n9024 ) & (wr )  ;
assign n9026 =  ( n9025 ) ? ( n5325 ) : ( iram_29 ) ;
assign n9027 = wr_addr[7:7] ;
assign n9028 =  ( n9027 ) == ( bv_1_0_n53 )  ;
assign n9029 =  ( wr_addr ) == ( bv_8_30_n129 )  ;
assign n9030 =  ( n9028 ) & (n9029 )  ;
assign n9031 =  ( n9030 ) & (wr )  ;
assign n9032 =  ( n9031 ) ? ( n4782 ) : ( iram_30 ) ;
assign n9033 = wr_addr[7:7] ;
assign n9034 =  ( n9033 ) == ( bv_1_0_n53 )  ;
assign n9035 =  ( wr_addr ) == ( bv_8_30_n129 )  ;
assign n9036 =  ( n9034 ) & (n9035 )  ;
assign n9037 =  ( n9036 ) & (wr )  ;
assign n9038 =  ( n9037 ) ? ( n4841 ) : ( iram_30 ) ;
assign n9039 = wr_addr[7:7] ;
assign n9040 =  ( n9039 ) == ( bv_1_0_n53 )  ;
assign n9041 =  ( wr_addr ) == ( bv_8_30_n129 )  ;
assign n9042 =  ( n9040 ) & (n9041 )  ;
assign n9043 =  ( n9042 ) & (wr )  ;
assign n9044 =  ( n9043 ) ? ( n5449 ) : ( iram_30 ) ;
assign n9045 = wr_addr[7:7] ;
assign n9046 =  ( n9045 ) == ( bv_1_0_n53 )  ;
assign n9047 =  ( wr_addr ) == ( bv_8_30_n129 )  ;
assign n9048 =  ( n9046 ) & (n9047 )  ;
assign n9049 =  ( n9048 ) & (wr )  ;
assign n9050 =  ( n9049 ) ? ( n4906 ) : ( iram_30 ) ;
assign n9051 = wr_addr[7:7] ;
assign n9052 =  ( n9051 ) == ( bv_1_0_n53 )  ;
assign n9053 =  ( wr_addr ) == ( bv_8_30_n129 )  ;
assign n9054 =  ( n9052 ) & (n9053 )  ;
assign n9055 =  ( n9054 ) & (wr )  ;
assign n9056 =  ( n9055 ) ? ( n5485 ) : ( iram_30 ) ;
assign n9057 = wr_addr[7:7] ;
assign n9058 =  ( n9057 ) == ( bv_1_0_n53 )  ;
assign n9059 =  ( wr_addr ) == ( bv_8_30_n129 )  ;
assign n9060 =  ( n9058 ) & (n9059 )  ;
assign n9061 =  ( n9060 ) & (wr )  ;
assign n9062 =  ( n9061 ) ? ( n5512 ) : ( iram_30 ) ;
assign n9063 = wr_addr[7:7] ;
assign n9064 =  ( n9063 ) == ( bv_1_0_n53 )  ;
assign n9065 =  ( wr_addr ) == ( bv_8_30_n129 )  ;
assign n9066 =  ( n9064 ) & (n9065 )  ;
assign n9067 =  ( n9066 ) & (wr )  ;
assign n9068 =  ( n9067 ) ? ( bv_8_0_n69 ) : ( iram_30 ) ;
assign n9069 = wr_addr[7:7] ;
assign n9070 =  ( n9069 ) == ( bv_1_0_n53 )  ;
assign n9071 =  ( wr_addr ) == ( bv_8_30_n129 )  ;
assign n9072 =  ( n9070 ) & (n9071 )  ;
assign n9073 =  ( n9072 ) & (wr )  ;
assign n9074 =  ( n9073 ) ? ( n5071 ) : ( iram_30 ) ;
assign n9075 = wr_addr[7:7] ;
assign n9076 =  ( n9075 ) == ( bv_1_0_n53 )  ;
assign n9077 =  ( wr_addr ) == ( bv_8_30_n129 )  ;
assign n9078 =  ( n9076 ) & (n9077 )  ;
assign n9079 =  ( n9078 ) & (wr )  ;
assign n9080 =  ( n9079 ) ? ( n5096 ) : ( iram_30 ) ;
assign n9081 = wr_addr[7:7] ;
assign n9082 =  ( n9081 ) == ( bv_1_0_n53 )  ;
assign n9083 =  ( wr_addr ) == ( bv_8_30_n129 )  ;
assign n9084 =  ( n9082 ) & (n9083 )  ;
assign n9085 =  ( n9084 ) & (wr )  ;
assign n9086 =  ( n9085 ) ? ( n5123 ) : ( iram_30 ) ;
assign n9087 = wr_addr[7:7] ;
assign n9088 =  ( n9087 ) == ( bv_1_0_n53 )  ;
assign n9089 =  ( wr_addr ) == ( bv_8_30_n129 )  ;
assign n9090 =  ( n9088 ) & (n9089 )  ;
assign n9091 =  ( n9090 ) & (wr )  ;
assign n9092 =  ( n9091 ) ? ( n5165 ) : ( iram_30 ) ;
assign n9093 = wr_addr[7:7] ;
assign n9094 =  ( n9093 ) == ( bv_1_0_n53 )  ;
assign n9095 =  ( wr_addr ) == ( bv_8_30_n129 )  ;
assign n9096 =  ( n9094 ) & (n9095 )  ;
assign n9097 =  ( n9096 ) & (wr )  ;
assign n9098 =  ( n9097 ) ? ( n5204 ) : ( iram_30 ) ;
assign n9099 = wr_addr[7:7] ;
assign n9100 =  ( n9099 ) == ( bv_1_0_n53 )  ;
assign n9101 =  ( wr_addr ) == ( bv_8_30_n129 )  ;
assign n9102 =  ( n9100 ) & (n9101 )  ;
assign n9103 =  ( n9102 ) & (wr )  ;
assign n9104 =  ( n9103 ) ? ( n5262 ) : ( iram_30 ) ;
assign n9105 = wr_addr[7:7] ;
assign n9106 =  ( n9105 ) == ( bv_1_0_n53 )  ;
assign n9107 =  ( wr_addr ) == ( bv_8_30_n129 )  ;
assign n9108 =  ( n9106 ) & (n9107 )  ;
assign n9109 =  ( n9108 ) & (wr )  ;
assign n9110 =  ( n9109 ) ? ( n5298 ) : ( iram_30 ) ;
assign n9111 = wr_addr[7:7] ;
assign n9112 =  ( n9111 ) == ( bv_1_0_n53 )  ;
assign n9113 =  ( wr_addr ) == ( bv_8_30_n129 )  ;
assign n9114 =  ( n9112 ) & (n9113 )  ;
assign n9115 =  ( n9114 ) & (wr )  ;
assign n9116 =  ( n9115 ) ? ( n5325 ) : ( iram_30 ) ;
assign n9117 = wr_addr[7:7] ;
assign n9118 =  ( n9117 ) == ( bv_1_0_n53 )  ;
assign n9119 =  ( wr_addr ) == ( bv_8_31_n131 )  ;
assign n9120 =  ( n9118 ) & (n9119 )  ;
assign n9121 =  ( n9120 ) & (wr )  ;
assign n9122 =  ( n9121 ) ? ( n4782 ) : ( iram_31 ) ;
assign n9123 = wr_addr[7:7] ;
assign n9124 =  ( n9123 ) == ( bv_1_0_n53 )  ;
assign n9125 =  ( wr_addr ) == ( bv_8_31_n131 )  ;
assign n9126 =  ( n9124 ) & (n9125 )  ;
assign n9127 =  ( n9126 ) & (wr )  ;
assign n9128 =  ( n9127 ) ? ( n4841 ) : ( iram_31 ) ;
assign n9129 = wr_addr[7:7] ;
assign n9130 =  ( n9129 ) == ( bv_1_0_n53 )  ;
assign n9131 =  ( wr_addr ) == ( bv_8_31_n131 )  ;
assign n9132 =  ( n9130 ) & (n9131 )  ;
assign n9133 =  ( n9132 ) & (wr )  ;
assign n9134 =  ( n9133 ) ? ( n5449 ) : ( iram_31 ) ;
assign n9135 = wr_addr[7:7] ;
assign n9136 =  ( n9135 ) == ( bv_1_0_n53 )  ;
assign n9137 =  ( wr_addr ) == ( bv_8_31_n131 )  ;
assign n9138 =  ( n9136 ) & (n9137 )  ;
assign n9139 =  ( n9138 ) & (wr )  ;
assign n9140 =  ( n9139 ) ? ( n4906 ) : ( iram_31 ) ;
assign n9141 = wr_addr[7:7] ;
assign n9142 =  ( n9141 ) == ( bv_1_0_n53 )  ;
assign n9143 =  ( wr_addr ) == ( bv_8_31_n131 )  ;
assign n9144 =  ( n9142 ) & (n9143 )  ;
assign n9145 =  ( n9144 ) & (wr )  ;
assign n9146 =  ( n9145 ) ? ( n5485 ) : ( iram_31 ) ;
assign n9147 = wr_addr[7:7] ;
assign n9148 =  ( n9147 ) == ( bv_1_0_n53 )  ;
assign n9149 =  ( wr_addr ) == ( bv_8_31_n131 )  ;
assign n9150 =  ( n9148 ) & (n9149 )  ;
assign n9151 =  ( n9150 ) & (wr )  ;
assign n9152 =  ( n9151 ) ? ( n5512 ) : ( iram_31 ) ;
assign n9153 = wr_addr[7:7] ;
assign n9154 =  ( n9153 ) == ( bv_1_0_n53 )  ;
assign n9155 =  ( wr_addr ) == ( bv_8_31_n131 )  ;
assign n9156 =  ( n9154 ) & (n9155 )  ;
assign n9157 =  ( n9156 ) & (wr )  ;
assign n9158 =  ( n9157 ) ? ( bv_8_0_n69 ) : ( iram_31 ) ;
assign n9159 = wr_addr[7:7] ;
assign n9160 =  ( n9159 ) == ( bv_1_0_n53 )  ;
assign n9161 =  ( wr_addr ) == ( bv_8_31_n131 )  ;
assign n9162 =  ( n9160 ) & (n9161 )  ;
assign n9163 =  ( n9162 ) & (wr )  ;
assign n9164 =  ( n9163 ) ? ( n5071 ) : ( iram_31 ) ;
assign n9165 = wr_addr[7:7] ;
assign n9166 =  ( n9165 ) == ( bv_1_0_n53 )  ;
assign n9167 =  ( wr_addr ) == ( bv_8_31_n131 )  ;
assign n9168 =  ( n9166 ) & (n9167 )  ;
assign n9169 =  ( n9168 ) & (wr )  ;
assign n9170 =  ( n9169 ) ? ( n5096 ) : ( iram_31 ) ;
assign n9171 = wr_addr[7:7] ;
assign n9172 =  ( n9171 ) == ( bv_1_0_n53 )  ;
assign n9173 =  ( wr_addr ) == ( bv_8_31_n131 )  ;
assign n9174 =  ( n9172 ) & (n9173 )  ;
assign n9175 =  ( n9174 ) & (wr )  ;
assign n9176 =  ( n9175 ) ? ( n5123 ) : ( iram_31 ) ;
assign n9177 = wr_addr[7:7] ;
assign n9178 =  ( n9177 ) == ( bv_1_0_n53 )  ;
assign n9179 =  ( wr_addr ) == ( bv_8_31_n131 )  ;
assign n9180 =  ( n9178 ) & (n9179 )  ;
assign n9181 =  ( n9180 ) & (wr )  ;
assign n9182 =  ( n9181 ) ? ( n5165 ) : ( iram_31 ) ;
assign n9183 = wr_addr[7:7] ;
assign n9184 =  ( n9183 ) == ( bv_1_0_n53 )  ;
assign n9185 =  ( wr_addr ) == ( bv_8_31_n131 )  ;
assign n9186 =  ( n9184 ) & (n9185 )  ;
assign n9187 =  ( n9186 ) & (wr )  ;
assign n9188 =  ( n9187 ) ? ( n5204 ) : ( iram_31 ) ;
assign n9189 = wr_addr[7:7] ;
assign n9190 =  ( n9189 ) == ( bv_1_0_n53 )  ;
assign n9191 =  ( wr_addr ) == ( bv_8_31_n131 )  ;
assign n9192 =  ( n9190 ) & (n9191 )  ;
assign n9193 =  ( n9192 ) & (wr )  ;
assign n9194 =  ( n9193 ) ? ( n5262 ) : ( iram_31 ) ;
assign n9195 = wr_addr[7:7] ;
assign n9196 =  ( n9195 ) == ( bv_1_0_n53 )  ;
assign n9197 =  ( wr_addr ) == ( bv_8_31_n131 )  ;
assign n9198 =  ( n9196 ) & (n9197 )  ;
assign n9199 =  ( n9198 ) & (wr )  ;
assign n9200 =  ( n9199 ) ? ( n5298 ) : ( iram_31 ) ;
assign n9201 = wr_addr[7:7] ;
assign n9202 =  ( n9201 ) == ( bv_1_0_n53 )  ;
assign n9203 =  ( wr_addr ) == ( bv_8_31_n131 )  ;
assign n9204 =  ( n9202 ) & (n9203 )  ;
assign n9205 =  ( n9204 ) & (wr )  ;
assign n9206 =  ( n9205 ) ? ( n5325 ) : ( iram_31 ) ;
assign n9207 = wr_addr[7:7] ;
assign n9208 =  ( n9207 ) == ( bv_1_0_n53 )  ;
assign n9209 =  ( wr_addr ) == ( bv_8_32_n133 )  ;
assign n9210 =  ( n9208 ) & (n9209 )  ;
assign n9211 =  ( n9210 ) & (wr )  ;
assign n9212 =  ( n9211 ) ? ( n4782 ) : ( iram_32 ) ;
assign n9213 = wr_addr[7:7] ;
assign n9214 =  ( n9213 ) == ( bv_1_0_n53 )  ;
assign n9215 =  ( wr_addr ) == ( bv_8_32_n133 )  ;
assign n9216 =  ( n9214 ) & (n9215 )  ;
assign n9217 =  ( n9216 ) & (wr )  ;
assign n9218 =  ( n9217 ) ? ( n4841 ) : ( iram_32 ) ;
assign n9219 = wr_addr[7:7] ;
assign n9220 =  ( n9219 ) == ( bv_1_0_n53 )  ;
assign n9221 =  ( wr_addr ) == ( bv_8_32_n133 )  ;
assign n9222 =  ( n9220 ) & (n9221 )  ;
assign n9223 =  ( n9222 ) & (wr )  ;
assign n9224 =  ( n9223 ) ? ( n5449 ) : ( iram_32 ) ;
assign n9225 = wr_addr[7:7] ;
assign n9226 =  ( n9225 ) == ( bv_1_0_n53 )  ;
assign n9227 =  ( wr_addr ) == ( bv_8_32_n133 )  ;
assign n9228 =  ( n9226 ) & (n9227 )  ;
assign n9229 =  ( n9228 ) & (wr )  ;
assign n9230 =  ( n9229 ) ? ( n4906 ) : ( iram_32 ) ;
assign n9231 = wr_addr[7:7] ;
assign n9232 =  ( n9231 ) == ( bv_1_0_n53 )  ;
assign n9233 =  ( wr_addr ) == ( bv_8_32_n133 )  ;
assign n9234 =  ( n9232 ) & (n9233 )  ;
assign n9235 =  ( n9234 ) & (wr )  ;
assign n9236 =  ( n9235 ) ? ( n5485 ) : ( iram_32 ) ;
assign n9237 = wr_addr[7:7] ;
assign n9238 =  ( n9237 ) == ( bv_1_0_n53 )  ;
assign n9239 =  ( wr_addr ) == ( bv_8_32_n133 )  ;
assign n9240 =  ( n9238 ) & (n9239 )  ;
assign n9241 =  ( n9240 ) & (wr )  ;
assign n9242 =  ( n9241 ) ? ( n5512 ) : ( iram_32 ) ;
assign n9243 = wr_addr[7:7] ;
assign n9244 =  ( n9243 ) == ( bv_1_0_n53 )  ;
assign n9245 =  ( wr_addr ) == ( bv_8_32_n133 )  ;
assign n9246 =  ( n9244 ) & (n9245 )  ;
assign n9247 =  ( n9246 ) & (wr )  ;
assign n9248 =  ( n9247 ) ? ( bv_8_0_n69 ) : ( iram_32 ) ;
assign n9249 = wr_addr[7:7] ;
assign n9250 =  ( n9249 ) == ( bv_1_0_n53 )  ;
assign n9251 =  ( wr_addr ) == ( bv_8_32_n133 )  ;
assign n9252 =  ( n9250 ) & (n9251 )  ;
assign n9253 =  ( n9252 ) & (wr )  ;
assign n9254 =  ( n9253 ) ? ( n5071 ) : ( iram_32 ) ;
assign n9255 = wr_addr[7:7] ;
assign n9256 =  ( n9255 ) == ( bv_1_0_n53 )  ;
assign n9257 =  ( wr_addr ) == ( bv_8_32_n133 )  ;
assign n9258 =  ( n9256 ) & (n9257 )  ;
assign n9259 =  ( n9258 ) & (wr )  ;
assign n9260 =  ( n9259 ) ? ( n5096 ) : ( iram_32 ) ;
assign n9261 = wr_addr[7:7] ;
assign n9262 =  ( n9261 ) == ( bv_1_0_n53 )  ;
assign n9263 =  ( wr_addr ) == ( bv_8_32_n133 )  ;
assign n9264 =  ( n9262 ) & (n9263 )  ;
assign n9265 =  ( n9264 ) & (wr )  ;
assign n9266 =  ( n9265 ) ? ( n5123 ) : ( iram_32 ) ;
assign n9267 = wr_addr[7:7] ;
assign n9268 =  ( n9267 ) == ( bv_1_0_n53 )  ;
assign n9269 =  ( wr_addr ) == ( bv_8_32_n133 )  ;
assign n9270 =  ( n9268 ) & (n9269 )  ;
assign n9271 =  ( n9270 ) & (wr )  ;
assign n9272 =  ( n9271 ) ? ( n5165 ) : ( iram_32 ) ;
assign n9273 = wr_addr[7:7] ;
assign n9274 =  ( n9273 ) == ( bv_1_0_n53 )  ;
assign n9275 =  ( wr_addr ) == ( bv_8_32_n133 )  ;
assign n9276 =  ( n9274 ) & (n9275 )  ;
assign n9277 =  ( n9276 ) & (wr )  ;
assign n9278 =  ( n9277 ) ? ( n5204 ) : ( iram_32 ) ;
assign n9279 = wr_addr[7:7] ;
assign n9280 =  ( n9279 ) == ( bv_1_0_n53 )  ;
assign n9281 =  ( wr_addr ) == ( bv_8_32_n133 )  ;
assign n9282 =  ( n9280 ) & (n9281 )  ;
assign n9283 =  ( n9282 ) & (wr )  ;
assign n9284 =  ( n9283 ) ? ( n5262 ) : ( iram_32 ) ;
assign n9285 = wr_addr[7:7] ;
assign n9286 =  ( n9285 ) == ( bv_1_0_n53 )  ;
assign n9287 =  ( wr_addr ) == ( bv_8_32_n133 )  ;
assign n9288 =  ( n9286 ) & (n9287 )  ;
assign n9289 =  ( n9288 ) & (wr )  ;
assign n9290 =  ( n9289 ) ? ( n5298 ) : ( iram_32 ) ;
assign n9291 = wr_addr[7:7] ;
assign n9292 =  ( n9291 ) == ( bv_1_0_n53 )  ;
assign n9293 =  ( wr_addr ) == ( bv_8_32_n133 )  ;
assign n9294 =  ( n9292 ) & (n9293 )  ;
assign n9295 =  ( n9294 ) & (wr )  ;
assign n9296 =  ( n9295 ) ? ( n5325 ) : ( iram_32 ) ;
assign n9297 = wr_addr[7:7] ;
assign n9298 =  ( n9297 ) == ( bv_1_0_n53 )  ;
assign n9299 =  ( wr_addr ) == ( bv_8_33_n135 )  ;
assign n9300 =  ( n9298 ) & (n9299 )  ;
assign n9301 =  ( n9300 ) & (wr )  ;
assign n9302 =  ( n9301 ) ? ( n4782 ) : ( iram_33 ) ;
assign n9303 = wr_addr[7:7] ;
assign n9304 =  ( n9303 ) == ( bv_1_0_n53 )  ;
assign n9305 =  ( wr_addr ) == ( bv_8_33_n135 )  ;
assign n9306 =  ( n9304 ) & (n9305 )  ;
assign n9307 =  ( n9306 ) & (wr )  ;
assign n9308 =  ( n9307 ) ? ( n4841 ) : ( iram_33 ) ;
assign n9309 = wr_addr[7:7] ;
assign n9310 =  ( n9309 ) == ( bv_1_0_n53 )  ;
assign n9311 =  ( wr_addr ) == ( bv_8_33_n135 )  ;
assign n9312 =  ( n9310 ) & (n9311 )  ;
assign n9313 =  ( n9312 ) & (wr )  ;
assign n9314 =  ( n9313 ) ? ( n5449 ) : ( iram_33 ) ;
assign n9315 = wr_addr[7:7] ;
assign n9316 =  ( n9315 ) == ( bv_1_0_n53 )  ;
assign n9317 =  ( wr_addr ) == ( bv_8_33_n135 )  ;
assign n9318 =  ( n9316 ) & (n9317 )  ;
assign n9319 =  ( n9318 ) & (wr )  ;
assign n9320 =  ( n9319 ) ? ( n4906 ) : ( iram_33 ) ;
assign n9321 = wr_addr[7:7] ;
assign n9322 =  ( n9321 ) == ( bv_1_0_n53 )  ;
assign n9323 =  ( wr_addr ) == ( bv_8_33_n135 )  ;
assign n9324 =  ( n9322 ) & (n9323 )  ;
assign n9325 =  ( n9324 ) & (wr )  ;
assign n9326 =  ( n9325 ) ? ( n5485 ) : ( iram_33 ) ;
assign n9327 = wr_addr[7:7] ;
assign n9328 =  ( n9327 ) == ( bv_1_0_n53 )  ;
assign n9329 =  ( wr_addr ) == ( bv_8_33_n135 )  ;
assign n9330 =  ( n9328 ) & (n9329 )  ;
assign n9331 =  ( n9330 ) & (wr )  ;
assign n9332 =  ( n9331 ) ? ( n5512 ) : ( iram_33 ) ;
assign n9333 = wr_addr[7:7] ;
assign n9334 =  ( n9333 ) == ( bv_1_0_n53 )  ;
assign n9335 =  ( wr_addr ) == ( bv_8_33_n135 )  ;
assign n9336 =  ( n9334 ) & (n9335 )  ;
assign n9337 =  ( n9336 ) & (wr )  ;
assign n9338 =  ( n9337 ) ? ( bv_8_0_n69 ) : ( iram_33 ) ;
assign n9339 = wr_addr[7:7] ;
assign n9340 =  ( n9339 ) == ( bv_1_0_n53 )  ;
assign n9341 =  ( wr_addr ) == ( bv_8_33_n135 )  ;
assign n9342 =  ( n9340 ) & (n9341 )  ;
assign n9343 =  ( n9342 ) & (wr )  ;
assign n9344 =  ( n9343 ) ? ( n5071 ) : ( iram_33 ) ;
assign n9345 = wr_addr[7:7] ;
assign n9346 =  ( n9345 ) == ( bv_1_0_n53 )  ;
assign n9347 =  ( wr_addr ) == ( bv_8_33_n135 )  ;
assign n9348 =  ( n9346 ) & (n9347 )  ;
assign n9349 =  ( n9348 ) & (wr )  ;
assign n9350 =  ( n9349 ) ? ( n5096 ) : ( iram_33 ) ;
assign n9351 = wr_addr[7:7] ;
assign n9352 =  ( n9351 ) == ( bv_1_0_n53 )  ;
assign n9353 =  ( wr_addr ) == ( bv_8_33_n135 )  ;
assign n9354 =  ( n9352 ) & (n9353 )  ;
assign n9355 =  ( n9354 ) & (wr )  ;
assign n9356 =  ( n9355 ) ? ( n5123 ) : ( iram_33 ) ;
assign n9357 = wr_addr[7:7] ;
assign n9358 =  ( n9357 ) == ( bv_1_0_n53 )  ;
assign n9359 =  ( wr_addr ) == ( bv_8_33_n135 )  ;
assign n9360 =  ( n9358 ) & (n9359 )  ;
assign n9361 =  ( n9360 ) & (wr )  ;
assign n9362 =  ( n9361 ) ? ( n5165 ) : ( iram_33 ) ;
assign n9363 = wr_addr[7:7] ;
assign n9364 =  ( n9363 ) == ( bv_1_0_n53 )  ;
assign n9365 =  ( wr_addr ) == ( bv_8_33_n135 )  ;
assign n9366 =  ( n9364 ) & (n9365 )  ;
assign n9367 =  ( n9366 ) & (wr )  ;
assign n9368 =  ( n9367 ) ? ( n5204 ) : ( iram_33 ) ;
assign n9369 = wr_addr[7:7] ;
assign n9370 =  ( n9369 ) == ( bv_1_0_n53 )  ;
assign n9371 =  ( wr_addr ) == ( bv_8_33_n135 )  ;
assign n9372 =  ( n9370 ) & (n9371 )  ;
assign n9373 =  ( n9372 ) & (wr )  ;
assign n9374 =  ( n9373 ) ? ( n5262 ) : ( iram_33 ) ;
assign n9375 = wr_addr[7:7] ;
assign n9376 =  ( n9375 ) == ( bv_1_0_n53 )  ;
assign n9377 =  ( wr_addr ) == ( bv_8_33_n135 )  ;
assign n9378 =  ( n9376 ) & (n9377 )  ;
assign n9379 =  ( n9378 ) & (wr )  ;
assign n9380 =  ( n9379 ) ? ( n5298 ) : ( iram_33 ) ;
assign n9381 = wr_addr[7:7] ;
assign n9382 =  ( n9381 ) == ( bv_1_0_n53 )  ;
assign n9383 =  ( wr_addr ) == ( bv_8_33_n135 )  ;
assign n9384 =  ( n9382 ) & (n9383 )  ;
assign n9385 =  ( n9384 ) & (wr )  ;
assign n9386 =  ( n9385 ) ? ( n5325 ) : ( iram_33 ) ;
assign n9387 = wr_addr[7:7] ;
assign n9388 =  ( n9387 ) == ( bv_1_0_n53 )  ;
assign n9389 =  ( wr_addr ) == ( bv_8_34_n137 )  ;
assign n9390 =  ( n9388 ) & (n9389 )  ;
assign n9391 =  ( n9390 ) & (wr )  ;
assign n9392 =  ( n9391 ) ? ( n4782 ) : ( iram_34 ) ;
assign n9393 = wr_addr[7:7] ;
assign n9394 =  ( n9393 ) == ( bv_1_0_n53 )  ;
assign n9395 =  ( wr_addr ) == ( bv_8_34_n137 )  ;
assign n9396 =  ( n9394 ) & (n9395 )  ;
assign n9397 =  ( n9396 ) & (wr )  ;
assign n9398 =  ( n9397 ) ? ( n4841 ) : ( iram_34 ) ;
assign n9399 = wr_addr[7:7] ;
assign n9400 =  ( n9399 ) == ( bv_1_0_n53 )  ;
assign n9401 =  ( wr_addr ) == ( bv_8_34_n137 )  ;
assign n9402 =  ( n9400 ) & (n9401 )  ;
assign n9403 =  ( n9402 ) & (wr )  ;
assign n9404 =  ( n9403 ) ? ( n5449 ) : ( iram_34 ) ;
assign n9405 = wr_addr[7:7] ;
assign n9406 =  ( n9405 ) == ( bv_1_0_n53 )  ;
assign n9407 =  ( wr_addr ) == ( bv_8_34_n137 )  ;
assign n9408 =  ( n9406 ) & (n9407 )  ;
assign n9409 =  ( n9408 ) & (wr )  ;
assign n9410 =  ( n9409 ) ? ( n4906 ) : ( iram_34 ) ;
assign n9411 = wr_addr[7:7] ;
assign n9412 =  ( n9411 ) == ( bv_1_0_n53 )  ;
assign n9413 =  ( wr_addr ) == ( bv_8_34_n137 )  ;
assign n9414 =  ( n9412 ) & (n9413 )  ;
assign n9415 =  ( n9414 ) & (wr )  ;
assign n9416 =  ( n9415 ) ? ( n5485 ) : ( iram_34 ) ;
assign n9417 = wr_addr[7:7] ;
assign n9418 =  ( n9417 ) == ( bv_1_0_n53 )  ;
assign n9419 =  ( wr_addr ) == ( bv_8_34_n137 )  ;
assign n9420 =  ( n9418 ) & (n9419 )  ;
assign n9421 =  ( n9420 ) & (wr )  ;
assign n9422 =  ( n9421 ) ? ( n5512 ) : ( iram_34 ) ;
assign n9423 = wr_addr[7:7] ;
assign n9424 =  ( n9423 ) == ( bv_1_0_n53 )  ;
assign n9425 =  ( wr_addr ) == ( bv_8_34_n137 )  ;
assign n9426 =  ( n9424 ) & (n9425 )  ;
assign n9427 =  ( n9426 ) & (wr )  ;
assign n9428 =  ( n9427 ) ? ( bv_8_0_n69 ) : ( iram_34 ) ;
assign n9429 = wr_addr[7:7] ;
assign n9430 =  ( n9429 ) == ( bv_1_0_n53 )  ;
assign n9431 =  ( wr_addr ) == ( bv_8_34_n137 )  ;
assign n9432 =  ( n9430 ) & (n9431 )  ;
assign n9433 =  ( n9432 ) & (wr )  ;
assign n9434 =  ( n9433 ) ? ( n5071 ) : ( iram_34 ) ;
assign n9435 = wr_addr[7:7] ;
assign n9436 =  ( n9435 ) == ( bv_1_0_n53 )  ;
assign n9437 =  ( wr_addr ) == ( bv_8_34_n137 )  ;
assign n9438 =  ( n9436 ) & (n9437 )  ;
assign n9439 =  ( n9438 ) & (wr )  ;
assign n9440 =  ( n9439 ) ? ( n5096 ) : ( iram_34 ) ;
assign n9441 = wr_addr[7:7] ;
assign n9442 =  ( n9441 ) == ( bv_1_0_n53 )  ;
assign n9443 =  ( wr_addr ) == ( bv_8_34_n137 )  ;
assign n9444 =  ( n9442 ) & (n9443 )  ;
assign n9445 =  ( n9444 ) & (wr )  ;
assign n9446 =  ( n9445 ) ? ( n5123 ) : ( iram_34 ) ;
assign n9447 = wr_addr[7:7] ;
assign n9448 =  ( n9447 ) == ( bv_1_0_n53 )  ;
assign n9449 =  ( wr_addr ) == ( bv_8_34_n137 )  ;
assign n9450 =  ( n9448 ) & (n9449 )  ;
assign n9451 =  ( n9450 ) & (wr )  ;
assign n9452 =  ( n9451 ) ? ( n5165 ) : ( iram_34 ) ;
assign n9453 = wr_addr[7:7] ;
assign n9454 =  ( n9453 ) == ( bv_1_0_n53 )  ;
assign n9455 =  ( wr_addr ) == ( bv_8_34_n137 )  ;
assign n9456 =  ( n9454 ) & (n9455 )  ;
assign n9457 =  ( n9456 ) & (wr )  ;
assign n9458 =  ( n9457 ) ? ( n5204 ) : ( iram_34 ) ;
assign n9459 = wr_addr[7:7] ;
assign n9460 =  ( n9459 ) == ( bv_1_0_n53 )  ;
assign n9461 =  ( wr_addr ) == ( bv_8_34_n137 )  ;
assign n9462 =  ( n9460 ) & (n9461 )  ;
assign n9463 =  ( n9462 ) & (wr )  ;
assign n9464 =  ( n9463 ) ? ( n5262 ) : ( iram_34 ) ;
assign n9465 = wr_addr[7:7] ;
assign n9466 =  ( n9465 ) == ( bv_1_0_n53 )  ;
assign n9467 =  ( wr_addr ) == ( bv_8_34_n137 )  ;
assign n9468 =  ( n9466 ) & (n9467 )  ;
assign n9469 =  ( n9468 ) & (wr )  ;
assign n9470 =  ( n9469 ) ? ( n5298 ) : ( iram_34 ) ;
assign n9471 = wr_addr[7:7] ;
assign n9472 =  ( n9471 ) == ( bv_1_0_n53 )  ;
assign n9473 =  ( wr_addr ) == ( bv_8_34_n137 )  ;
assign n9474 =  ( n9472 ) & (n9473 )  ;
assign n9475 =  ( n9474 ) & (wr )  ;
assign n9476 =  ( n9475 ) ? ( n5325 ) : ( iram_34 ) ;
assign n9477 = wr_addr[7:7] ;
assign n9478 =  ( n9477 ) == ( bv_1_0_n53 )  ;
assign n9479 =  ( wr_addr ) == ( bv_8_35_n139 )  ;
assign n9480 =  ( n9478 ) & (n9479 )  ;
assign n9481 =  ( n9480 ) & (wr )  ;
assign n9482 =  ( n9481 ) ? ( n4782 ) : ( iram_35 ) ;
assign n9483 = wr_addr[7:7] ;
assign n9484 =  ( n9483 ) == ( bv_1_0_n53 )  ;
assign n9485 =  ( wr_addr ) == ( bv_8_35_n139 )  ;
assign n9486 =  ( n9484 ) & (n9485 )  ;
assign n9487 =  ( n9486 ) & (wr )  ;
assign n9488 =  ( n9487 ) ? ( n4841 ) : ( iram_35 ) ;
assign n9489 = wr_addr[7:7] ;
assign n9490 =  ( n9489 ) == ( bv_1_0_n53 )  ;
assign n9491 =  ( wr_addr ) == ( bv_8_35_n139 )  ;
assign n9492 =  ( n9490 ) & (n9491 )  ;
assign n9493 =  ( n9492 ) & (wr )  ;
assign n9494 =  ( n9493 ) ? ( n5449 ) : ( iram_35 ) ;
assign n9495 = wr_addr[7:7] ;
assign n9496 =  ( n9495 ) == ( bv_1_0_n53 )  ;
assign n9497 =  ( wr_addr ) == ( bv_8_35_n139 )  ;
assign n9498 =  ( n9496 ) & (n9497 )  ;
assign n9499 =  ( n9498 ) & (wr )  ;
assign n9500 =  ( n9499 ) ? ( n4906 ) : ( iram_35 ) ;
assign n9501 = wr_addr[7:7] ;
assign n9502 =  ( n9501 ) == ( bv_1_0_n53 )  ;
assign n9503 =  ( wr_addr ) == ( bv_8_35_n139 )  ;
assign n9504 =  ( n9502 ) & (n9503 )  ;
assign n9505 =  ( n9504 ) & (wr )  ;
assign n9506 =  ( n9505 ) ? ( n5485 ) : ( iram_35 ) ;
assign n9507 = wr_addr[7:7] ;
assign n9508 =  ( n9507 ) == ( bv_1_0_n53 )  ;
assign n9509 =  ( wr_addr ) == ( bv_8_35_n139 )  ;
assign n9510 =  ( n9508 ) & (n9509 )  ;
assign n9511 =  ( n9510 ) & (wr )  ;
assign n9512 =  ( n9511 ) ? ( n5512 ) : ( iram_35 ) ;
assign n9513 = wr_addr[7:7] ;
assign n9514 =  ( n9513 ) == ( bv_1_0_n53 )  ;
assign n9515 =  ( wr_addr ) == ( bv_8_35_n139 )  ;
assign n9516 =  ( n9514 ) & (n9515 )  ;
assign n9517 =  ( n9516 ) & (wr )  ;
assign n9518 =  ( n9517 ) ? ( bv_8_0_n69 ) : ( iram_35 ) ;
assign n9519 = wr_addr[7:7] ;
assign n9520 =  ( n9519 ) == ( bv_1_0_n53 )  ;
assign n9521 =  ( wr_addr ) == ( bv_8_35_n139 )  ;
assign n9522 =  ( n9520 ) & (n9521 )  ;
assign n9523 =  ( n9522 ) & (wr )  ;
assign n9524 =  ( n9523 ) ? ( n5071 ) : ( iram_35 ) ;
assign n9525 = wr_addr[7:7] ;
assign n9526 =  ( n9525 ) == ( bv_1_0_n53 )  ;
assign n9527 =  ( wr_addr ) == ( bv_8_35_n139 )  ;
assign n9528 =  ( n9526 ) & (n9527 )  ;
assign n9529 =  ( n9528 ) & (wr )  ;
assign n9530 =  ( n9529 ) ? ( n5096 ) : ( iram_35 ) ;
assign n9531 = wr_addr[7:7] ;
assign n9532 =  ( n9531 ) == ( bv_1_0_n53 )  ;
assign n9533 =  ( wr_addr ) == ( bv_8_35_n139 )  ;
assign n9534 =  ( n9532 ) & (n9533 )  ;
assign n9535 =  ( n9534 ) & (wr )  ;
assign n9536 =  ( n9535 ) ? ( n5123 ) : ( iram_35 ) ;
assign n9537 = wr_addr[7:7] ;
assign n9538 =  ( n9537 ) == ( bv_1_0_n53 )  ;
assign n9539 =  ( wr_addr ) == ( bv_8_35_n139 )  ;
assign n9540 =  ( n9538 ) & (n9539 )  ;
assign n9541 =  ( n9540 ) & (wr )  ;
assign n9542 =  ( n9541 ) ? ( n5165 ) : ( iram_35 ) ;
assign n9543 = wr_addr[7:7] ;
assign n9544 =  ( n9543 ) == ( bv_1_0_n53 )  ;
assign n9545 =  ( wr_addr ) == ( bv_8_35_n139 )  ;
assign n9546 =  ( n9544 ) & (n9545 )  ;
assign n9547 =  ( n9546 ) & (wr )  ;
assign n9548 =  ( n9547 ) ? ( n5204 ) : ( iram_35 ) ;
assign n9549 = wr_addr[7:7] ;
assign n9550 =  ( n9549 ) == ( bv_1_0_n53 )  ;
assign n9551 =  ( wr_addr ) == ( bv_8_35_n139 )  ;
assign n9552 =  ( n9550 ) & (n9551 )  ;
assign n9553 =  ( n9552 ) & (wr )  ;
assign n9554 =  ( n9553 ) ? ( n5262 ) : ( iram_35 ) ;
assign n9555 = wr_addr[7:7] ;
assign n9556 =  ( n9555 ) == ( bv_1_0_n53 )  ;
assign n9557 =  ( wr_addr ) == ( bv_8_35_n139 )  ;
assign n9558 =  ( n9556 ) & (n9557 )  ;
assign n9559 =  ( n9558 ) & (wr )  ;
assign n9560 =  ( n9559 ) ? ( n5298 ) : ( iram_35 ) ;
assign n9561 = wr_addr[7:7] ;
assign n9562 =  ( n9561 ) == ( bv_1_0_n53 )  ;
assign n9563 =  ( wr_addr ) == ( bv_8_35_n139 )  ;
assign n9564 =  ( n9562 ) & (n9563 )  ;
assign n9565 =  ( n9564 ) & (wr )  ;
assign n9566 =  ( n9565 ) ? ( n5325 ) : ( iram_35 ) ;
assign n9567 = wr_addr[7:7] ;
assign n9568 =  ( n9567 ) == ( bv_1_0_n53 )  ;
assign n9569 =  ( wr_addr ) == ( bv_8_36_n141 )  ;
assign n9570 =  ( n9568 ) & (n9569 )  ;
assign n9571 =  ( n9570 ) & (wr )  ;
assign n9572 =  ( n9571 ) ? ( n4782 ) : ( iram_36 ) ;
assign n9573 = wr_addr[7:7] ;
assign n9574 =  ( n9573 ) == ( bv_1_0_n53 )  ;
assign n9575 =  ( wr_addr ) == ( bv_8_36_n141 )  ;
assign n9576 =  ( n9574 ) & (n9575 )  ;
assign n9577 =  ( n9576 ) & (wr )  ;
assign n9578 =  ( n9577 ) ? ( n4841 ) : ( iram_36 ) ;
assign n9579 = wr_addr[7:7] ;
assign n9580 =  ( n9579 ) == ( bv_1_0_n53 )  ;
assign n9581 =  ( wr_addr ) == ( bv_8_36_n141 )  ;
assign n9582 =  ( n9580 ) & (n9581 )  ;
assign n9583 =  ( n9582 ) & (wr )  ;
assign n9584 =  ( n9583 ) ? ( n5449 ) : ( iram_36 ) ;
assign n9585 = wr_addr[7:7] ;
assign n9586 =  ( n9585 ) == ( bv_1_0_n53 )  ;
assign n9587 =  ( wr_addr ) == ( bv_8_36_n141 )  ;
assign n9588 =  ( n9586 ) & (n9587 )  ;
assign n9589 =  ( n9588 ) & (wr )  ;
assign n9590 =  ( n9589 ) ? ( n4906 ) : ( iram_36 ) ;
assign n9591 = wr_addr[7:7] ;
assign n9592 =  ( n9591 ) == ( bv_1_0_n53 )  ;
assign n9593 =  ( wr_addr ) == ( bv_8_36_n141 )  ;
assign n9594 =  ( n9592 ) & (n9593 )  ;
assign n9595 =  ( n9594 ) & (wr )  ;
assign n9596 =  ( n9595 ) ? ( n5485 ) : ( iram_36 ) ;
assign n9597 = wr_addr[7:7] ;
assign n9598 =  ( n9597 ) == ( bv_1_0_n53 )  ;
assign n9599 =  ( wr_addr ) == ( bv_8_36_n141 )  ;
assign n9600 =  ( n9598 ) & (n9599 )  ;
assign n9601 =  ( n9600 ) & (wr )  ;
assign n9602 =  ( n9601 ) ? ( n5512 ) : ( iram_36 ) ;
assign n9603 = wr_addr[7:7] ;
assign n9604 =  ( n9603 ) == ( bv_1_0_n53 )  ;
assign n9605 =  ( wr_addr ) == ( bv_8_36_n141 )  ;
assign n9606 =  ( n9604 ) & (n9605 )  ;
assign n9607 =  ( n9606 ) & (wr )  ;
assign n9608 =  ( n9607 ) ? ( bv_8_0_n69 ) : ( iram_36 ) ;
assign n9609 = wr_addr[7:7] ;
assign n9610 =  ( n9609 ) == ( bv_1_0_n53 )  ;
assign n9611 =  ( wr_addr ) == ( bv_8_36_n141 )  ;
assign n9612 =  ( n9610 ) & (n9611 )  ;
assign n9613 =  ( n9612 ) & (wr )  ;
assign n9614 =  ( n9613 ) ? ( n5071 ) : ( iram_36 ) ;
assign n9615 = wr_addr[7:7] ;
assign n9616 =  ( n9615 ) == ( bv_1_0_n53 )  ;
assign n9617 =  ( wr_addr ) == ( bv_8_36_n141 )  ;
assign n9618 =  ( n9616 ) & (n9617 )  ;
assign n9619 =  ( n9618 ) & (wr )  ;
assign n9620 =  ( n9619 ) ? ( n5096 ) : ( iram_36 ) ;
assign n9621 = wr_addr[7:7] ;
assign n9622 =  ( n9621 ) == ( bv_1_0_n53 )  ;
assign n9623 =  ( wr_addr ) == ( bv_8_36_n141 )  ;
assign n9624 =  ( n9622 ) & (n9623 )  ;
assign n9625 =  ( n9624 ) & (wr )  ;
assign n9626 =  ( n9625 ) ? ( n5123 ) : ( iram_36 ) ;
assign n9627 = wr_addr[7:7] ;
assign n9628 =  ( n9627 ) == ( bv_1_0_n53 )  ;
assign n9629 =  ( wr_addr ) == ( bv_8_36_n141 )  ;
assign n9630 =  ( n9628 ) & (n9629 )  ;
assign n9631 =  ( n9630 ) & (wr )  ;
assign n9632 =  ( n9631 ) ? ( n5165 ) : ( iram_36 ) ;
assign n9633 = wr_addr[7:7] ;
assign n9634 =  ( n9633 ) == ( bv_1_0_n53 )  ;
assign n9635 =  ( wr_addr ) == ( bv_8_36_n141 )  ;
assign n9636 =  ( n9634 ) & (n9635 )  ;
assign n9637 =  ( n9636 ) & (wr )  ;
assign n9638 =  ( n9637 ) ? ( n5204 ) : ( iram_36 ) ;
assign n9639 = wr_addr[7:7] ;
assign n9640 =  ( n9639 ) == ( bv_1_0_n53 )  ;
assign n9641 =  ( wr_addr ) == ( bv_8_36_n141 )  ;
assign n9642 =  ( n9640 ) & (n9641 )  ;
assign n9643 =  ( n9642 ) & (wr )  ;
assign n9644 =  ( n9643 ) ? ( n5262 ) : ( iram_36 ) ;
assign n9645 = wr_addr[7:7] ;
assign n9646 =  ( n9645 ) == ( bv_1_0_n53 )  ;
assign n9647 =  ( wr_addr ) == ( bv_8_36_n141 )  ;
assign n9648 =  ( n9646 ) & (n9647 )  ;
assign n9649 =  ( n9648 ) & (wr )  ;
assign n9650 =  ( n9649 ) ? ( n5298 ) : ( iram_36 ) ;
assign n9651 = wr_addr[7:7] ;
assign n9652 =  ( n9651 ) == ( bv_1_0_n53 )  ;
assign n9653 =  ( wr_addr ) == ( bv_8_36_n141 )  ;
assign n9654 =  ( n9652 ) & (n9653 )  ;
assign n9655 =  ( n9654 ) & (wr )  ;
assign n9656 =  ( n9655 ) ? ( n5325 ) : ( iram_36 ) ;
assign n9657 = wr_addr[7:7] ;
assign n9658 =  ( n9657 ) == ( bv_1_0_n53 )  ;
assign n9659 =  ( wr_addr ) == ( bv_8_37_n143 )  ;
assign n9660 =  ( n9658 ) & (n9659 )  ;
assign n9661 =  ( n9660 ) & (wr )  ;
assign n9662 =  ( n9661 ) ? ( n4782 ) : ( iram_37 ) ;
assign n9663 = wr_addr[7:7] ;
assign n9664 =  ( n9663 ) == ( bv_1_0_n53 )  ;
assign n9665 =  ( wr_addr ) == ( bv_8_37_n143 )  ;
assign n9666 =  ( n9664 ) & (n9665 )  ;
assign n9667 =  ( n9666 ) & (wr )  ;
assign n9668 =  ( n9667 ) ? ( n4841 ) : ( iram_37 ) ;
assign n9669 = wr_addr[7:7] ;
assign n9670 =  ( n9669 ) == ( bv_1_0_n53 )  ;
assign n9671 =  ( wr_addr ) == ( bv_8_37_n143 )  ;
assign n9672 =  ( n9670 ) & (n9671 )  ;
assign n9673 =  ( n9672 ) & (wr )  ;
assign n9674 =  ( n9673 ) ? ( n5449 ) : ( iram_37 ) ;
assign n9675 = wr_addr[7:7] ;
assign n9676 =  ( n9675 ) == ( bv_1_0_n53 )  ;
assign n9677 =  ( wr_addr ) == ( bv_8_37_n143 )  ;
assign n9678 =  ( n9676 ) & (n9677 )  ;
assign n9679 =  ( n9678 ) & (wr )  ;
assign n9680 =  ( n9679 ) ? ( n4906 ) : ( iram_37 ) ;
assign n9681 = wr_addr[7:7] ;
assign n9682 =  ( n9681 ) == ( bv_1_0_n53 )  ;
assign n9683 =  ( wr_addr ) == ( bv_8_37_n143 )  ;
assign n9684 =  ( n9682 ) & (n9683 )  ;
assign n9685 =  ( n9684 ) & (wr )  ;
assign n9686 =  ( n9685 ) ? ( n5485 ) : ( iram_37 ) ;
assign n9687 = wr_addr[7:7] ;
assign n9688 =  ( n9687 ) == ( bv_1_0_n53 )  ;
assign n9689 =  ( wr_addr ) == ( bv_8_37_n143 )  ;
assign n9690 =  ( n9688 ) & (n9689 )  ;
assign n9691 =  ( n9690 ) & (wr )  ;
assign n9692 =  ( n9691 ) ? ( n5512 ) : ( iram_37 ) ;
assign n9693 = wr_addr[7:7] ;
assign n9694 =  ( n9693 ) == ( bv_1_0_n53 )  ;
assign n9695 =  ( wr_addr ) == ( bv_8_37_n143 )  ;
assign n9696 =  ( n9694 ) & (n9695 )  ;
assign n9697 =  ( n9696 ) & (wr )  ;
assign n9698 =  ( n9697 ) ? ( bv_8_0_n69 ) : ( iram_37 ) ;
assign n9699 = wr_addr[7:7] ;
assign n9700 =  ( n9699 ) == ( bv_1_0_n53 )  ;
assign n9701 =  ( wr_addr ) == ( bv_8_37_n143 )  ;
assign n9702 =  ( n9700 ) & (n9701 )  ;
assign n9703 =  ( n9702 ) & (wr )  ;
assign n9704 =  ( n9703 ) ? ( n5071 ) : ( iram_37 ) ;
assign n9705 = wr_addr[7:7] ;
assign n9706 =  ( n9705 ) == ( bv_1_0_n53 )  ;
assign n9707 =  ( wr_addr ) == ( bv_8_37_n143 )  ;
assign n9708 =  ( n9706 ) & (n9707 )  ;
assign n9709 =  ( n9708 ) & (wr )  ;
assign n9710 =  ( n9709 ) ? ( n5096 ) : ( iram_37 ) ;
assign n9711 = wr_addr[7:7] ;
assign n9712 =  ( n9711 ) == ( bv_1_0_n53 )  ;
assign n9713 =  ( wr_addr ) == ( bv_8_37_n143 )  ;
assign n9714 =  ( n9712 ) & (n9713 )  ;
assign n9715 =  ( n9714 ) & (wr )  ;
assign n9716 =  ( n9715 ) ? ( n5123 ) : ( iram_37 ) ;
assign n9717 = wr_addr[7:7] ;
assign n9718 =  ( n9717 ) == ( bv_1_0_n53 )  ;
assign n9719 =  ( wr_addr ) == ( bv_8_37_n143 )  ;
assign n9720 =  ( n9718 ) & (n9719 )  ;
assign n9721 =  ( n9720 ) & (wr )  ;
assign n9722 =  ( n9721 ) ? ( n5165 ) : ( iram_37 ) ;
assign n9723 = wr_addr[7:7] ;
assign n9724 =  ( n9723 ) == ( bv_1_0_n53 )  ;
assign n9725 =  ( wr_addr ) == ( bv_8_37_n143 )  ;
assign n9726 =  ( n9724 ) & (n9725 )  ;
assign n9727 =  ( n9726 ) & (wr )  ;
assign n9728 =  ( n9727 ) ? ( n5204 ) : ( iram_37 ) ;
assign n9729 = wr_addr[7:7] ;
assign n9730 =  ( n9729 ) == ( bv_1_0_n53 )  ;
assign n9731 =  ( wr_addr ) == ( bv_8_37_n143 )  ;
assign n9732 =  ( n9730 ) & (n9731 )  ;
assign n9733 =  ( n9732 ) & (wr )  ;
assign n9734 =  ( n9733 ) ? ( n5262 ) : ( iram_37 ) ;
assign n9735 = wr_addr[7:7] ;
assign n9736 =  ( n9735 ) == ( bv_1_0_n53 )  ;
assign n9737 =  ( wr_addr ) == ( bv_8_37_n143 )  ;
assign n9738 =  ( n9736 ) & (n9737 )  ;
assign n9739 =  ( n9738 ) & (wr )  ;
assign n9740 =  ( n9739 ) ? ( n5298 ) : ( iram_37 ) ;
assign n9741 = wr_addr[7:7] ;
assign n9742 =  ( n9741 ) == ( bv_1_0_n53 )  ;
assign n9743 =  ( wr_addr ) == ( bv_8_37_n143 )  ;
assign n9744 =  ( n9742 ) & (n9743 )  ;
assign n9745 =  ( n9744 ) & (wr )  ;
assign n9746 =  ( n9745 ) ? ( n5325 ) : ( iram_37 ) ;
assign n9747 = wr_addr[7:7] ;
assign n9748 =  ( n9747 ) == ( bv_1_0_n53 )  ;
assign n9749 =  ( wr_addr ) == ( bv_8_38_n145 )  ;
assign n9750 =  ( n9748 ) & (n9749 )  ;
assign n9751 =  ( n9750 ) & (wr )  ;
assign n9752 =  ( n9751 ) ? ( n4782 ) : ( iram_38 ) ;
assign n9753 = wr_addr[7:7] ;
assign n9754 =  ( n9753 ) == ( bv_1_0_n53 )  ;
assign n9755 =  ( wr_addr ) == ( bv_8_38_n145 )  ;
assign n9756 =  ( n9754 ) & (n9755 )  ;
assign n9757 =  ( n9756 ) & (wr )  ;
assign n9758 =  ( n9757 ) ? ( n4841 ) : ( iram_38 ) ;
assign n9759 = wr_addr[7:7] ;
assign n9760 =  ( n9759 ) == ( bv_1_0_n53 )  ;
assign n9761 =  ( wr_addr ) == ( bv_8_38_n145 )  ;
assign n9762 =  ( n9760 ) & (n9761 )  ;
assign n9763 =  ( n9762 ) & (wr )  ;
assign n9764 =  ( n9763 ) ? ( n5449 ) : ( iram_38 ) ;
assign n9765 = wr_addr[7:7] ;
assign n9766 =  ( n9765 ) == ( bv_1_0_n53 )  ;
assign n9767 =  ( wr_addr ) == ( bv_8_38_n145 )  ;
assign n9768 =  ( n9766 ) & (n9767 )  ;
assign n9769 =  ( n9768 ) & (wr )  ;
assign n9770 =  ( n9769 ) ? ( n4906 ) : ( iram_38 ) ;
assign n9771 = wr_addr[7:7] ;
assign n9772 =  ( n9771 ) == ( bv_1_0_n53 )  ;
assign n9773 =  ( wr_addr ) == ( bv_8_38_n145 )  ;
assign n9774 =  ( n9772 ) & (n9773 )  ;
assign n9775 =  ( n9774 ) & (wr )  ;
assign n9776 =  ( n9775 ) ? ( n5485 ) : ( iram_38 ) ;
assign n9777 = wr_addr[7:7] ;
assign n9778 =  ( n9777 ) == ( bv_1_0_n53 )  ;
assign n9779 =  ( wr_addr ) == ( bv_8_38_n145 )  ;
assign n9780 =  ( n9778 ) & (n9779 )  ;
assign n9781 =  ( n9780 ) & (wr )  ;
assign n9782 =  ( n9781 ) ? ( n5512 ) : ( iram_38 ) ;
assign n9783 = wr_addr[7:7] ;
assign n9784 =  ( n9783 ) == ( bv_1_0_n53 )  ;
assign n9785 =  ( wr_addr ) == ( bv_8_38_n145 )  ;
assign n9786 =  ( n9784 ) & (n9785 )  ;
assign n9787 =  ( n9786 ) & (wr )  ;
assign n9788 =  ( n9787 ) ? ( bv_8_0_n69 ) : ( iram_38 ) ;
assign n9789 = wr_addr[7:7] ;
assign n9790 =  ( n9789 ) == ( bv_1_0_n53 )  ;
assign n9791 =  ( wr_addr ) == ( bv_8_38_n145 )  ;
assign n9792 =  ( n9790 ) & (n9791 )  ;
assign n9793 =  ( n9792 ) & (wr )  ;
assign n9794 =  ( n9793 ) ? ( n5071 ) : ( iram_38 ) ;
assign n9795 = wr_addr[7:7] ;
assign n9796 =  ( n9795 ) == ( bv_1_0_n53 )  ;
assign n9797 =  ( wr_addr ) == ( bv_8_38_n145 )  ;
assign n9798 =  ( n9796 ) & (n9797 )  ;
assign n9799 =  ( n9798 ) & (wr )  ;
assign n9800 =  ( n9799 ) ? ( n5096 ) : ( iram_38 ) ;
assign n9801 = wr_addr[7:7] ;
assign n9802 =  ( n9801 ) == ( bv_1_0_n53 )  ;
assign n9803 =  ( wr_addr ) == ( bv_8_38_n145 )  ;
assign n9804 =  ( n9802 ) & (n9803 )  ;
assign n9805 =  ( n9804 ) & (wr )  ;
assign n9806 =  ( n9805 ) ? ( n5123 ) : ( iram_38 ) ;
assign n9807 = wr_addr[7:7] ;
assign n9808 =  ( n9807 ) == ( bv_1_0_n53 )  ;
assign n9809 =  ( wr_addr ) == ( bv_8_38_n145 )  ;
assign n9810 =  ( n9808 ) & (n9809 )  ;
assign n9811 =  ( n9810 ) & (wr )  ;
assign n9812 =  ( n9811 ) ? ( n5165 ) : ( iram_38 ) ;
assign n9813 = wr_addr[7:7] ;
assign n9814 =  ( n9813 ) == ( bv_1_0_n53 )  ;
assign n9815 =  ( wr_addr ) == ( bv_8_38_n145 )  ;
assign n9816 =  ( n9814 ) & (n9815 )  ;
assign n9817 =  ( n9816 ) & (wr )  ;
assign n9818 =  ( n9817 ) ? ( n5204 ) : ( iram_38 ) ;
assign n9819 = wr_addr[7:7] ;
assign n9820 =  ( n9819 ) == ( bv_1_0_n53 )  ;
assign n9821 =  ( wr_addr ) == ( bv_8_38_n145 )  ;
assign n9822 =  ( n9820 ) & (n9821 )  ;
assign n9823 =  ( n9822 ) & (wr )  ;
assign n9824 =  ( n9823 ) ? ( n5262 ) : ( iram_38 ) ;
assign n9825 = wr_addr[7:7] ;
assign n9826 =  ( n9825 ) == ( bv_1_0_n53 )  ;
assign n9827 =  ( wr_addr ) == ( bv_8_38_n145 )  ;
assign n9828 =  ( n9826 ) & (n9827 )  ;
assign n9829 =  ( n9828 ) & (wr )  ;
assign n9830 =  ( n9829 ) ? ( n5298 ) : ( iram_38 ) ;
assign n9831 = wr_addr[7:7] ;
assign n9832 =  ( n9831 ) == ( bv_1_0_n53 )  ;
assign n9833 =  ( wr_addr ) == ( bv_8_38_n145 )  ;
assign n9834 =  ( n9832 ) & (n9833 )  ;
assign n9835 =  ( n9834 ) & (wr )  ;
assign n9836 =  ( n9835 ) ? ( n5325 ) : ( iram_38 ) ;
assign n9837 = wr_addr[7:7] ;
assign n9838 =  ( n9837 ) == ( bv_1_0_n53 )  ;
assign n9839 =  ( wr_addr ) == ( bv_8_39_n147 )  ;
assign n9840 =  ( n9838 ) & (n9839 )  ;
assign n9841 =  ( n9840 ) & (wr )  ;
assign n9842 =  ( n9841 ) ? ( n4782 ) : ( iram_39 ) ;
assign n9843 = wr_addr[7:7] ;
assign n9844 =  ( n9843 ) == ( bv_1_0_n53 )  ;
assign n9845 =  ( wr_addr ) == ( bv_8_39_n147 )  ;
assign n9846 =  ( n9844 ) & (n9845 )  ;
assign n9847 =  ( n9846 ) & (wr )  ;
assign n9848 =  ( n9847 ) ? ( n4841 ) : ( iram_39 ) ;
assign n9849 = wr_addr[7:7] ;
assign n9850 =  ( n9849 ) == ( bv_1_0_n53 )  ;
assign n9851 =  ( wr_addr ) == ( bv_8_39_n147 )  ;
assign n9852 =  ( n9850 ) & (n9851 )  ;
assign n9853 =  ( n9852 ) & (wr )  ;
assign n9854 =  ( n9853 ) ? ( n5449 ) : ( iram_39 ) ;
assign n9855 = wr_addr[7:7] ;
assign n9856 =  ( n9855 ) == ( bv_1_0_n53 )  ;
assign n9857 =  ( wr_addr ) == ( bv_8_39_n147 )  ;
assign n9858 =  ( n9856 ) & (n9857 )  ;
assign n9859 =  ( n9858 ) & (wr )  ;
assign n9860 =  ( n9859 ) ? ( n4906 ) : ( iram_39 ) ;
assign n9861 = wr_addr[7:7] ;
assign n9862 =  ( n9861 ) == ( bv_1_0_n53 )  ;
assign n9863 =  ( wr_addr ) == ( bv_8_39_n147 )  ;
assign n9864 =  ( n9862 ) & (n9863 )  ;
assign n9865 =  ( n9864 ) & (wr )  ;
assign n9866 =  ( n9865 ) ? ( n5485 ) : ( iram_39 ) ;
assign n9867 = wr_addr[7:7] ;
assign n9868 =  ( n9867 ) == ( bv_1_0_n53 )  ;
assign n9869 =  ( wr_addr ) == ( bv_8_39_n147 )  ;
assign n9870 =  ( n9868 ) & (n9869 )  ;
assign n9871 =  ( n9870 ) & (wr )  ;
assign n9872 =  ( n9871 ) ? ( n5512 ) : ( iram_39 ) ;
assign n9873 = wr_addr[7:7] ;
assign n9874 =  ( n9873 ) == ( bv_1_0_n53 )  ;
assign n9875 =  ( wr_addr ) == ( bv_8_39_n147 )  ;
assign n9876 =  ( n9874 ) & (n9875 )  ;
assign n9877 =  ( n9876 ) & (wr )  ;
assign n9878 =  ( n9877 ) ? ( bv_8_0_n69 ) : ( iram_39 ) ;
assign n9879 = wr_addr[7:7] ;
assign n9880 =  ( n9879 ) == ( bv_1_0_n53 )  ;
assign n9881 =  ( wr_addr ) == ( bv_8_39_n147 )  ;
assign n9882 =  ( n9880 ) & (n9881 )  ;
assign n9883 =  ( n9882 ) & (wr )  ;
assign n9884 =  ( n9883 ) ? ( n5071 ) : ( iram_39 ) ;
assign n9885 = wr_addr[7:7] ;
assign n9886 =  ( n9885 ) == ( bv_1_0_n53 )  ;
assign n9887 =  ( wr_addr ) == ( bv_8_39_n147 )  ;
assign n9888 =  ( n9886 ) & (n9887 )  ;
assign n9889 =  ( n9888 ) & (wr )  ;
assign n9890 =  ( n9889 ) ? ( n5096 ) : ( iram_39 ) ;
assign n9891 = wr_addr[7:7] ;
assign n9892 =  ( n9891 ) == ( bv_1_0_n53 )  ;
assign n9893 =  ( wr_addr ) == ( bv_8_39_n147 )  ;
assign n9894 =  ( n9892 ) & (n9893 )  ;
assign n9895 =  ( n9894 ) & (wr )  ;
assign n9896 =  ( n9895 ) ? ( n5123 ) : ( iram_39 ) ;
assign n9897 = wr_addr[7:7] ;
assign n9898 =  ( n9897 ) == ( bv_1_0_n53 )  ;
assign n9899 =  ( wr_addr ) == ( bv_8_39_n147 )  ;
assign n9900 =  ( n9898 ) & (n9899 )  ;
assign n9901 =  ( n9900 ) & (wr )  ;
assign n9902 =  ( n9901 ) ? ( n5165 ) : ( iram_39 ) ;
assign n9903 = wr_addr[7:7] ;
assign n9904 =  ( n9903 ) == ( bv_1_0_n53 )  ;
assign n9905 =  ( wr_addr ) == ( bv_8_39_n147 )  ;
assign n9906 =  ( n9904 ) & (n9905 )  ;
assign n9907 =  ( n9906 ) & (wr )  ;
assign n9908 =  ( n9907 ) ? ( n5204 ) : ( iram_39 ) ;
assign n9909 = wr_addr[7:7] ;
assign n9910 =  ( n9909 ) == ( bv_1_0_n53 )  ;
assign n9911 =  ( wr_addr ) == ( bv_8_39_n147 )  ;
assign n9912 =  ( n9910 ) & (n9911 )  ;
assign n9913 =  ( n9912 ) & (wr )  ;
assign n9914 =  ( n9913 ) ? ( n5262 ) : ( iram_39 ) ;
assign n9915 = wr_addr[7:7] ;
assign n9916 =  ( n9915 ) == ( bv_1_0_n53 )  ;
assign n9917 =  ( wr_addr ) == ( bv_8_39_n147 )  ;
assign n9918 =  ( n9916 ) & (n9917 )  ;
assign n9919 =  ( n9918 ) & (wr )  ;
assign n9920 =  ( n9919 ) ? ( n5298 ) : ( iram_39 ) ;
assign n9921 = wr_addr[7:7] ;
assign n9922 =  ( n9921 ) == ( bv_1_0_n53 )  ;
assign n9923 =  ( wr_addr ) == ( bv_8_39_n147 )  ;
assign n9924 =  ( n9922 ) & (n9923 )  ;
assign n9925 =  ( n9924 ) & (wr )  ;
assign n9926 =  ( n9925 ) ? ( n5325 ) : ( iram_39 ) ;
assign n9927 = wr_addr[7:7] ;
assign n9928 =  ( n9927 ) == ( bv_1_0_n53 )  ;
assign n9929 =  ( wr_addr ) == ( bv_8_40_n149 )  ;
assign n9930 =  ( n9928 ) & (n9929 )  ;
assign n9931 =  ( n9930 ) & (wr )  ;
assign n9932 =  ( n9931 ) ? ( n4782 ) : ( iram_40 ) ;
assign n9933 = wr_addr[7:7] ;
assign n9934 =  ( n9933 ) == ( bv_1_0_n53 )  ;
assign n9935 =  ( wr_addr ) == ( bv_8_40_n149 )  ;
assign n9936 =  ( n9934 ) & (n9935 )  ;
assign n9937 =  ( n9936 ) & (wr )  ;
assign n9938 =  ( n9937 ) ? ( n4841 ) : ( iram_40 ) ;
assign n9939 = wr_addr[7:7] ;
assign n9940 =  ( n9939 ) == ( bv_1_0_n53 )  ;
assign n9941 =  ( wr_addr ) == ( bv_8_40_n149 )  ;
assign n9942 =  ( n9940 ) & (n9941 )  ;
assign n9943 =  ( n9942 ) & (wr )  ;
assign n9944 =  ( n9943 ) ? ( n5449 ) : ( iram_40 ) ;
assign n9945 = wr_addr[7:7] ;
assign n9946 =  ( n9945 ) == ( bv_1_0_n53 )  ;
assign n9947 =  ( wr_addr ) == ( bv_8_40_n149 )  ;
assign n9948 =  ( n9946 ) & (n9947 )  ;
assign n9949 =  ( n9948 ) & (wr )  ;
assign n9950 =  ( n9949 ) ? ( n4906 ) : ( iram_40 ) ;
assign n9951 = wr_addr[7:7] ;
assign n9952 =  ( n9951 ) == ( bv_1_0_n53 )  ;
assign n9953 =  ( wr_addr ) == ( bv_8_40_n149 )  ;
assign n9954 =  ( n9952 ) & (n9953 )  ;
assign n9955 =  ( n9954 ) & (wr )  ;
assign n9956 =  ( n9955 ) ? ( n5485 ) : ( iram_40 ) ;
assign n9957 = wr_addr[7:7] ;
assign n9958 =  ( n9957 ) == ( bv_1_0_n53 )  ;
assign n9959 =  ( wr_addr ) == ( bv_8_40_n149 )  ;
assign n9960 =  ( n9958 ) & (n9959 )  ;
assign n9961 =  ( n9960 ) & (wr )  ;
assign n9962 =  ( n9961 ) ? ( n5512 ) : ( iram_40 ) ;
assign n9963 = wr_addr[7:7] ;
assign n9964 =  ( n9963 ) == ( bv_1_0_n53 )  ;
assign n9965 =  ( wr_addr ) == ( bv_8_40_n149 )  ;
assign n9966 =  ( n9964 ) & (n9965 )  ;
assign n9967 =  ( n9966 ) & (wr )  ;
assign n9968 =  ( n9967 ) ? ( bv_8_0_n69 ) : ( iram_40 ) ;
assign n9969 = wr_addr[7:7] ;
assign n9970 =  ( n9969 ) == ( bv_1_0_n53 )  ;
assign n9971 =  ( wr_addr ) == ( bv_8_40_n149 )  ;
assign n9972 =  ( n9970 ) & (n9971 )  ;
assign n9973 =  ( n9972 ) & (wr )  ;
assign n9974 =  ( n9973 ) ? ( n5071 ) : ( iram_40 ) ;
assign n9975 = wr_addr[7:7] ;
assign n9976 =  ( n9975 ) == ( bv_1_0_n53 )  ;
assign n9977 =  ( wr_addr ) == ( bv_8_40_n149 )  ;
assign n9978 =  ( n9976 ) & (n9977 )  ;
assign n9979 =  ( n9978 ) & (wr )  ;
assign n9980 =  ( n9979 ) ? ( n5096 ) : ( iram_40 ) ;
assign n9981 = wr_addr[7:7] ;
assign n9982 =  ( n9981 ) == ( bv_1_0_n53 )  ;
assign n9983 =  ( wr_addr ) == ( bv_8_40_n149 )  ;
assign n9984 =  ( n9982 ) & (n9983 )  ;
assign n9985 =  ( n9984 ) & (wr )  ;
assign n9986 =  ( n9985 ) ? ( n5123 ) : ( iram_40 ) ;
assign n9987 = wr_addr[7:7] ;
assign n9988 =  ( n9987 ) == ( bv_1_0_n53 )  ;
assign n9989 =  ( wr_addr ) == ( bv_8_40_n149 )  ;
assign n9990 =  ( n9988 ) & (n9989 )  ;
assign n9991 =  ( n9990 ) & (wr )  ;
assign n9992 =  ( n9991 ) ? ( n5165 ) : ( iram_40 ) ;
assign n9993 = wr_addr[7:7] ;
assign n9994 =  ( n9993 ) == ( bv_1_0_n53 )  ;
assign n9995 =  ( wr_addr ) == ( bv_8_40_n149 )  ;
assign n9996 =  ( n9994 ) & (n9995 )  ;
assign n9997 =  ( n9996 ) & (wr )  ;
assign n9998 =  ( n9997 ) ? ( n5204 ) : ( iram_40 ) ;
assign n9999 = wr_addr[7:7] ;
assign n10000 =  ( n9999 ) == ( bv_1_0_n53 )  ;
assign n10001 =  ( wr_addr ) == ( bv_8_40_n149 )  ;
assign n10002 =  ( n10000 ) & (n10001 )  ;
assign n10003 =  ( n10002 ) & (wr )  ;
assign n10004 =  ( n10003 ) ? ( n5262 ) : ( iram_40 ) ;
assign n10005 = wr_addr[7:7] ;
assign n10006 =  ( n10005 ) == ( bv_1_0_n53 )  ;
assign n10007 =  ( wr_addr ) == ( bv_8_40_n149 )  ;
assign n10008 =  ( n10006 ) & (n10007 )  ;
assign n10009 =  ( n10008 ) & (wr )  ;
assign n10010 =  ( n10009 ) ? ( n5298 ) : ( iram_40 ) ;
assign n10011 = wr_addr[7:7] ;
assign n10012 =  ( n10011 ) == ( bv_1_0_n53 )  ;
assign n10013 =  ( wr_addr ) == ( bv_8_40_n149 )  ;
assign n10014 =  ( n10012 ) & (n10013 )  ;
assign n10015 =  ( n10014 ) & (wr )  ;
assign n10016 =  ( n10015 ) ? ( n5325 ) : ( iram_40 ) ;
assign n10017 = wr_addr[7:7] ;
assign n10018 =  ( n10017 ) == ( bv_1_0_n53 )  ;
assign n10019 =  ( wr_addr ) == ( bv_8_41_n151 )  ;
assign n10020 =  ( n10018 ) & (n10019 )  ;
assign n10021 =  ( n10020 ) & (wr )  ;
assign n10022 =  ( n10021 ) ? ( n4782 ) : ( iram_41 ) ;
assign n10023 = wr_addr[7:7] ;
assign n10024 =  ( n10023 ) == ( bv_1_0_n53 )  ;
assign n10025 =  ( wr_addr ) == ( bv_8_41_n151 )  ;
assign n10026 =  ( n10024 ) & (n10025 )  ;
assign n10027 =  ( n10026 ) & (wr )  ;
assign n10028 =  ( n10027 ) ? ( n4841 ) : ( iram_41 ) ;
assign n10029 = wr_addr[7:7] ;
assign n10030 =  ( n10029 ) == ( bv_1_0_n53 )  ;
assign n10031 =  ( wr_addr ) == ( bv_8_41_n151 )  ;
assign n10032 =  ( n10030 ) & (n10031 )  ;
assign n10033 =  ( n10032 ) & (wr )  ;
assign n10034 =  ( n10033 ) ? ( n5449 ) : ( iram_41 ) ;
assign n10035 = wr_addr[7:7] ;
assign n10036 =  ( n10035 ) == ( bv_1_0_n53 )  ;
assign n10037 =  ( wr_addr ) == ( bv_8_41_n151 )  ;
assign n10038 =  ( n10036 ) & (n10037 )  ;
assign n10039 =  ( n10038 ) & (wr )  ;
assign n10040 =  ( n10039 ) ? ( n4906 ) : ( iram_41 ) ;
assign n10041 = wr_addr[7:7] ;
assign n10042 =  ( n10041 ) == ( bv_1_0_n53 )  ;
assign n10043 =  ( wr_addr ) == ( bv_8_41_n151 )  ;
assign n10044 =  ( n10042 ) & (n10043 )  ;
assign n10045 =  ( n10044 ) & (wr )  ;
assign n10046 =  ( n10045 ) ? ( n5485 ) : ( iram_41 ) ;
assign n10047 = wr_addr[7:7] ;
assign n10048 =  ( n10047 ) == ( bv_1_0_n53 )  ;
assign n10049 =  ( wr_addr ) == ( bv_8_41_n151 )  ;
assign n10050 =  ( n10048 ) & (n10049 )  ;
assign n10051 =  ( n10050 ) & (wr )  ;
assign n10052 =  ( n10051 ) ? ( n5512 ) : ( iram_41 ) ;
assign n10053 = wr_addr[7:7] ;
assign n10054 =  ( n10053 ) == ( bv_1_0_n53 )  ;
assign n10055 =  ( wr_addr ) == ( bv_8_41_n151 )  ;
assign n10056 =  ( n10054 ) & (n10055 )  ;
assign n10057 =  ( n10056 ) & (wr )  ;
assign n10058 =  ( n10057 ) ? ( bv_8_0_n69 ) : ( iram_41 ) ;
assign n10059 = wr_addr[7:7] ;
assign n10060 =  ( n10059 ) == ( bv_1_0_n53 )  ;
assign n10061 =  ( wr_addr ) == ( bv_8_41_n151 )  ;
assign n10062 =  ( n10060 ) & (n10061 )  ;
assign n10063 =  ( n10062 ) & (wr )  ;
assign n10064 =  ( n10063 ) ? ( n5071 ) : ( iram_41 ) ;
assign n10065 = wr_addr[7:7] ;
assign n10066 =  ( n10065 ) == ( bv_1_0_n53 )  ;
assign n10067 =  ( wr_addr ) == ( bv_8_41_n151 )  ;
assign n10068 =  ( n10066 ) & (n10067 )  ;
assign n10069 =  ( n10068 ) & (wr )  ;
assign n10070 =  ( n10069 ) ? ( n5096 ) : ( iram_41 ) ;
assign n10071 = wr_addr[7:7] ;
assign n10072 =  ( n10071 ) == ( bv_1_0_n53 )  ;
assign n10073 =  ( wr_addr ) == ( bv_8_41_n151 )  ;
assign n10074 =  ( n10072 ) & (n10073 )  ;
assign n10075 =  ( n10074 ) & (wr )  ;
assign n10076 =  ( n10075 ) ? ( n5123 ) : ( iram_41 ) ;
assign n10077 = wr_addr[7:7] ;
assign n10078 =  ( n10077 ) == ( bv_1_0_n53 )  ;
assign n10079 =  ( wr_addr ) == ( bv_8_41_n151 )  ;
assign n10080 =  ( n10078 ) & (n10079 )  ;
assign n10081 =  ( n10080 ) & (wr )  ;
assign n10082 =  ( n10081 ) ? ( n5165 ) : ( iram_41 ) ;
assign n10083 = wr_addr[7:7] ;
assign n10084 =  ( n10083 ) == ( bv_1_0_n53 )  ;
assign n10085 =  ( wr_addr ) == ( bv_8_41_n151 )  ;
assign n10086 =  ( n10084 ) & (n10085 )  ;
assign n10087 =  ( n10086 ) & (wr )  ;
assign n10088 =  ( n10087 ) ? ( n5204 ) : ( iram_41 ) ;
assign n10089 = wr_addr[7:7] ;
assign n10090 =  ( n10089 ) == ( bv_1_0_n53 )  ;
assign n10091 =  ( wr_addr ) == ( bv_8_41_n151 )  ;
assign n10092 =  ( n10090 ) & (n10091 )  ;
assign n10093 =  ( n10092 ) & (wr )  ;
assign n10094 =  ( n10093 ) ? ( n5262 ) : ( iram_41 ) ;
assign n10095 = wr_addr[7:7] ;
assign n10096 =  ( n10095 ) == ( bv_1_0_n53 )  ;
assign n10097 =  ( wr_addr ) == ( bv_8_41_n151 )  ;
assign n10098 =  ( n10096 ) & (n10097 )  ;
assign n10099 =  ( n10098 ) & (wr )  ;
assign n10100 =  ( n10099 ) ? ( n5298 ) : ( iram_41 ) ;
assign n10101 = wr_addr[7:7] ;
assign n10102 =  ( n10101 ) == ( bv_1_0_n53 )  ;
assign n10103 =  ( wr_addr ) == ( bv_8_41_n151 )  ;
assign n10104 =  ( n10102 ) & (n10103 )  ;
assign n10105 =  ( n10104 ) & (wr )  ;
assign n10106 =  ( n10105 ) ? ( n5325 ) : ( iram_41 ) ;
assign n10107 = wr_addr[7:7] ;
assign n10108 =  ( n10107 ) == ( bv_1_0_n53 )  ;
assign n10109 =  ( wr_addr ) == ( bv_8_42_n153 )  ;
assign n10110 =  ( n10108 ) & (n10109 )  ;
assign n10111 =  ( n10110 ) & (wr )  ;
assign n10112 =  ( n10111 ) ? ( n4782 ) : ( iram_42 ) ;
assign n10113 = wr_addr[7:7] ;
assign n10114 =  ( n10113 ) == ( bv_1_0_n53 )  ;
assign n10115 =  ( wr_addr ) == ( bv_8_42_n153 )  ;
assign n10116 =  ( n10114 ) & (n10115 )  ;
assign n10117 =  ( n10116 ) & (wr )  ;
assign n10118 =  ( n10117 ) ? ( n4841 ) : ( iram_42 ) ;
assign n10119 = wr_addr[7:7] ;
assign n10120 =  ( n10119 ) == ( bv_1_0_n53 )  ;
assign n10121 =  ( wr_addr ) == ( bv_8_42_n153 )  ;
assign n10122 =  ( n10120 ) & (n10121 )  ;
assign n10123 =  ( n10122 ) & (wr )  ;
assign n10124 =  ( n10123 ) ? ( n5449 ) : ( iram_42 ) ;
assign n10125 = wr_addr[7:7] ;
assign n10126 =  ( n10125 ) == ( bv_1_0_n53 )  ;
assign n10127 =  ( wr_addr ) == ( bv_8_42_n153 )  ;
assign n10128 =  ( n10126 ) & (n10127 )  ;
assign n10129 =  ( n10128 ) & (wr )  ;
assign n10130 =  ( n10129 ) ? ( n4906 ) : ( iram_42 ) ;
assign n10131 = wr_addr[7:7] ;
assign n10132 =  ( n10131 ) == ( bv_1_0_n53 )  ;
assign n10133 =  ( wr_addr ) == ( bv_8_42_n153 )  ;
assign n10134 =  ( n10132 ) & (n10133 )  ;
assign n10135 =  ( n10134 ) & (wr )  ;
assign n10136 =  ( n10135 ) ? ( n5485 ) : ( iram_42 ) ;
assign n10137 = wr_addr[7:7] ;
assign n10138 =  ( n10137 ) == ( bv_1_0_n53 )  ;
assign n10139 =  ( wr_addr ) == ( bv_8_42_n153 )  ;
assign n10140 =  ( n10138 ) & (n10139 )  ;
assign n10141 =  ( n10140 ) & (wr )  ;
assign n10142 =  ( n10141 ) ? ( n5512 ) : ( iram_42 ) ;
assign n10143 = wr_addr[7:7] ;
assign n10144 =  ( n10143 ) == ( bv_1_0_n53 )  ;
assign n10145 =  ( wr_addr ) == ( bv_8_42_n153 )  ;
assign n10146 =  ( n10144 ) & (n10145 )  ;
assign n10147 =  ( n10146 ) & (wr )  ;
assign n10148 =  ( n10147 ) ? ( bv_8_0_n69 ) : ( iram_42 ) ;
assign n10149 = wr_addr[7:7] ;
assign n10150 =  ( n10149 ) == ( bv_1_0_n53 )  ;
assign n10151 =  ( wr_addr ) == ( bv_8_42_n153 )  ;
assign n10152 =  ( n10150 ) & (n10151 )  ;
assign n10153 =  ( n10152 ) & (wr )  ;
assign n10154 =  ( n10153 ) ? ( n5071 ) : ( iram_42 ) ;
assign n10155 = wr_addr[7:7] ;
assign n10156 =  ( n10155 ) == ( bv_1_0_n53 )  ;
assign n10157 =  ( wr_addr ) == ( bv_8_42_n153 )  ;
assign n10158 =  ( n10156 ) & (n10157 )  ;
assign n10159 =  ( n10158 ) & (wr )  ;
assign n10160 =  ( n10159 ) ? ( n5096 ) : ( iram_42 ) ;
assign n10161 = wr_addr[7:7] ;
assign n10162 =  ( n10161 ) == ( bv_1_0_n53 )  ;
assign n10163 =  ( wr_addr ) == ( bv_8_42_n153 )  ;
assign n10164 =  ( n10162 ) & (n10163 )  ;
assign n10165 =  ( n10164 ) & (wr )  ;
assign n10166 =  ( n10165 ) ? ( n5123 ) : ( iram_42 ) ;
assign n10167 = wr_addr[7:7] ;
assign n10168 =  ( n10167 ) == ( bv_1_0_n53 )  ;
assign n10169 =  ( wr_addr ) == ( bv_8_42_n153 )  ;
assign n10170 =  ( n10168 ) & (n10169 )  ;
assign n10171 =  ( n10170 ) & (wr )  ;
assign n10172 =  ( n10171 ) ? ( n5165 ) : ( iram_42 ) ;
assign n10173 = wr_addr[7:7] ;
assign n10174 =  ( n10173 ) == ( bv_1_0_n53 )  ;
assign n10175 =  ( wr_addr ) == ( bv_8_42_n153 )  ;
assign n10176 =  ( n10174 ) & (n10175 )  ;
assign n10177 =  ( n10176 ) & (wr )  ;
assign n10178 =  ( n10177 ) ? ( n5204 ) : ( iram_42 ) ;
assign n10179 = wr_addr[7:7] ;
assign n10180 =  ( n10179 ) == ( bv_1_0_n53 )  ;
assign n10181 =  ( wr_addr ) == ( bv_8_42_n153 )  ;
assign n10182 =  ( n10180 ) & (n10181 )  ;
assign n10183 =  ( n10182 ) & (wr )  ;
assign n10184 =  ( n10183 ) ? ( n5262 ) : ( iram_42 ) ;
assign n10185 = wr_addr[7:7] ;
assign n10186 =  ( n10185 ) == ( bv_1_0_n53 )  ;
assign n10187 =  ( wr_addr ) == ( bv_8_42_n153 )  ;
assign n10188 =  ( n10186 ) & (n10187 )  ;
assign n10189 =  ( n10188 ) & (wr )  ;
assign n10190 =  ( n10189 ) ? ( n5298 ) : ( iram_42 ) ;
assign n10191 = wr_addr[7:7] ;
assign n10192 =  ( n10191 ) == ( bv_1_0_n53 )  ;
assign n10193 =  ( wr_addr ) == ( bv_8_42_n153 )  ;
assign n10194 =  ( n10192 ) & (n10193 )  ;
assign n10195 =  ( n10194 ) & (wr )  ;
assign n10196 =  ( n10195 ) ? ( n5325 ) : ( iram_42 ) ;
assign n10197 = wr_addr[7:7] ;
assign n10198 =  ( n10197 ) == ( bv_1_0_n53 )  ;
assign n10199 =  ( wr_addr ) == ( bv_8_43_n155 )  ;
assign n10200 =  ( n10198 ) & (n10199 )  ;
assign n10201 =  ( n10200 ) & (wr )  ;
assign n10202 =  ( n10201 ) ? ( n4782 ) : ( iram_43 ) ;
assign n10203 = wr_addr[7:7] ;
assign n10204 =  ( n10203 ) == ( bv_1_0_n53 )  ;
assign n10205 =  ( wr_addr ) == ( bv_8_43_n155 )  ;
assign n10206 =  ( n10204 ) & (n10205 )  ;
assign n10207 =  ( n10206 ) & (wr )  ;
assign n10208 =  ( n10207 ) ? ( n4841 ) : ( iram_43 ) ;
assign n10209 = wr_addr[7:7] ;
assign n10210 =  ( n10209 ) == ( bv_1_0_n53 )  ;
assign n10211 =  ( wr_addr ) == ( bv_8_43_n155 )  ;
assign n10212 =  ( n10210 ) & (n10211 )  ;
assign n10213 =  ( n10212 ) & (wr )  ;
assign n10214 =  ( n10213 ) ? ( n5449 ) : ( iram_43 ) ;
assign n10215 = wr_addr[7:7] ;
assign n10216 =  ( n10215 ) == ( bv_1_0_n53 )  ;
assign n10217 =  ( wr_addr ) == ( bv_8_43_n155 )  ;
assign n10218 =  ( n10216 ) & (n10217 )  ;
assign n10219 =  ( n10218 ) & (wr )  ;
assign n10220 =  ( n10219 ) ? ( n4906 ) : ( iram_43 ) ;
assign n10221 = wr_addr[7:7] ;
assign n10222 =  ( n10221 ) == ( bv_1_0_n53 )  ;
assign n10223 =  ( wr_addr ) == ( bv_8_43_n155 )  ;
assign n10224 =  ( n10222 ) & (n10223 )  ;
assign n10225 =  ( n10224 ) & (wr )  ;
assign n10226 =  ( n10225 ) ? ( n5485 ) : ( iram_43 ) ;
assign n10227 = wr_addr[7:7] ;
assign n10228 =  ( n10227 ) == ( bv_1_0_n53 )  ;
assign n10229 =  ( wr_addr ) == ( bv_8_43_n155 )  ;
assign n10230 =  ( n10228 ) & (n10229 )  ;
assign n10231 =  ( n10230 ) & (wr )  ;
assign n10232 =  ( n10231 ) ? ( n5512 ) : ( iram_43 ) ;
assign n10233 = wr_addr[7:7] ;
assign n10234 =  ( n10233 ) == ( bv_1_0_n53 )  ;
assign n10235 =  ( wr_addr ) == ( bv_8_43_n155 )  ;
assign n10236 =  ( n10234 ) & (n10235 )  ;
assign n10237 =  ( n10236 ) & (wr )  ;
assign n10238 =  ( n10237 ) ? ( bv_8_0_n69 ) : ( iram_43 ) ;
assign n10239 = wr_addr[7:7] ;
assign n10240 =  ( n10239 ) == ( bv_1_0_n53 )  ;
assign n10241 =  ( wr_addr ) == ( bv_8_43_n155 )  ;
assign n10242 =  ( n10240 ) & (n10241 )  ;
assign n10243 =  ( n10242 ) & (wr )  ;
assign n10244 =  ( n10243 ) ? ( n5071 ) : ( iram_43 ) ;
assign n10245 = wr_addr[7:7] ;
assign n10246 =  ( n10245 ) == ( bv_1_0_n53 )  ;
assign n10247 =  ( wr_addr ) == ( bv_8_43_n155 )  ;
assign n10248 =  ( n10246 ) & (n10247 )  ;
assign n10249 =  ( n10248 ) & (wr )  ;
assign n10250 =  ( n10249 ) ? ( n5096 ) : ( iram_43 ) ;
assign n10251 = wr_addr[7:7] ;
assign n10252 =  ( n10251 ) == ( bv_1_0_n53 )  ;
assign n10253 =  ( wr_addr ) == ( bv_8_43_n155 )  ;
assign n10254 =  ( n10252 ) & (n10253 )  ;
assign n10255 =  ( n10254 ) & (wr )  ;
assign n10256 =  ( n10255 ) ? ( n5123 ) : ( iram_43 ) ;
assign n10257 = wr_addr[7:7] ;
assign n10258 =  ( n10257 ) == ( bv_1_0_n53 )  ;
assign n10259 =  ( wr_addr ) == ( bv_8_43_n155 )  ;
assign n10260 =  ( n10258 ) & (n10259 )  ;
assign n10261 =  ( n10260 ) & (wr )  ;
assign n10262 =  ( n10261 ) ? ( n5165 ) : ( iram_43 ) ;
assign n10263 = wr_addr[7:7] ;
assign n10264 =  ( n10263 ) == ( bv_1_0_n53 )  ;
assign n10265 =  ( wr_addr ) == ( bv_8_43_n155 )  ;
assign n10266 =  ( n10264 ) & (n10265 )  ;
assign n10267 =  ( n10266 ) & (wr )  ;
assign n10268 =  ( n10267 ) ? ( n5204 ) : ( iram_43 ) ;
assign n10269 = wr_addr[7:7] ;
assign n10270 =  ( n10269 ) == ( bv_1_0_n53 )  ;
assign n10271 =  ( wr_addr ) == ( bv_8_43_n155 )  ;
assign n10272 =  ( n10270 ) & (n10271 )  ;
assign n10273 =  ( n10272 ) & (wr )  ;
assign n10274 =  ( n10273 ) ? ( n5262 ) : ( iram_43 ) ;
assign n10275 = wr_addr[7:7] ;
assign n10276 =  ( n10275 ) == ( bv_1_0_n53 )  ;
assign n10277 =  ( wr_addr ) == ( bv_8_43_n155 )  ;
assign n10278 =  ( n10276 ) & (n10277 )  ;
assign n10279 =  ( n10278 ) & (wr )  ;
assign n10280 =  ( n10279 ) ? ( n5298 ) : ( iram_43 ) ;
assign n10281 = wr_addr[7:7] ;
assign n10282 =  ( n10281 ) == ( bv_1_0_n53 )  ;
assign n10283 =  ( wr_addr ) == ( bv_8_43_n155 )  ;
assign n10284 =  ( n10282 ) & (n10283 )  ;
assign n10285 =  ( n10284 ) & (wr )  ;
assign n10286 =  ( n10285 ) ? ( n5325 ) : ( iram_43 ) ;
assign n10287 = wr_addr[7:7] ;
assign n10288 =  ( n10287 ) == ( bv_1_0_n53 )  ;
assign n10289 =  ( wr_addr ) == ( bv_8_44_n157 )  ;
assign n10290 =  ( n10288 ) & (n10289 )  ;
assign n10291 =  ( n10290 ) & (wr )  ;
assign n10292 =  ( n10291 ) ? ( n4782 ) : ( iram_44 ) ;
assign n10293 = wr_addr[7:7] ;
assign n10294 =  ( n10293 ) == ( bv_1_0_n53 )  ;
assign n10295 =  ( wr_addr ) == ( bv_8_44_n157 )  ;
assign n10296 =  ( n10294 ) & (n10295 )  ;
assign n10297 =  ( n10296 ) & (wr )  ;
assign n10298 =  ( n10297 ) ? ( n4841 ) : ( iram_44 ) ;
assign n10299 = wr_addr[7:7] ;
assign n10300 =  ( n10299 ) == ( bv_1_0_n53 )  ;
assign n10301 =  ( wr_addr ) == ( bv_8_44_n157 )  ;
assign n10302 =  ( n10300 ) & (n10301 )  ;
assign n10303 =  ( n10302 ) & (wr )  ;
assign n10304 =  ( n10303 ) ? ( n5449 ) : ( iram_44 ) ;
assign n10305 = wr_addr[7:7] ;
assign n10306 =  ( n10305 ) == ( bv_1_0_n53 )  ;
assign n10307 =  ( wr_addr ) == ( bv_8_44_n157 )  ;
assign n10308 =  ( n10306 ) & (n10307 )  ;
assign n10309 =  ( n10308 ) & (wr )  ;
assign n10310 =  ( n10309 ) ? ( n4906 ) : ( iram_44 ) ;
assign n10311 = wr_addr[7:7] ;
assign n10312 =  ( n10311 ) == ( bv_1_0_n53 )  ;
assign n10313 =  ( wr_addr ) == ( bv_8_44_n157 )  ;
assign n10314 =  ( n10312 ) & (n10313 )  ;
assign n10315 =  ( n10314 ) & (wr )  ;
assign n10316 =  ( n10315 ) ? ( n5485 ) : ( iram_44 ) ;
assign n10317 = wr_addr[7:7] ;
assign n10318 =  ( n10317 ) == ( bv_1_0_n53 )  ;
assign n10319 =  ( wr_addr ) == ( bv_8_44_n157 )  ;
assign n10320 =  ( n10318 ) & (n10319 )  ;
assign n10321 =  ( n10320 ) & (wr )  ;
assign n10322 =  ( n10321 ) ? ( n5512 ) : ( iram_44 ) ;
assign n10323 = wr_addr[7:7] ;
assign n10324 =  ( n10323 ) == ( bv_1_0_n53 )  ;
assign n10325 =  ( wr_addr ) == ( bv_8_44_n157 )  ;
assign n10326 =  ( n10324 ) & (n10325 )  ;
assign n10327 =  ( n10326 ) & (wr )  ;
assign n10328 =  ( n10327 ) ? ( bv_8_0_n69 ) : ( iram_44 ) ;
assign n10329 = wr_addr[7:7] ;
assign n10330 =  ( n10329 ) == ( bv_1_0_n53 )  ;
assign n10331 =  ( wr_addr ) == ( bv_8_44_n157 )  ;
assign n10332 =  ( n10330 ) & (n10331 )  ;
assign n10333 =  ( n10332 ) & (wr )  ;
assign n10334 =  ( n10333 ) ? ( n5071 ) : ( iram_44 ) ;
assign n10335 = wr_addr[7:7] ;
assign n10336 =  ( n10335 ) == ( bv_1_0_n53 )  ;
assign n10337 =  ( wr_addr ) == ( bv_8_44_n157 )  ;
assign n10338 =  ( n10336 ) & (n10337 )  ;
assign n10339 =  ( n10338 ) & (wr )  ;
assign n10340 =  ( n10339 ) ? ( n5096 ) : ( iram_44 ) ;
assign n10341 = wr_addr[7:7] ;
assign n10342 =  ( n10341 ) == ( bv_1_0_n53 )  ;
assign n10343 =  ( wr_addr ) == ( bv_8_44_n157 )  ;
assign n10344 =  ( n10342 ) & (n10343 )  ;
assign n10345 =  ( n10344 ) & (wr )  ;
assign n10346 =  ( n10345 ) ? ( n5123 ) : ( iram_44 ) ;
assign n10347 = wr_addr[7:7] ;
assign n10348 =  ( n10347 ) == ( bv_1_0_n53 )  ;
assign n10349 =  ( wr_addr ) == ( bv_8_44_n157 )  ;
assign n10350 =  ( n10348 ) & (n10349 )  ;
assign n10351 =  ( n10350 ) & (wr )  ;
assign n10352 =  ( n10351 ) ? ( n5165 ) : ( iram_44 ) ;
assign n10353 = wr_addr[7:7] ;
assign n10354 =  ( n10353 ) == ( bv_1_0_n53 )  ;
assign n10355 =  ( wr_addr ) == ( bv_8_44_n157 )  ;
assign n10356 =  ( n10354 ) & (n10355 )  ;
assign n10357 =  ( n10356 ) & (wr )  ;
assign n10358 =  ( n10357 ) ? ( n5204 ) : ( iram_44 ) ;
assign n10359 = wr_addr[7:7] ;
assign n10360 =  ( n10359 ) == ( bv_1_0_n53 )  ;
assign n10361 =  ( wr_addr ) == ( bv_8_44_n157 )  ;
assign n10362 =  ( n10360 ) & (n10361 )  ;
assign n10363 =  ( n10362 ) & (wr )  ;
assign n10364 =  ( n10363 ) ? ( n5262 ) : ( iram_44 ) ;
assign n10365 = wr_addr[7:7] ;
assign n10366 =  ( n10365 ) == ( bv_1_0_n53 )  ;
assign n10367 =  ( wr_addr ) == ( bv_8_44_n157 )  ;
assign n10368 =  ( n10366 ) & (n10367 )  ;
assign n10369 =  ( n10368 ) & (wr )  ;
assign n10370 =  ( n10369 ) ? ( n5298 ) : ( iram_44 ) ;
assign n10371 = wr_addr[7:7] ;
assign n10372 =  ( n10371 ) == ( bv_1_0_n53 )  ;
assign n10373 =  ( wr_addr ) == ( bv_8_44_n157 )  ;
assign n10374 =  ( n10372 ) & (n10373 )  ;
assign n10375 =  ( n10374 ) & (wr )  ;
assign n10376 =  ( n10375 ) ? ( n5325 ) : ( iram_44 ) ;
assign n10377 = wr_addr[7:7] ;
assign n10378 =  ( n10377 ) == ( bv_1_0_n53 )  ;
assign n10379 =  ( wr_addr ) == ( bv_8_45_n159 )  ;
assign n10380 =  ( n10378 ) & (n10379 )  ;
assign n10381 =  ( n10380 ) & (wr )  ;
assign n10382 =  ( n10381 ) ? ( n4782 ) : ( iram_45 ) ;
assign n10383 = wr_addr[7:7] ;
assign n10384 =  ( n10383 ) == ( bv_1_0_n53 )  ;
assign n10385 =  ( wr_addr ) == ( bv_8_45_n159 )  ;
assign n10386 =  ( n10384 ) & (n10385 )  ;
assign n10387 =  ( n10386 ) & (wr )  ;
assign n10388 =  ( n10387 ) ? ( n4841 ) : ( iram_45 ) ;
assign n10389 = wr_addr[7:7] ;
assign n10390 =  ( n10389 ) == ( bv_1_0_n53 )  ;
assign n10391 =  ( wr_addr ) == ( bv_8_45_n159 )  ;
assign n10392 =  ( n10390 ) & (n10391 )  ;
assign n10393 =  ( n10392 ) & (wr )  ;
assign n10394 =  ( n10393 ) ? ( n5449 ) : ( iram_45 ) ;
assign n10395 = wr_addr[7:7] ;
assign n10396 =  ( n10395 ) == ( bv_1_0_n53 )  ;
assign n10397 =  ( wr_addr ) == ( bv_8_45_n159 )  ;
assign n10398 =  ( n10396 ) & (n10397 )  ;
assign n10399 =  ( n10398 ) & (wr )  ;
assign n10400 =  ( n10399 ) ? ( n4906 ) : ( iram_45 ) ;
assign n10401 = wr_addr[7:7] ;
assign n10402 =  ( n10401 ) == ( bv_1_0_n53 )  ;
assign n10403 =  ( wr_addr ) == ( bv_8_45_n159 )  ;
assign n10404 =  ( n10402 ) & (n10403 )  ;
assign n10405 =  ( n10404 ) & (wr )  ;
assign n10406 =  ( n10405 ) ? ( n5485 ) : ( iram_45 ) ;
assign n10407 = wr_addr[7:7] ;
assign n10408 =  ( n10407 ) == ( bv_1_0_n53 )  ;
assign n10409 =  ( wr_addr ) == ( bv_8_45_n159 )  ;
assign n10410 =  ( n10408 ) & (n10409 )  ;
assign n10411 =  ( n10410 ) & (wr )  ;
assign n10412 =  ( n10411 ) ? ( n5512 ) : ( iram_45 ) ;
assign n10413 = wr_addr[7:7] ;
assign n10414 =  ( n10413 ) == ( bv_1_0_n53 )  ;
assign n10415 =  ( wr_addr ) == ( bv_8_45_n159 )  ;
assign n10416 =  ( n10414 ) & (n10415 )  ;
assign n10417 =  ( n10416 ) & (wr )  ;
assign n10418 =  ( n10417 ) ? ( bv_8_0_n69 ) : ( iram_45 ) ;
assign n10419 = wr_addr[7:7] ;
assign n10420 =  ( n10419 ) == ( bv_1_0_n53 )  ;
assign n10421 =  ( wr_addr ) == ( bv_8_45_n159 )  ;
assign n10422 =  ( n10420 ) & (n10421 )  ;
assign n10423 =  ( n10422 ) & (wr )  ;
assign n10424 =  ( n10423 ) ? ( n5071 ) : ( iram_45 ) ;
assign n10425 = wr_addr[7:7] ;
assign n10426 =  ( n10425 ) == ( bv_1_0_n53 )  ;
assign n10427 =  ( wr_addr ) == ( bv_8_45_n159 )  ;
assign n10428 =  ( n10426 ) & (n10427 )  ;
assign n10429 =  ( n10428 ) & (wr )  ;
assign n10430 =  ( n10429 ) ? ( n5096 ) : ( iram_45 ) ;
assign n10431 = wr_addr[7:7] ;
assign n10432 =  ( n10431 ) == ( bv_1_0_n53 )  ;
assign n10433 =  ( wr_addr ) == ( bv_8_45_n159 )  ;
assign n10434 =  ( n10432 ) & (n10433 )  ;
assign n10435 =  ( n10434 ) & (wr )  ;
assign n10436 =  ( n10435 ) ? ( n5123 ) : ( iram_45 ) ;
assign n10437 = wr_addr[7:7] ;
assign n10438 =  ( n10437 ) == ( bv_1_0_n53 )  ;
assign n10439 =  ( wr_addr ) == ( bv_8_45_n159 )  ;
assign n10440 =  ( n10438 ) & (n10439 )  ;
assign n10441 =  ( n10440 ) & (wr )  ;
assign n10442 =  ( n10441 ) ? ( n5165 ) : ( iram_45 ) ;
assign n10443 = wr_addr[7:7] ;
assign n10444 =  ( n10443 ) == ( bv_1_0_n53 )  ;
assign n10445 =  ( wr_addr ) == ( bv_8_45_n159 )  ;
assign n10446 =  ( n10444 ) & (n10445 )  ;
assign n10447 =  ( n10446 ) & (wr )  ;
assign n10448 =  ( n10447 ) ? ( n5204 ) : ( iram_45 ) ;
assign n10449 = wr_addr[7:7] ;
assign n10450 =  ( n10449 ) == ( bv_1_0_n53 )  ;
assign n10451 =  ( wr_addr ) == ( bv_8_45_n159 )  ;
assign n10452 =  ( n10450 ) & (n10451 )  ;
assign n10453 =  ( n10452 ) & (wr )  ;
assign n10454 =  ( n10453 ) ? ( n5262 ) : ( iram_45 ) ;
assign n10455 = wr_addr[7:7] ;
assign n10456 =  ( n10455 ) == ( bv_1_0_n53 )  ;
assign n10457 =  ( wr_addr ) == ( bv_8_45_n159 )  ;
assign n10458 =  ( n10456 ) & (n10457 )  ;
assign n10459 =  ( n10458 ) & (wr )  ;
assign n10460 =  ( n10459 ) ? ( n5298 ) : ( iram_45 ) ;
assign n10461 = wr_addr[7:7] ;
assign n10462 =  ( n10461 ) == ( bv_1_0_n53 )  ;
assign n10463 =  ( wr_addr ) == ( bv_8_45_n159 )  ;
assign n10464 =  ( n10462 ) & (n10463 )  ;
assign n10465 =  ( n10464 ) & (wr )  ;
assign n10466 =  ( n10465 ) ? ( n5325 ) : ( iram_45 ) ;
assign n10467 = wr_addr[7:7] ;
assign n10468 =  ( n10467 ) == ( bv_1_0_n53 )  ;
assign n10469 =  ( wr_addr ) == ( bv_8_46_n161 )  ;
assign n10470 =  ( n10468 ) & (n10469 )  ;
assign n10471 =  ( n10470 ) & (wr )  ;
assign n10472 =  ( n10471 ) ? ( n4782 ) : ( iram_46 ) ;
assign n10473 = wr_addr[7:7] ;
assign n10474 =  ( n10473 ) == ( bv_1_0_n53 )  ;
assign n10475 =  ( wr_addr ) == ( bv_8_46_n161 )  ;
assign n10476 =  ( n10474 ) & (n10475 )  ;
assign n10477 =  ( n10476 ) & (wr )  ;
assign n10478 =  ( n10477 ) ? ( n4841 ) : ( iram_46 ) ;
assign n10479 = wr_addr[7:7] ;
assign n10480 =  ( n10479 ) == ( bv_1_0_n53 )  ;
assign n10481 =  ( wr_addr ) == ( bv_8_46_n161 )  ;
assign n10482 =  ( n10480 ) & (n10481 )  ;
assign n10483 =  ( n10482 ) & (wr )  ;
assign n10484 =  ( n10483 ) ? ( n5449 ) : ( iram_46 ) ;
assign n10485 = wr_addr[7:7] ;
assign n10486 =  ( n10485 ) == ( bv_1_0_n53 )  ;
assign n10487 =  ( wr_addr ) == ( bv_8_46_n161 )  ;
assign n10488 =  ( n10486 ) & (n10487 )  ;
assign n10489 =  ( n10488 ) & (wr )  ;
assign n10490 =  ( n10489 ) ? ( n4906 ) : ( iram_46 ) ;
assign n10491 = wr_addr[7:7] ;
assign n10492 =  ( n10491 ) == ( bv_1_0_n53 )  ;
assign n10493 =  ( wr_addr ) == ( bv_8_46_n161 )  ;
assign n10494 =  ( n10492 ) & (n10493 )  ;
assign n10495 =  ( n10494 ) & (wr )  ;
assign n10496 =  ( n10495 ) ? ( n5485 ) : ( iram_46 ) ;
assign n10497 = wr_addr[7:7] ;
assign n10498 =  ( n10497 ) == ( bv_1_0_n53 )  ;
assign n10499 =  ( wr_addr ) == ( bv_8_46_n161 )  ;
assign n10500 =  ( n10498 ) & (n10499 )  ;
assign n10501 =  ( n10500 ) & (wr )  ;
assign n10502 =  ( n10501 ) ? ( n5512 ) : ( iram_46 ) ;
assign n10503 = wr_addr[7:7] ;
assign n10504 =  ( n10503 ) == ( bv_1_0_n53 )  ;
assign n10505 =  ( wr_addr ) == ( bv_8_46_n161 )  ;
assign n10506 =  ( n10504 ) & (n10505 )  ;
assign n10507 =  ( n10506 ) & (wr )  ;
assign n10508 =  ( n10507 ) ? ( bv_8_0_n69 ) : ( iram_46 ) ;
assign n10509 = wr_addr[7:7] ;
assign n10510 =  ( n10509 ) == ( bv_1_0_n53 )  ;
assign n10511 =  ( wr_addr ) == ( bv_8_46_n161 )  ;
assign n10512 =  ( n10510 ) & (n10511 )  ;
assign n10513 =  ( n10512 ) & (wr )  ;
assign n10514 =  ( n10513 ) ? ( n5071 ) : ( iram_46 ) ;
assign n10515 = wr_addr[7:7] ;
assign n10516 =  ( n10515 ) == ( bv_1_0_n53 )  ;
assign n10517 =  ( wr_addr ) == ( bv_8_46_n161 )  ;
assign n10518 =  ( n10516 ) & (n10517 )  ;
assign n10519 =  ( n10518 ) & (wr )  ;
assign n10520 =  ( n10519 ) ? ( n5096 ) : ( iram_46 ) ;
assign n10521 = wr_addr[7:7] ;
assign n10522 =  ( n10521 ) == ( bv_1_0_n53 )  ;
assign n10523 =  ( wr_addr ) == ( bv_8_46_n161 )  ;
assign n10524 =  ( n10522 ) & (n10523 )  ;
assign n10525 =  ( n10524 ) & (wr )  ;
assign n10526 =  ( n10525 ) ? ( n5123 ) : ( iram_46 ) ;
assign n10527 = wr_addr[7:7] ;
assign n10528 =  ( n10527 ) == ( bv_1_0_n53 )  ;
assign n10529 =  ( wr_addr ) == ( bv_8_46_n161 )  ;
assign n10530 =  ( n10528 ) & (n10529 )  ;
assign n10531 =  ( n10530 ) & (wr )  ;
assign n10532 =  ( n10531 ) ? ( n5165 ) : ( iram_46 ) ;
assign n10533 = wr_addr[7:7] ;
assign n10534 =  ( n10533 ) == ( bv_1_0_n53 )  ;
assign n10535 =  ( wr_addr ) == ( bv_8_46_n161 )  ;
assign n10536 =  ( n10534 ) & (n10535 )  ;
assign n10537 =  ( n10536 ) & (wr )  ;
assign n10538 =  ( n10537 ) ? ( n5204 ) : ( iram_46 ) ;
assign n10539 = wr_addr[7:7] ;
assign n10540 =  ( n10539 ) == ( bv_1_0_n53 )  ;
assign n10541 =  ( wr_addr ) == ( bv_8_46_n161 )  ;
assign n10542 =  ( n10540 ) & (n10541 )  ;
assign n10543 =  ( n10542 ) & (wr )  ;
assign n10544 =  ( n10543 ) ? ( n5262 ) : ( iram_46 ) ;
assign n10545 = wr_addr[7:7] ;
assign n10546 =  ( n10545 ) == ( bv_1_0_n53 )  ;
assign n10547 =  ( wr_addr ) == ( bv_8_46_n161 )  ;
assign n10548 =  ( n10546 ) & (n10547 )  ;
assign n10549 =  ( n10548 ) & (wr )  ;
assign n10550 =  ( n10549 ) ? ( n5298 ) : ( iram_46 ) ;
assign n10551 = wr_addr[7:7] ;
assign n10552 =  ( n10551 ) == ( bv_1_0_n53 )  ;
assign n10553 =  ( wr_addr ) == ( bv_8_46_n161 )  ;
assign n10554 =  ( n10552 ) & (n10553 )  ;
assign n10555 =  ( n10554 ) & (wr )  ;
assign n10556 =  ( n10555 ) ? ( n5325 ) : ( iram_46 ) ;
assign n10557 = wr_addr[7:7] ;
assign n10558 =  ( n10557 ) == ( bv_1_0_n53 )  ;
assign n10559 =  ( wr_addr ) == ( bv_8_47_n163 )  ;
assign n10560 =  ( n10558 ) & (n10559 )  ;
assign n10561 =  ( n10560 ) & (wr )  ;
assign n10562 =  ( n10561 ) ? ( n4782 ) : ( iram_47 ) ;
assign n10563 = wr_addr[7:7] ;
assign n10564 =  ( n10563 ) == ( bv_1_0_n53 )  ;
assign n10565 =  ( wr_addr ) == ( bv_8_47_n163 )  ;
assign n10566 =  ( n10564 ) & (n10565 )  ;
assign n10567 =  ( n10566 ) & (wr )  ;
assign n10568 =  ( n10567 ) ? ( n4841 ) : ( iram_47 ) ;
assign n10569 = wr_addr[7:7] ;
assign n10570 =  ( n10569 ) == ( bv_1_0_n53 )  ;
assign n10571 =  ( wr_addr ) == ( bv_8_47_n163 )  ;
assign n10572 =  ( n10570 ) & (n10571 )  ;
assign n10573 =  ( n10572 ) & (wr )  ;
assign n10574 =  ( n10573 ) ? ( n5449 ) : ( iram_47 ) ;
assign n10575 = wr_addr[7:7] ;
assign n10576 =  ( n10575 ) == ( bv_1_0_n53 )  ;
assign n10577 =  ( wr_addr ) == ( bv_8_47_n163 )  ;
assign n10578 =  ( n10576 ) & (n10577 )  ;
assign n10579 =  ( n10578 ) & (wr )  ;
assign n10580 =  ( n10579 ) ? ( n4906 ) : ( iram_47 ) ;
assign n10581 = wr_addr[7:7] ;
assign n10582 =  ( n10581 ) == ( bv_1_0_n53 )  ;
assign n10583 =  ( wr_addr ) == ( bv_8_47_n163 )  ;
assign n10584 =  ( n10582 ) & (n10583 )  ;
assign n10585 =  ( n10584 ) & (wr )  ;
assign n10586 =  ( n10585 ) ? ( n5485 ) : ( iram_47 ) ;
assign n10587 = wr_addr[7:7] ;
assign n10588 =  ( n10587 ) == ( bv_1_0_n53 )  ;
assign n10589 =  ( wr_addr ) == ( bv_8_47_n163 )  ;
assign n10590 =  ( n10588 ) & (n10589 )  ;
assign n10591 =  ( n10590 ) & (wr )  ;
assign n10592 =  ( n10591 ) ? ( n5512 ) : ( iram_47 ) ;
assign n10593 = wr_addr[7:7] ;
assign n10594 =  ( n10593 ) == ( bv_1_0_n53 )  ;
assign n10595 =  ( wr_addr ) == ( bv_8_47_n163 )  ;
assign n10596 =  ( n10594 ) & (n10595 )  ;
assign n10597 =  ( n10596 ) & (wr )  ;
assign n10598 =  ( n10597 ) ? ( bv_8_0_n69 ) : ( iram_47 ) ;
assign n10599 = wr_addr[7:7] ;
assign n10600 =  ( n10599 ) == ( bv_1_0_n53 )  ;
assign n10601 =  ( wr_addr ) == ( bv_8_47_n163 )  ;
assign n10602 =  ( n10600 ) & (n10601 )  ;
assign n10603 =  ( n10602 ) & (wr )  ;
assign n10604 =  ( n10603 ) ? ( n5071 ) : ( iram_47 ) ;
assign n10605 = wr_addr[7:7] ;
assign n10606 =  ( n10605 ) == ( bv_1_0_n53 )  ;
assign n10607 =  ( wr_addr ) == ( bv_8_47_n163 )  ;
assign n10608 =  ( n10606 ) & (n10607 )  ;
assign n10609 =  ( n10608 ) & (wr )  ;
assign n10610 =  ( n10609 ) ? ( n5096 ) : ( iram_47 ) ;
assign n10611 = wr_addr[7:7] ;
assign n10612 =  ( n10611 ) == ( bv_1_0_n53 )  ;
assign n10613 =  ( wr_addr ) == ( bv_8_47_n163 )  ;
assign n10614 =  ( n10612 ) & (n10613 )  ;
assign n10615 =  ( n10614 ) & (wr )  ;
assign n10616 =  ( n10615 ) ? ( n5123 ) : ( iram_47 ) ;
assign n10617 = wr_addr[7:7] ;
assign n10618 =  ( n10617 ) == ( bv_1_0_n53 )  ;
assign n10619 =  ( wr_addr ) == ( bv_8_47_n163 )  ;
assign n10620 =  ( n10618 ) & (n10619 )  ;
assign n10621 =  ( n10620 ) & (wr )  ;
assign n10622 =  ( n10621 ) ? ( n5165 ) : ( iram_47 ) ;
assign n10623 = wr_addr[7:7] ;
assign n10624 =  ( n10623 ) == ( bv_1_0_n53 )  ;
assign n10625 =  ( wr_addr ) == ( bv_8_47_n163 )  ;
assign n10626 =  ( n10624 ) & (n10625 )  ;
assign n10627 =  ( n10626 ) & (wr )  ;
assign n10628 =  ( n10627 ) ? ( n5204 ) : ( iram_47 ) ;
assign n10629 = wr_addr[7:7] ;
assign n10630 =  ( n10629 ) == ( bv_1_0_n53 )  ;
assign n10631 =  ( wr_addr ) == ( bv_8_47_n163 )  ;
assign n10632 =  ( n10630 ) & (n10631 )  ;
assign n10633 =  ( n10632 ) & (wr )  ;
assign n10634 =  ( n10633 ) ? ( n5262 ) : ( iram_47 ) ;
assign n10635 = wr_addr[7:7] ;
assign n10636 =  ( n10635 ) == ( bv_1_0_n53 )  ;
assign n10637 =  ( wr_addr ) == ( bv_8_47_n163 )  ;
assign n10638 =  ( n10636 ) & (n10637 )  ;
assign n10639 =  ( n10638 ) & (wr )  ;
assign n10640 =  ( n10639 ) ? ( n5298 ) : ( iram_47 ) ;
assign n10641 = wr_addr[7:7] ;
assign n10642 =  ( n10641 ) == ( bv_1_0_n53 )  ;
assign n10643 =  ( wr_addr ) == ( bv_8_47_n163 )  ;
assign n10644 =  ( n10642 ) & (n10643 )  ;
assign n10645 =  ( n10644 ) & (wr )  ;
assign n10646 =  ( n10645 ) ? ( n5325 ) : ( iram_47 ) ;
assign n10647 = wr_addr[7:7] ;
assign n10648 =  ( n10647 ) == ( bv_1_0_n53 )  ;
assign n10649 =  ( wr_addr ) == ( bv_8_48_n165 )  ;
assign n10650 =  ( n10648 ) & (n10649 )  ;
assign n10651 =  ( n10650 ) & (wr )  ;
assign n10652 =  ( n10651 ) ? ( n4782 ) : ( iram_48 ) ;
assign n10653 = wr_addr[7:7] ;
assign n10654 =  ( n10653 ) == ( bv_1_0_n53 )  ;
assign n10655 =  ( wr_addr ) == ( bv_8_48_n165 )  ;
assign n10656 =  ( n10654 ) & (n10655 )  ;
assign n10657 =  ( n10656 ) & (wr )  ;
assign n10658 =  ( n10657 ) ? ( n4841 ) : ( iram_48 ) ;
assign n10659 = wr_addr[7:7] ;
assign n10660 =  ( n10659 ) == ( bv_1_0_n53 )  ;
assign n10661 =  ( wr_addr ) == ( bv_8_48_n165 )  ;
assign n10662 =  ( n10660 ) & (n10661 )  ;
assign n10663 =  ( n10662 ) & (wr )  ;
assign n10664 =  ( n10663 ) ? ( n5449 ) : ( iram_48 ) ;
assign n10665 = wr_addr[7:7] ;
assign n10666 =  ( n10665 ) == ( bv_1_0_n53 )  ;
assign n10667 =  ( wr_addr ) == ( bv_8_48_n165 )  ;
assign n10668 =  ( n10666 ) & (n10667 )  ;
assign n10669 =  ( n10668 ) & (wr )  ;
assign n10670 =  ( n10669 ) ? ( n4906 ) : ( iram_48 ) ;
assign n10671 = wr_addr[7:7] ;
assign n10672 =  ( n10671 ) == ( bv_1_0_n53 )  ;
assign n10673 =  ( wr_addr ) == ( bv_8_48_n165 )  ;
assign n10674 =  ( n10672 ) & (n10673 )  ;
assign n10675 =  ( n10674 ) & (wr )  ;
assign n10676 =  ( n10675 ) ? ( n5485 ) : ( iram_48 ) ;
assign n10677 = wr_addr[7:7] ;
assign n10678 =  ( n10677 ) == ( bv_1_0_n53 )  ;
assign n10679 =  ( wr_addr ) == ( bv_8_48_n165 )  ;
assign n10680 =  ( n10678 ) & (n10679 )  ;
assign n10681 =  ( n10680 ) & (wr )  ;
assign n10682 =  ( n10681 ) ? ( n5512 ) : ( iram_48 ) ;
assign n10683 = wr_addr[7:7] ;
assign n10684 =  ( n10683 ) == ( bv_1_0_n53 )  ;
assign n10685 =  ( wr_addr ) == ( bv_8_48_n165 )  ;
assign n10686 =  ( n10684 ) & (n10685 )  ;
assign n10687 =  ( n10686 ) & (wr )  ;
assign n10688 =  ( n10687 ) ? ( bv_8_0_n69 ) : ( iram_48 ) ;
assign n10689 = wr_addr[7:7] ;
assign n10690 =  ( n10689 ) == ( bv_1_0_n53 )  ;
assign n10691 =  ( wr_addr ) == ( bv_8_48_n165 )  ;
assign n10692 =  ( n10690 ) & (n10691 )  ;
assign n10693 =  ( n10692 ) & (wr )  ;
assign n10694 =  ( n10693 ) ? ( n5071 ) : ( iram_48 ) ;
assign n10695 = wr_addr[7:7] ;
assign n10696 =  ( n10695 ) == ( bv_1_0_n53 )  ;
assign n10697 =  ( wr_addr ) == ( bv_8_48_n165 )  ;
assign n10698 =  ( n10696 ) & (n10697 )  ;
assign n10699 =  ( n10698 ) & (wr )  ;
assign n10700 =  ( n10699 ) ? ( n5096 ) : ( iram_48 ) ;
assign n10701 = wr_addr[7:7] ;
assign n10702 =  ( n10701 ) == ( bv_1_0_n53 )  ;
assign n10703 =  ( wr_addr ) == ( bv_8_48_n165 )  ;
assign n10704 =  ( n10702 ) & (n10703 )  ;
assign n10705 =  ( n10704 ) & (wr )  ;
assign n10706 =  ( n10705 ) ? ( n5123 ) : ( iram_48 ) ;
assign n10707 = wr_addr[7:7] ;
assign n10708 =  ( n10707 ) == ( bv_1_0_n53 )  ;
assign n10709 =  ( wr_addr ) == ( bv_8_48_n165 )  ;
assign n10710 =  ( n10708 ) & (n10709 )  ;
assign n10711 =  ( n10710 ) & (wr )  ;
assign n10712 =  ( n10711 ) ? ( n5165 ) : ( iram_48 ) ;
assign n10713 = wr_addr[7:7] ;
assign n10714 =  ( n10713 ) == ( bv_1_0_n53 )  ;
assign n10715 =  ( wr_addr ) == ( bv_8_48_n165 )  ;
assign n10716 =  ( n10714 ) & (n10715 )  ;
assign n10717 =  ( n10716 ) & (wr )  ;
assign n10718 =  ( n10717 ) ? ( n5204 ) : ( iram_48 ) ;
assign n10719 = wr_addr[7:7] ;
assign n10720 =  ( n10719 ) == ( bv_1_0_n53 )  ;
assign n10721 =  ( wr_addr ) == ( bv_8_48_n165 )  ;
assign n10722 =  ( n10720 ) & (n10721 )  ;
assign n10723 =  ( n10722 ) & (wr )  ;
assign n10724 =  ( n10723 ) ? ( n5262 ) : ( iram_48 ) ;
assign n10725 = wr_addr[7:7] ;
assign n10726 =  ( n10725 ) == ( bv_1_0_n53 )  ;
assign n10727 =  ( wr_addr ) == ( bv_8_48_n165 )  ;
assign n10728 =  ( n10726 ) & (n10727 )  ;
assign n10729 =  ( n10728 ) & (wr )  ;
assign n10730 =  ( n10729 ) ? ( n5298 ) : ( iram_48 ) ;
assign n10731 = wr_addr[7:7] ;
assign n10732 =  ( n10731 ) == ( bv_1_0_n53 )  ;
assign n10733 =  ( wr_addr ) == ( bv_8_48_n165 )  ;
assign n10734 =  ( n10732 ) & (n10733 )  ;
assign n10735 =  ( n10734 ) & (wr )  ;
assign n10736 =  ( n10735 ) ? ( n5325 ) : ( iram_48 ) ;
assign n10737 = wr_addr[7:7] ;
assign n10738 =  ( n10737 ) == ( bv_1_0_n53 )  ;
assign n10739 =  ( wr_addr ) == ( bv_8_49_n167 )  ;
assign n10740 =  ( n10738 ) & (n10739 )  ;
assign n10741 =  ( n10740 ) & (wr )  ;
assign n10742 =  ( n10741 ) ? ( n4782 ) : ( iram_49 ) ;
assign n10743 = wr_addr[7:7] ;
assign n10744 =  ( n10743 ) == ( bv_1_0_n53 )  ;
assign n10745 =  ( wr_addr ) == ( bv_8_49_n167 )  ;
assign n10746 =  ( n10744 ) & (n10745 )  ;
assign n10747 =  ( n10746 ) & (wr )  ;
assign n10748 =  ( n10747 ) ? ( n4841 ) : ( iram_49 ) ;
assign n10749 = wr_addr[7:7] ;
assign n10750 =  ( n10749 ) == ( bv_1_0_n53 )  ;
assign n10751 =  ( wr_addr ) == ( bv_8_49_n167 )  ;
assign n10752 =  ( n10750 ) & (n10751 )  ;
assign n10753 =  ( n10752 ) & (wr )  ;
assign n10754 =  ( n10753 ) ? ( n5449 ) : ( iram_49 ) ;
assign n10755 = wr_addr[7:7] ;
assign n10756 =  ( n10755 ) == ( bv_1_0_n53 )  ;
assign n10757 =  ( wr_addr ) == ( bv_8_49_n167 )  ;
assign n10758 =  ( n10756 ) & (n10757 )  ;
assign n10759 =  ( n10758 ) & (wr )  ;
assign n10760 =  ( n10759 ) ? ( n4906 ) : ( iram_49 ) ;
assign n10761 = wr_addr[7:7] ;
assign n10762 =  ( n10761 ) == ( bv_1_0_n53 )  ;
assign n10763 =  ( wr_addr ) == ( bv_8_49_n167 )  ;
assign n10764 =  ( n10762 ) & (n10763 )  ;
assign n10765 =  ( n10764 ) & (wr )  ;
assign n10766 =  ( n10765 ) ? ( n5485 ) : ( iram_49 ) ;
assign n10767 = wr_addr[7:7] ;
assign n10768 =  ( n10767 ) == ( bv_1_0_n53 )  ;
assign n10769 =  ( wr_addr ) == ( bv_8_49_n167 )  ;
assign n10770 =  ( n10768 ) & (n10769 )  ;
assign n10771 =  ( n10770 ) & (wr )  ;
assign n10772 =  ( n10771 ) ? ( n5512 ) : ( iram_49 ) ;
assign n10773 = wr_addr[7:7] ;
assign n10774 =  ( n10773 ) == ( bv_1_0_n53 )  ;
assign n10775 =  ( wr_addr ) == ( bv_8_49_n167 )  ;
assign n10776 =  ( n10774 ) & (n10775 )  ;
assign n10777 =  ( n10776 ) & (wr )  ;
assign n10778 =  ( n10777 ) ? ( bv_8_0_n69 ) : ( iram_49 ) ;
assign n10779 = wr_addr[7:7] ;
assign n10780 =  ( n10779 ) == ( bv_1_0_n53 )  ;
assign n10781 =  ( wr_addr ) == ( bv_8_49_n167 )  ;
assign n10782 =  ( n10780 ) & (n10781 )  ;
assign n10783 =  ( n10782 ) & (wr )  ;
assign n10784 =  ( n10783 ) ? ( n5071 ) : ( iram_49 ) ;
assign n10785 = wr_addr[7:7] ;
assign n10786 =  ( n10785 ) == ( bv_1_0_n53 )  ;
assign n10787 =  ( wr_addr ) == ( bv_8_49_n167 )  ;
assign n10788 =  ( n10786 ) & (n10787 )  ;
assign n10789 =  ( n10788 ) & (wr )  ;
assign n10790 =  ( n10789 ) ? ( n5096 ) : ( iram_49 ) ;
assign n10791 = wr_addr[7:7] ;
assign n10792 =  ( n10791 ) == ( bv_1_0_n53 )  ;
assign n10793 =  ( wr_addr ) == ( bv_8_49_n167 )  ;
assign n10794 =  ( n10792 ) & (n10793 )  ;
assign n10795 =  ( n10794 ) & (wr )  ;
assign n10796 =  ( n10795 ) ? ( n5123 ) : ( iram_49 ) ;
assign n10797 = wr_addr[7:7] ;
assign n10798 =  ( n10797 ) == ( bv_1_0_n53 )  ;
assign n10799 =  ( wr_addr ) == ( bv_8_49_n167 )  ;
assign n10800 =  ( n10798 ) & (n10799 )  ;
assign n10801 =  ( n10800 ) & (wr )  ;
assign n10802 =  ( n10801 ) ? ( n5165 ) : ( iram_49 ) ;
assign n10803 = wr_addr[7:7] ;
assign n10804 =  ( n10803 ) == ( bv_1_0_n53 )  ;
assign n10805 =  ( wr_addr ) == ( bv_8_49_n167 )  ;
assign n10806 =  ( n10804 ) & (n10805 )  ;
assign n10807 =  ( n10806 ) & (wr )  ;
assign n10808 =  ( n10807 ) ? ( n5204 ) : ( iram_49 ) ;
assign n10809 = wr_addr[7:7] ;
assign n10810 =  ( n10809 ) == ( bv_1_0_n53 )  ;
assign n10811 =  ( wr_addr ) == ( bv_8_49_n167 )  ;
assign n10812 =  ( n10810 ) & (n10811 )  ;
assign n10813 =  ( n10812 ) & (wr )  ;
assign n10814 =  ( n10813 ) ? ( n5262 ) : ( iram_49 ) ;
assign n10815 = wr_addr[7:7] ;
assign n10816 =  ( n10815 ) == ( bv_1_0_n53 )  ;
assign n10817 =  ( wr_addr ) == ( bv_8_49_n167 )  ;
assign n10818 =  ( n10816 ) & (n10817 )  ;
assign n10819 =  ( n10818 ) & (wr )  ;
assign n10820 =  ( n10819 ) ? ( n5298 ) : ( iram_49 ) ;
assign n10821 = wr_addr[7:7] ;
assign n10822 =  ( n10821 ) == ( bv_1_0_n53 )  ;
assign n10823 =  ( wr_addr ) == ( bv_8_49_n167 )  ;
assign n10824 =  ( n10822 ) & (n10823 )  ;
assign n10825 =  ( n10824 ) & (wr )  ;
assign n10826 =  ( n10825 ) ? ( n5325 ) : ( iram_49 ) ;
assign n10827 = wr_addr[7:7] ;
assign n10828 =  ( n10827 ) == ( bv_1_0_n53 )  ;
assign n10829 =  ( wr_addr ) == ( bv_8_50_n169 )  ;
assign n10830 =  ( n10828 ) & (n10829 )  ;
assign n10831 =  ( n10830 ) & (wr )  ;
assign n10832 =  ( n10831 ) ? ( n4782 ) : ( iram_50 ) ;
assign n10833 = wr_addr[7:7] ;
assign n10834 =  ( n10833 ) == ( bv_1_0_n53 )  ;
assign n10835 =  ( wr_addr ) == ( bv_8_50_n169 )  ;
assign n10836 =  ( n10834 ) & (n10835 )  ;
assign n10837 =  ( n10836 ) & (wr )  ;
assign n10838 =  ( n10837 ) ? ( n4841 ) : ( iram_50 ) ;
assign n10839 = wr_addr[7:7] ;
assign n10840 =  ( n10839 ) == ( bv_1_0_n53 )  ;
assign n10841 =  ( wr_addr ) == ( bv_8_50_n169 )  ;
assign n10842 =  ( n10840 ) & (n10841 )  ;
assign n10843 =  ( n10842 ) & (wr )  ;
assign n10844 =  ( n10843 ) ? ( n5449 ) : ( iram_50 ) ;
assign n10845 = wr_addr[7:7] ;
assign n10846 =  ( n10845 ) == ( bv_1_0_n53 )  ;
assign n10847 =  ( wr_addr ) == ( bv_8_50_n169 )  ;
assign n10848 =  ( n10846 ) & (n10847 )  ;
assign n10849 =  ( n10848 ) & (wr )  ;
assign n10850 =  ( n10849 ) ? ( n4906 ) : ( iram_50 ) ;
assign n10851 = wr_addr[7:7] ;
assign n10852 =  ( n10851 ) == ( bv_1_0_n53 )  ;
assign n10853 =  ( wr_addr ) == ( bv_8_50_n169 )  ;
assign n10854 =  ( n10852 ) & (n10853 )  ;
assign n10855 =  ( n10854 ) & (wr )  ;
assign n10856 =  ( n10855 ) ? ( n5485 ) : ( iram_50 ) ;
assign n10857 = wr_addr[7:7] ;
assign n10858 =  ( n10857 ) == ( bv_1_0_n53 )  ;
assign n10859 =  ( wr_addr ) == ( bv_8_50_n169 )  ;
assign n10860 =  ( n10858 ) & (n10859 )  ;
assign n10861 =  ( n10860 ) & (wr )  ;
assign n10862 =  ( n10861 ) ? ( n5512 ) : ( iram_50 ) ;
assign n10863 = wr_addr[7:7] ;
assign n10864 =  ( n10863 ) == ( bv_1_0_n53 )  ;
assign n10865 =  ( wr_addr ) == ( bv_8_50_n169 )  ;
assign n10866 =  ( n10864 ) & (n10865 )  ;
assign n10867 =  ( n10866 ) & (wr )  ;
assign n10868 =  ( n10867 ) ? ( bv_8_0_n69 ) : ( iram_50 ) ;
assign n10869 = wr_addr[7:7] ;
assign n10870 =  ( n10869 ) == ( bv_1_0_n53 )  ;
assign n10871 =  ( wr_addr ) == ( bv_8_50_n169 )  ;
assign n10872 =  ( n10870 ) & (n10871 )  ;
assign n10873 =  ( n10872 ) & (wr )  ;
assign n10874 =  ( n10873 ) ? ( n5071 ) : ( iram_50 ) ;
assign n10875 = wr_addr[7:7] ;
assign n10876 =  ( n10875 ) == ( bv_1_0_n53 )  ;
assign n10877 =  ( wr_addr ) == ( bv_8_50_n169 )  ;
assign n10878 =  ( n10876 ) & (n10877 )  ;
assign n10879 =  ( n10878 ) & (wr )  ;
assign n10880 =  ( n10879 ) ? ( n5096 ) : ( iram_50 ) ;
assign n10881 = wr_addr[7:7] ;
assign n10882 =  ( n10881 ) == ( bv_1_0_n53 )  ;
assign n10883 =  ( wr_addr ) == ( bv_8_50_n169 )  ;
assign n10884 =  ( n10882 ) & (n10883 )  ;
assign n10885 =  ( n10884 ) & (wr )  ;
assign n10886 =  ( n10885 ) ? ( n5123 ) : ( iram_50 ) ;
assign n10887 = wr_addr[7:7] ;
assign n10888 =  ( n10887 ) == ( bv_1_0_n53 )  ;
assign n10889 =  ( wr_addr ) == ( bv_8_50_n169 )  ;
assign n10890 =  ( n10888 ) & (n10889 )  ;
assign n10891 =  ( n10890 ) & (wr )  ;
assign n10892 =  ( n10891 ) ? ( n5165 ) : ( iram_50 ) ;
assign n10893 = wr_addr[7:7] ;
assign n10894 =  ( n10893 ) == ( bv_1_0_n53 )  ;
assign n10895 =  ( wr_addr ) == ( bv_8_50_n169 )  ;
assign n10896 =  ( n10894 ) & (n10895 )  ;
assign n10897 =  ( n10896 ) & (wr )  ;
assign n10898 =  ( n10897 ) ? ( n5204 ) : ( iram_50 ) ;
assign n10899 = wr_addr[7:7] ;
assign n10900 =  ( n10899 ) == ( bv_1_0_n53 )  ;
assign n10901 =  ( wr_addr ) == ( bv_8_50_n169 )  ;
assign n10902 =  ( n10900 ) & (n10901 )  ;
assign n10903 =  ( n10902 ) & (wr )  ;
assign n10904 =  ( n10903 ) ? ( n5262 ) : ( iram_50 ) ;
assign n10905 = wr_addr[7:7] ;
assign n10906 =  ( n10905 ) == ( bv_1_0_n53 )  ;
assign n10907 =  ( wr_addr ) == ( bv_8_50_n169 )  ;
assign n10908 =  ( n10906 ) & (n10907 )  ;
assign n10909 =  ( n10908 ) & (wr )  ;
assign n10910 =  ( n10909 ) ? ( n5298 ) : ( iram_50 ) ;
assign n10911 = wr_addr[7:7] ;
assign n10912 =  ( n10911 ) == ( bv_1_0_n53 )  ;
assign n10913 =  ( wr_addr ) == ( bv_8_50_n169 )  ;
assign n10914 =  ( n10912 ) & (n10913 )  ;
assign n10915 =  ( n10914 ) & (wr )  ;
assign n10916 =  ( n10915 ) ? ( n5325 ) : ( iram_50 ) ;
assign n10917 = wr_addr[7:7] ;
assign n10918 =  ( n10917 ) == ( bv_1_0_n53 )  ;
assign n10919 =  ( wr_addr ) == ( bv_8_51_n171 )  ;
assign n10920 =  ( n10918 ) & (n10919 )  ;
assign n10921 =  ( n10920 ) & (wr )  ;
assign n10922 =  ( n10921 ) ? ( n4782 ) : ( iram_51 ) ;
assign n10923 = wr_addr[7:7] ;
assign n10924 =  ( n10923 ) == ( bv_1_0_n53 )  ;
assign n10925 =  ( wr_addr ) == ( bv_8_51_n171 )  ;
assign n10926 =  ( n10924 ) & (n10925 )  ;
assign n10927 =  ( n10926 ) & (wr )  ;
assign n10928 =  ( n10927 ) ? ( n4841 ) : ( iram_51 ) ;
assign n10929 = wr_addr[7:7] ;
assign n10930 =  ( n10929 ) == ( bv_1_0_n53 )  ;
assign n10931 =  ( wr_addr ) == ( bv_8_51_n171 )  ;
assign n10932 =  ( n10930 ) & (n10931 )  ;
assign n10933 =  ( n10932 ) & (wr )  ;
assign n10934 =  ( n10933 ) ? ( n5449 ) : ( iram_51 ) ;
assign n10935 = wr_addr[7:7] ;
assign n10936 =  ( n10935 ) == ( bv_1_0_n53 )  ;
assign n10937 =  ( wr_addr ) == ( bv_8_51_n171 )  ;
assign n10938 =  ( n10936 ) & (n10937 )  ;
assign n10939 =  ( n10938 ) & (wr )  ;
assign n10940 =  ( n10939 ) ? ( n4906 ) : ( iram_51 ) ;
assign n10941 = wr_addr[7:7] ;
assign n10942 =  ( n10941 ) == ( bv_1_0_n53 )  ;
assign n10943 =  ( wr_addr ) == ( bv_8_51_n171 )  ;
assign n10944 =  ( n10942 ) & (n10943 )  ;
assign n10945 =  ( n10944 ) & (wr )  ;
assign n10946 =  ( n10945 ) ? ( n5485 ) : ( iram_51 ) ;
assign n10947 = wr_addr[7:7] ;
assign n10948 =  ( n10947 ) == ( bv_1_0_n53 )  ;
assign n10949 =  ( wr_addr ) == ( bv_8_51_n171 )  ;
assign n10950 =  ( n10948 ) & (n10949 )  ;
assign n10951 =  ( n10950 ) & (wr )  ;
assign n10952 =  ( n10951 ) ? ( n5512 ) : ( iram_51 ) ;
assign n10953 = wr_addr[7:7] ;
assign n10954 =  ( n10953 ) == ( bv_1_0_n53 )  ;
assign n10955 =  ( wr_addr ) == ( bv_8_51_n171 )  ;
assign n10956 =  ( n10954 ) & (n10955 )  ;
assign n10957 =  ( n10956 ) & (wr )  ;
assign n10958 =  ( n10957 ) ? ( bv_8_0_n69 ) : ( iram_51 ) ;
assign n10959 = wr_addr[7:7] ;
assign n10960 =  ( n10959 ) == ( bv_1_0_n53 )  ;
assign n10961 =  ( wr_addr ) == ( bv_8_51_n171 )  ;
assign n10962 =  ( n10960 ) & (n10961 )  ;
assign n10963 =  ( n10962 ) & (wr )  ;
assign n10964 =  ( n10963 ) ? ( n5071 ) : ( iram_51 ) ;
assign n10965 = wr_addr[7:7] ;
assign n10966 =  ( n10965 ) == ( bv_1_0_n53 )  ;
assign n10967 =  ( wr_addr ) == ( bv_8_51_n171 )  ;
assign n10968 =  ( n10966 ) & (n10967 )  ;
assign n10969 =  ( n10968 ) & (wr )  ;
assign n10970 =  ( n10969 ) ? ( n5096 ) : ( iram_51 ) ;
assign n10971 = wr_addr[7:7] ;
assign n10972 =  ( n10971 ) == ( bv_1_0_n53 )  ;
assign n10973 =  ( wr_addr ) == ( bv_8_51_n171 )  ;
assign n10974 =  ( n10972 ) & (n10973 )  ;
assign n10975 =  ( n10974 ) & (wr )  ;
assign n10976 =  ( n10975 ) ? ( n5123 ) : ( iram_51 ) ;
assign n10977 = wr_addr[7:7] ;
assign n10978 =  ( n10977 ) == ( bv_1_0_n53 )  ;
assign n10979 =  ( wr_addr ) == ( bv_8_51_n171 )  ;
assign n10980 =  ( n10978 ) & (n10979 )  ;
assign n10981 =  ( n10980 ) & (wr )  ;
assign n10982 =  ( n10981 ) ? ( n5165 ) : ( iram_51 ) ;
assign n10983 = wr_addr[7:7] ;
assign n10984 =  ( n10983 ) == ( bv_1_0_n53 )  ;
assign n10985 =  ( wr_addr ) == ( bv_8_51_n171 )  ;
assign n10986 =  ( n10984 ) & (n10985 )  ;
assign n10987 =  ( n10986 ) & (wr )  ;
assign n10988 =  ( n10987 ) ? ( n5204 ) : ( iram_51 ) ;
assign n10989 = wr_addr[7:7] ;
assign n10990 =  ( n10989 ) == ( bv_1_0_n53 )  ;
assign n10991 =  ( wr_addr ) == ( bv_8_51_n171 )  ;
assign n10992 =  ( n10990 ) & (n10991 )  ;
assign n10993 =  ( n10992 ) & (wr )  ;
assign n10994 =  ( n10993 ) ? ( n5262 ) : ( iram_51 ) ;
assign n10995 = wr_addr[7:7] ;
assign n10996 =  ( n10995 ) == ( bv_1_0_n53 )  ;
assign n10997 =  ( wr_addr ) == ( bv_8_51_n171 )  ;
assign n10998 =  ( n10996 ) & (n10997 )  ;
assign n10999 =  ( n10998 ) & (wr )  ;
assign n11000 =  ( n10999 ) ? ( n5298 ) : ( iram_51 ) ;
assign n11001 = wr_addr[7:7] ;
assign n11002 =  ( n11001 ) == ( bv_1_0_n53 )  ;
assign n11003 =  ( wr_addr ) == ( bv_8_51_n171 )  ;
assign n11004 =  ( n11002 ) & (n11003 )  ;
assign n11005 =  ( n11004 ) & (wr )  ;
assign n11006 =  ( n11005 ) ? ( n5325 ) : ( iram_51 ) ;
assign n11007 = wr_addr[7:7] ;
assign n11008 =  ( n11007 ) == ( bv_1_0_n53 )  ;
assign n11009 =  ( wr_addr ) == ( bv_8_52_n173 )  ;
assign n11010 =  ( n11008 ) & (n11009 )  ;
assign n11011 =  ( n11010 ) & (wr )  ;
assign n11012 =  ( n11011 ) ? ( n4782 ) : ( iram_52 ) ;
assign n11013 = wr_addr[7:7] ;
assign n11014 =  ( n11013 ) == ( bv_1_0_n53 )  ;
assign n11015 =  ( wr_addr ) == ( bv_8_52_n173 )  ;
assign n11016 =  ( n11014 ) & (n11015 )  ;
assign n11017 =  ( n11016 ) & (wr )  ;
assign n11018 =  ( n11017 ) ? ( n4841 ) : ( iram_52 ) ;
assign n11019 = wr_addr[7:7] ;
assign n11020 =  ( n11019 ) == ( bv_1_0_n53 )  ;
assign n11021 =  ( wr_addr ) == ( bv_8_52_n173 )  ;
assign n11022 =  ( n11020 ) & (n11021 )  ;
assign n11023 =  ( n11022 ) & (wr )  ;
assign n11024 =  ( n11023 ) ? ( n5449 ) : ( iram_52 ) ;
assign n11025 = wr_addr[7:7] ;
assign n11026 =  ( n11025 ) == ( bv_1_0_n53 )  ;
assign n11027 =  ( wr_addr ) == ( bv_8_52_n173 )  ;
assign n11028 =  ( n11026 ) & (n11027 )  ;
assign n11029 =  ( n11028 ) & (wr )  ;
assign n11030 =  ( n11029 ) ? ( n4906 ) : ( iram_52 ) ;
assign n11031 = wr_addr[7:7] ;
assign n11032 =  ( n11031 ) == ( bv_1_0_n53 )  ;
assign n11033 =  ( wr_addr ) == ( bv_8_52_n173 )  ;
assign n11034 =  ( n11032 ) & (n11033 )  ;
assign n11035 =  ( n11034 ) & (wr )  ;
assign n11036 =  ( n11035 ) ? ( n5485 ) : ( iram_52 ) ;
assign n11037 = wr_addr[7:7] ;
assign n11038 =  ( n11037 ) == ( bv_1_0_n53 )  ;
assign n11039 =  ( wr_addr ) == ( bv_8_52_n173 )  ;
assign n11040 =  ( n11038 ) & (n11039 )  ;
assign n11041 =  ( n11040 ) & (wr )  ;
assign n11042 =  ( n11041 ) ? ( n5512 ) : ( iram_52 ) ;
assign n11043 = wr_addr[7:7] ;
assign n11044 =  ( n11043 ) == ( bv_1_0_n53 )  ;
assign n11045 =  ( wr_addr ) == ( bv_8_52_n173 )  ;
assign n11046 =  ( n11044 ) & (n11045 )  ;
assign n11047 =  ( n11046 ) & (wr )  ;
assign n11048 =  ( n11047 ) ? ( bv_8_0_n69 ) : ( iram_52 ) ;
assign n11049 = wr_addr[7:7] ;
assign n11050 =  ( n11049 ) == ( bv_1_0_n53 )  ;
assign n11051 =  ( wr_addr ) == ( bv_8_52_n173 )  ;
assign n11052 =  ( n11050 ) & (n11051 )  ;
assign n11053 =  ( n11052 ) & (wr )  ;
assign n11054 =  ( n11053 ) ? ( n5071 ) : ( iram_52 ) ;
assign n11055 = wr_addr[7:7] ;
assign n11056 =  ( n11055 ) == ( bv_1_0_n53 )  ;
assign n11057 =  ( wr_addr ) == ( bv_8_52_n173 )  ;
assign n11058 =  ( n11056 ) & (n11057 )  ;
assign n11059 =  ( n11058 ) & (wr )  ;
assign n11060 =  ( n11059 ) ? ( n5096 ) : ( iram_52 ) ;
assign n11061 = wr_addr[7:7] ;
assign n11062 =  ( n11061 ) == ( bv_1_0_n53 )  ;
assign n11063 =  ( wr_addr ) == ( bv_8_52_n173 )  ;
assign n11064 =  ( n11062 ) & (n11063 )  ;
assign n11065 =  ( n11064 ) & (wr )  ;
assign n11066 =  ( n11065 ) ? ( n5123 ) : ( iram_52 ) ;
assign n11067 = wr_addr[7:7] ;
assign n11068 =  ( n11067 ) == ( bv_1_0_n53 )  ;
assign n11069 =  ( wr_addr ) == ( bv_8_52_n173 )  ;
assign n11070 =  ( n11068 ) & (n11069 )  ;
assign n11071 =  ( n11070 ) & (wr )  ;
assign n11072 =  ( n11071 ) ? ( n5165 ) : ( iram_52 ) ;
assign n11073 = wr_addr[7:7] ;
assign n11074 =  ( n11073 ) == ( bv_1_0_n53 )  ;
assign n11075 =  ( wr_addr ) == ( bv_8_52_n173 )  ;
assign n11076 =  ( n11074 ) & (n11075 )  ;
assign n11077 =  ( n11076 ) & (wr )  ;
assign n11078 =  ( n11077 ) ? ( n5204 ) : ( iram_52 ) ;
assign n11079 = wr_addr[7:7] ;
assign n11080 =  ( n11079 ) == ( bv_1_0_n53 )  ;
assign n11081 =  ( wr_addr ) == ( bv_8_52_n173 )  ;
assign n11082 =  ( n11080 ) & (n11081 )  ;
assign n11083 =  ( n11082 ) & (wr )  ;
assign n11084 =  ( n11083 ) ? ( n5262 ) : ( iram_52 ) ;
assign n11085 = wr_addr[7:7] ;
assign n11086 =  ( n11085 ) == ( bv_1_0_n53 )  ;
assign n11087 =  ( wr_addr ) == ( bv_8_52_n173 )  ;
assign n11088 =  ( n11086 ) & (n11087 )  ;
assign n11089 =  ( n11088 ) & (wr )  ;
assign n11090 =  ( n11089 ) ? ( n5298 ) : ( iram_52 ) ;
assign n11091 = wr_addr[7:7] ;
assign n11092 =  ( n11091 ) == ( bv_1_0_n53 )  ;
assign n11093 =  ( wr_addr ) == ( bv_8_52_n173 )  ;
assign n11094 =  ( n11092 ) & (n11093 )  ;
assign n11095 =  ( n11094 ) & (wr )  ;
assign n11096 =  ( n11095 ) ? ( n5325 ) : ( iram_52 ) ;
assign n11097 = wr_addr[7:7] ;
assign n11098 =  ( n11097 ) == ( bv_1_0_n53 )  ;
assign n11099 =  ( wr_addr ) == ( bv_8_53_n175 )  ;
assign n11100 =  ( n11098 ) & (n11099 )  ;
assign n11101 =  ( n11100 ) & (wr )  ;
assign n11102 =  ( n11101 ) ? ( n4782 ) : ( iram_53 ) ;
assign n11103 = wr_addr[7:7] ;
assign n11104 =  ( n11103 ) == ( bv_1_0_n53 )  ;
assign n11105 =  ( wr_addr ) == ( bv_8_53_n175 )  ;
assign n11106 =  ( n11104 ) & (n11105 )  ;
assign n11107 =  ( n11106 ) & (wr )  ;
assign n11108 =  ( n11107 ) ? ( n4841 ) : ( iram_53 ) ;
assign n11109 = wr_addr[7:7] ;
assign n11110 =  ( n11109 ) == ( bv_1_0_n53 )  ;
assign n11111 =  ( wr_addr ) == ( bv_8_53_n175 )  ;
assign n11112 =  ( n11110 ) & (n11111 )  ;
assign n11113 =  ( n11112 ) & (wr )  ;
assign n11114 =  ( n11113 ) ? ( n5449 ) : ( iram_53 ) ;
assign n11115 = wr_addr[7:7] ;
assign n11116 =  ( n11115 ) == ( bv_1_0_n53 )  ;
assign n11117 =  ( wr_addr ) == ( bv_8_53_n175 )  ;
assign n11118 =  ( n11116 ) & (n11117 )  ;
assign n11119 =  ( n11118 ) & (wr )  ;
assign n11120 =  ( n11119 ) ? ( n4906 ) : ( iram_53 ) ;
assign n11121 = wr_addr[7:7] ;
assign n11122 =  ( n11121 ) == ( bv_1_0_n53 )  ;
assign n11123 =  ( wr_addr ) == ( bv_8_53_n175 )  ;
assign n11124 =  ( n11122 ) & (n11123 )  ;
assign n11125 =  ( n11124 ) & (wr )  ;
assign n11126 =  ( n11125 ) ? ( n5485 ) : ( iram_53 ) ;
assign n11127 = wr_addr[7:7] ;
assign n11128 =  ( n11127 ) == ( bv_1_0_n53 )  ;
assign n11129 =  ( wr_addr ) == ( bv_8_53_n175 )  ;
assign n11130 =  ( n11128 ) & (n11129 )  ;
assign n11131 =  ( n11130 ) & (wr )  ;
assign n11132 =  ( n11131 ) ? ( n5512 ) : ( iram_53 ) ;
assign n11133 = wr_addr[7:7] ;
assign n11134 =  ( n11133 ) == ( bv_1_0_n53 )  ;
assign n11135 =  ( wr_addr ) == ( bv_8_53_n175 )  ;
assign n11136 =  ( n11134 ) & (n11135 )  ;
assign n11137 =  ( n11136 ) & (wr )  ;
assign n11138 =  ( n11137 ) ? ( bv_8_0_n69 ) : ( iram_53 ) ;
assign n11139 = wr_addr[7:7] ;
assign n11140 =  ( n11139 ) == ( bv_1_0_n53 )  ;
assign n11141 =  ( wr_addr ) == ( bv_8_53_n175 )  ;
assign n11142 =  ( n11140 ) & (n11141 )  ;
assign n11143 =  ( n11142 ) & (wr )  ;
assign n11144 =  ( n11143 ) ? ( n5071 ) : ( iram_53 ) ;
assign n11145 = wr_addr[7:7] ;
assign n11146 =  ( n11145 ) == ( bv_1_0_n53 )  ;
assign n11147 =  ( wr_addr ) == ( bv_8_53_n175 )  ;
assign n11148 =  ( n11146 ) & (n11147 )  ;
assign n11149 =  ( n11148 ) & (wr )  ;
assign n11150 =  ( n11149 ) ? ( n5096 ) : ( iram_53 ) ;
assign n11151 = wr_addr[7:7] ;
assign n11152 =  ( n11151 ) == ( bv_1_0_n53 )  ;
assign n11153 =  ( wr_addr ) == ( bv_8_53_n175 )  ;
assign n11154 =  ( n11152 ) & (n11153 )  ;
assign n11155 =  ( n11154 ) & (wr )  ;
assign n11156 =  ( n11155 ) ? ( n5123 ) : ( iram_53 ) ;
assign n11157 = wr_addr[7:7] ;
assign n11158 =  ( n11157 ) == ( bv_1_0_n53 )  ;
assign n11159 =  ( wr_addr ) == ( bv_8_53_n175 )  ;
assign n11160 =  ( n11158 ) & (n11159 )  ;
assign n11161 =  ( n11160 ) & (wr )  ;
assign n11162 =  ( n11161 ) ? ( n5165 ) : ( iram_53 ) ;
assign n11163 = wr_addr[7:7] ;
assign n11164 =  ( n11163 ) == ( bv_1_0_n53 )  ;
assign n11165 =  ( wr_addr ) == ( bv_8_53_n175 )  ;
assign n11166 =  ( n11164 ) & (n11165 )  ;
assign n11167 =  ( n11166 ) & (wr )  ;
assign n11168 =  ( n11167 ) ? ( n5204 ) : ( iram_53 ) ;
assign n11169 = wr_addr[7:7] ;
assign n11170 =  ( n11169 ) == ( bv_1_0_n53 )  ;
assign n11171 =  ( wr_addr ) == ( bv_8_53_n175 )  ;
assign n11172 =  ( n11170 ) & (n11171 )  ;
assign n11173 =  ( n11172 ) & (wr )  ;
assign n11174 =  ( n11173 ) ? ( n5262 ) : ( iram_53 ) ;
assign n11175 = wr_addr[7:7] ;
assign n11176 =  ( n11175 ) == ( bv_1_0_n53 )  ;
assign n11177 =  ( wr_addr ) == ( bv_8_53_n175 )  ;
assign n11178 =  ( n11176 ) & (n11177 )  ;
assign n11179 =  ( n11178 ) & (wr )  ;
assign n11180 =  ( n11179 ) ? ( n5298 ) : ( iram_53 ) ;
assign n11181 = wr_addr[7:7] ;
assign n11182 =  ( n11181 ) == ( bv_1_0_n53 )  ;
assign n11183 =  ( wr_addr ) == ( bv_8_53_n175 )  ;
assign n11184 =  ( n11182 ) & (n11183 )  ;
assign n11185 =  ( n11184 ) & (wr )  ;
assign n11186 =  ( n11185 ) ? ( n5325 ) : ( iram_53 ) ;
assign n11187 = wr_addr[7:7] ;
assign n11188 =  ( n11187 ) == ( bv_1_0_n53 )  ;
assign n11189 =  ( wr_addr ) == ( bv_8_54_n177 )  ;
assign n11190 =  ( n11188 ) & (n11189 )  ;
assign n11191 =  ( n11190 ) & (wr )  ;
assign n11192 =  ( n11191 ) ? ( n4782 ) : ( iram_54 ) ;
assign n11193 = wr_addr[7:7] ;
assign n11194 =  ( n11193 ) == ( bv_1_0_n53 )  ;
assign n11195 =  ( wr_addr ) == ( bv_8_54_n177 )  ;
assign n11196 =  ( n11194 ) & (n11195 )  ;
assign n11197 =  ( n11196 ) & (wr )  ;
assign n11198 =  ( n11197 ) ? ( n4841 ) : ( iram_54 ) ;
assign n11199 = wr_addr[7:7] ;
assign n11200 =  ( n11199 ) == ( bv_1_0_n53 )  ;
assign n11201 =  ( wr_addr ) == ( bv_8_54_n177 )  ;
assign n11202 =  ( n11200 ) & (n11201 )  ;
assign n11203 =  ( n11202 ) & (wr )  ;
assign n11204 =  ( n11203 ) ? ( n5449 ) : ( iram_54 ) ;
assign n11205 = wr_addr[7:7] ;
assign n11206 =  ( n11205 ) == ( bv_1_0_n53 )  ;
assign n11207 =  ( wr_addr ) == ( bv_8_54_n177 )  ;
assign n11208 =  ( n11206 ) & (n11207 )  ;
assign n11209 =  ( n11208 ) & (wr )  ;
assign n11210 =  ( n11209 ) ? ( n4906 ) : ( iram_54 ) ;
assign n11211 = wr_addr[7:7] ;
assign n11212 =  ( n11211 ) == ( bv_1_0_n53 )  ;
assign n11213 =  ( wr_addr ) == ( bv_8_54_n177 )  ;
assign n11214 =  ( n11212 ) & (n11213 )  ;
assign n11215 =  ( n11214 ) & (wr )  ;
assign n11216 =  ( n11215 ) ? ( n5485 ) : ( iram_54 ) ;
assign n11217 = wr_addr[7:7] ;
assign n11218 =  ( n11217 ) == ( bv_1_0_n53 )  ;
assign n11219 =  ( wr_addr ) == ( bv_8_54_n177 )  ;
assign n11220 =  ( n11218 ) & (n11219 )  ;
assign n11221 =  ( n11220 ) & (wr )  ;
assign n11222 =  ( n11221 ) ? ( n5512 ) : ( iram_54 ) ;
assign n11223 = wr_addr[7:7] ;
assign n11224 =  ( n11223 ) == ( bv_1_0_n53 )  ;
assign n11225 =  ( wr_addr ) == ( bv_8_54_n177 )  ;
assign n11226 =  ( n11224 ) & (n11225 )  ;
assign n11227 =  ( n11226 ) & (wr )  ;
assign n11228 =  ( n11227 ) ? ( bv_8_0_n69 ) : ( iram_54 ) ;
assign n11229 = wr_addr[7:7] ;
assign n11230 =  ( n11229 ) == ( bv_1_0_n53 )  ;
assign n11231 =  ( wr_addr ) == ( bv_8_54_n177 )  ;
assign n11232 =  ( n11230 ) & (n11231 )  ;
assign n11233 =  ( n11232 ) & (wr )  ;
assign n11234 =  ( n11233 ) ? ( n5071 ) : ( iram_54 ) ;
assign n11235 = wr_addr[7:7] ;
assign n11236 =  ( n11235 ) == ( bv_1_0_n53 )  ;
assign n11237 =  ( wr_addr ) == ( bv_8_54_n177 )  ;
assign n11238 =  ( n11236 ) & (n11237 )  ;
assign n11239 =  ( n11238 ) & (wr )  ;
assign n11240 =  ( n11239 ) ? ( n5096 ) : ( iram_54 ) ;
assign n11241 = wr_addr[7:7] ;
assign n11242 =  ( n11241 ) == ( bv_1_0_n53 )  ;
assign n11243 =  ( wr_addr ) == ( bv_8_54_n177 )  ;
assign n11244 =  ( n11242 ) & (n11243 )  ;
assign n11245 =  ( n11244 ) & (wr )  ;
assign n11246 =  ( n11245 ) ? ( n5123 ) : ( iram_54 ) ;
assign n11247 = wr_addr[7:7] ;
assign n11248 =  ( n11247 ) == ( bv_1_0_n53 )  ;
assign n11249 =  ( wr_addr ) == ( bv_8_54_n177 )  ;
assign n11250 =  ( n11248 ) & (n11249 )  ;
assign n11251 =  ( n11250 ) & (wr )  ;
assign n11252 =  ( n11251 ) ? ( n5165 ) : ( iram_54 ) ;
assign n11253 = wr_addr[7:7] ;
assign n11254 =  ( n11253 ) == ( bv_1_0_n53 )  ;
assign n11255 =  ( wr_addr ) == ( bv_8_54_n177 )  ;
assign n11256 =  ( n11254 ) & (n11255 )  ;
assign n11257 =  ( n11256 ) & (wr )  ;
assign n11258 =  ( n11257 ) ? ( n5204 ) : ( iram_54 ) ;
assign n11259 = wr_addr[7:7] ;
assign n11260 =  ( n11259 ) == ( bv_1_0_n53 )  ;
assign n11261 =  ( wr_addr ) == ( bv_8_54_n177 )  ;
assign n11262 =  ( n11260 ) & (n11261 )  ;
assign n11263 =  ( n11262 ) & (wr )  ;
assign n11264 =  ( n11263 ) ? ( n5262 ) : ( iram_54 ) ;
assign n11265 = wr_addr[7:7] ;
assign n11266 =  ( n11265 ) == ( bv_1_0_n53 )  ;
assign n11267 =  ( wr_addr ) == ( bv_8_54_n177 )  ;
assign n11268 =  ( n11266 ) & (n11267 )  ;
assign n11269 =  ( n11268 ) & (wr )  ;
assign n11270 =  ( n11269 ) ? ( n5298 ) : ( iram_54 ) ;
assign n11271 = wr_addr[7:7] ;
assign n11272 =  ( n11271 ) == ( bv_1_0_n53 )  ;
assign n11273 =  ( wr_addr ) == ( bv_8_54_n177 )  ;
assign n11274 =  ( n11272 ) & (n11273 )  ;
assign n11275 =  ( n11274 ) & (wr )  ;
assign n11276 =  ( n11275 ) ? ( n5325 ) : ( iram_54 ) ;
assign n11277 = wr_addr[7:7] ;
assign n11278 =  ( n11277 ) == ( bv_1_0_n53 )  ;
assign n11279 =  ( wr_addr ) == ( bv_8_55_n179 )  ;
assign n11280 =  ( n11278 ) & (n11279 )  ;
assign n11281 =  ( n11280 ) & (wr )  ;
assign n11282 =  ( n11281 ) ? ( n4782 ) : ( iram_55 ) ;
assign n11283 = wr_addr[7:7] ;
assign n11284 =  ( n11283 ) == ( bv_1_0_n53 )  ;
assign n11285 =  ( wr_addr ) == ( bv_8_55_n179 )  ;
assign n11286 =  ( n11284 ) & (n11285 )  ;
assign n11287 =  ( n11286 ) & (wr )  ;
assign n11288 =  ( n11287 ) ? ( n4841 ) : ( iram_55 ) ;
assign n11289 = wr_addr[7:7] ;
assign n11290 =  ( n11289 ) == ( bv_1_0_n53 )  ;
assign n11291 =  ( wr_addr ) == ( bv_8_55_n179 )  ;
assign n11292 =  ( n11290 ) & (n11291 )  ;
assign n11293 =  ( n11292 ) & (wr )  ;
assign n11294 =  ( n11293 ) ? ( n5449 ) : ( iram_55 ) ;
assign n11295 = wr_addr[7:7] ;
assign n11296 =  ( n11295 ) == ( bv_1_0_n53 )  ;
assign n11297 =  ( wr_addr ) == ( bv_8_55_n179 )  ;
assign n11298 =  ( n11296 ) & (n11297 )  ;
assign n11299 =  ( n11298 ) & (wr )  ;
assign n11300 =  ( n11299 ) ? ( n4906 ) : ( iram_55 ) ;
assign n11301 = wr_addr[7:7] ;
assign n11302 =  ( n11301 ) == ( bv_1_0_n53 )  ;
assign n11303 =  ( wr_addr ) == ( bv_8_55_n179 )  ;
assign n11304 =  ( n11302 ) & (n11303 )  ;
assign n11305 =  ( n11304 ) & (wr )  ;
assign n11306 =  ( n11305 ) ? ( n5485 ) : ( iram_55 ) ;
assign n11307 = wr_addr[7:7] ;
assign n11308 =  ( n11307 ) == ( bv_1_0_n53 )  ;
assign n11309 =  ( wr_addr ) == ( bv_8_55_n179 )  ;
assign n11310 =  ( n11308 ) & (n11309 )  ;
assign n11311 =  ( n11310 ) & (wr )  ;
assign n11312 =  ( n11311 ) ? ( n5512 ) : ( iram_55 ) ;
assign n11313 = wr_addr[7:7] ;
assign n11314 =  ( n11313 ) == ( bv_1_0_n53 )  ;
assign n11315 =  ( wr_addr ) == ( bv_8_55_n179 )  ;
assign n11316 =  ( n11314 ) & (n11315 )  ;
assign n11317 =  ( n11316 ) & (wr )  ;
assign n11318 =  ( n11317 ) ? ( bv_8_0_n69 ) : ( iram_55 ) ;
assign n11319 = wr_addr[7:7] ;
assign n11320 =  ( n11319 ) == ( bv_1_0_n53 )  ;
assign n11321 =  ( wr_addr ) == ( bv_8_55_n179 )  ;
assign n11322 =  ( n11320 ) & (n11321 )  ;
assign n11323 =  ( n11322 ) & (wr )  ;
assign n11324 =  ( n11323 ) ? ( n5071 ) : ( iram_55 ) ;
assign n11325 = wr_addr[7:7] ;
assign n11326 =  ( n11325 ) == ( bv_1_0_n53 )  ;
assign n11327 =  ( wr_addr ) == ( bv_8_55_n179 )  ;
assign n11328 =  ( n11326 ) & (n11327 )  ;
assign n11329 =  ( n11328 ) & (wr )  ;
assign n11330 =  ( n11329 ) ? ( n5096 ) : ( iram_55 ) ;
assign n11331 = wr_addr[7:7] ;
assign n11332 =  ( n11331 ) == ( bv_1_0_n53 )  ;
assign n11333 =  ( wr_addr ) == ( bv_8_55_n179 )  ;
assign n11334 =  ( n11332 ) & (n11333 )  ;
assign n11335 =  ( n11334 ) & (wr )  ;
assign n11336 =  ( n11335 ) ? ( n5123 ) : ( iram_55 ) ;
assign n11337 = wr_addr[7:7] ;
assign n11338 =  ( n11337 ) == ( bv_1_0_n53 )  ;
assign n11339 =  ( wr_addr ) == ( bv_8_55_n179 )  ;
assign n11340 =  ( n11338 ) & (n11339 )  ;
assign n11341 =  ( n11340 ) & (wr )  ;
assign n11342 =  ( n11341 ) ? ( n5165 ) : ( iram_55 ) ;
assign n11343 = wr_addr[7:7] ;
assign n11344 =  ( n11343 ) == ( bv_1_0_n53 )  ;
assign n11345 =  ( wr_addr ) == ( bv_8_55_n179 )  ;
assign n11346 =  ( n11344 ) & (n11345 )  ;
assign n11347 =  ( n11346 ) & (wr )  ;
assign n11348 =  ( n11347 ) ? ( n5204 ) : ( iram_55 ) ;
assign n11349 = wr_addr[7:7] ;
assign n11350 =  ( n11349 ) == ( bv_1_0_n53 )  ;
assign n11351 =  ( wr_addr ) == ( bv_8_55_n179 )  ;
assign n11352 =  ( n11350 ) & (n11351 )  ;
assign n11353 =  ( n11352 ) & (wr )  ;
assign n11354 =  ( n11353 ) ? ( n5262 ) : ( iram_55 ) ;
assign n11355 = wr_addr[7:7] ;
assign n11356 =  ( n11355 ) == ( bv_1_0_n53 )  ;
assign n11357 =  ( wr_addr ) == ( bv_8_55_n179 )  ;
assign n11358 =  ( n11356 ) & (n11357 )  ;
assign n11359 =  ( n11358 ) & (wr )  ;
assign n11360 =  ( n11359 ) ? ( n5298 ) : ( iram_55 ) ;
assign n11361 = wr_addr[7:7] ;
assign n11362 =  ( n11361 ) == ( bv_1_0_n53 )  ;
assign n11363 =  ( wr_addr ) == ( bv_8_55_n179 )  ;
assign n11364 =  ( n11362 ) & (n11363 )  ;
assign n11365 =  ( n11364 ) & (wr )  ;
assign n11366 =  ( n11365 ) ? ( n5325 ) : ( iram_55 ) ;
assign n11367 = wr_addr[7:7] ;
assign n11368 =  ( n11367 ) == ( bv_1_0_n53 )  ;
assign n11369 =  ( wr_addr ) == ( bv_8_56_n181 )  ;
assign n11370 =  ( n11368 ) & (n11369 )  ;
assign n11371 =  ( n11370 ) & (wr )  ;
assign n11372 =  ( n11371 ) ? ( n4782 ) : ( iram_56 ) ;
assign n11373 = wr_addr[7:7] ;
assign n11374 =  ( n11373 ) == ( bv_1_0_n53 )  ;
assign n11375 =  ( wr_addr ) == ( bv_8_56_n181 )  ;
assign n11376 =  ( n11374 ) & (n11375 )  ;
assign n11377 =  ( n11376 ) & (wr )  ;
assign n11378 =  ( n11377 ) ? ( n4841 ) : ( iram_56 ) ;
assign n11379 = wr_addr[7:7] ;
assign n11380 =  ( n11379 ) == ( bv_1_0_n53 )  ;
assign n11381 =  ( wr_addr ) == ( bv_8_56_n181 )  ;
assign n11382 =  ( n11380 ) & (n11381 )  ;
assign n11383 =  ( n11382 ) & (wr )  ;
assign n11384 =  ( n11383 ) ? ( n5449 ) : ( iram_56 ) ;
assign n11385 = wr_addr[7:7] ;
assign n11386 =  ( n11385 ) == ( bv_1_0_n53 )  ;
assign n11387 =  ( wr_addr ) == ( bv_8_56_n181 )  ;
assign n11388 =  ( n11386 ) & (n11387 )  ;
assign n11389 =  ( n11388 ) & (wr )  ;
assign n11390 =  ( n11389 ) ? ( n4906 ) : ( iram_56 ) ;
assign n11391 = wr_addr[7:7] ;
assign n11392 =  ( n11391 ) == ( bv_1_0_n53 )  ;
assign n11393 =  ( wr_addr ) == ( bv_8_56_n181 )  ;
assign n11394 =  ( n11392 ) & (n11393 )  ;
assign n11395 =  ( n11394 ) & (wr )  ;
assign n11396 =  ( n11395 ) ? ( n5485 ) : ( iram_56 ) ;
assign n11397 = wr_addr[7:7] ;
assign n11398 =  ( n11397 ) == ( bv_1_0_n53 )  ;
assign n11399 =  ( wr_addr ) == ( bv_8_56_n181 )  ;
assign n11400 =  ( n11398 ) & (n11399 )  ;
assign n11401 =  ( n11400 ) & (wr )  ;
assign n11402 =  ( n11401 ) ? ( n5512 ) : ( iram_56 ) ;
assign n11403 = wr_addr[7:7] ;
assign n11404 =  ( n11403 ) == ( bv_1_0_n53 )  ;
assign n11405 =  ( wr_addr ) == ( bv_8_56_n181 )  ;
assign n11406 =  ( n11404 ) & (n11405 )  ;
assign n11407 =  ( n11406 ) & (wr )  ;
assign n11408 =  ( n11407 ) ? ( bv_8_0_n69 ) : ( iram_56 ) ;
assign n11409 = wr_addr[7:7] ;
assign n11410 =  ( n11409 ) == ( bv_1_0_n53 )  ;
assign n11411 =  ( wr_addr ) == ( bv_8_56_n181 )  ;
assign n11412 =  ( n11410 ) & (n11411 )  ;
assign n11413 =  ( n11412 ) & (wr )  ;
assign n11414 =  ( n11413 ) ? ( n5071 ) : ( iram_56 ) ;
assign n11415 = wr_addr[7:7] ;
assign n11416 =  ( n11415 ) == ( bv_1_0_n53 )  ;
assign n11417 =  ( wr_addr ) == ( bv_8_56_n181 )  ;
assign n11418 =  ( n11416 ) & (n11417 )  ;
assign n11419 =  ( n11418 ) & (wr )  ;
assign n11420 =  ( n11419 ) ? ( n5096 ) : ( iram_56 ) ;
assign n11421 = wr_addr[7:7] ;
assign n11422 =  ( n11421 ) == ( bv_1_0_n53 )  ;
assign n11423 =  ( wr_addr ) == ( bv_8_56_n181 )  ;
assign n11424 =  ( n11422 ) & (n11423 )  ;
assign n11425 =  ( n11424 ) & (wr )  ;
assign n11426 =  ( n11425 ) ? ( n5123 ) : ( iram_56 ) ;
assign n11427 = wr_addr[7:7] ;
assign n11428 =  ( n11427 ) == ( bv_1_0_n53 )  ;
assign n11429 =  ( wr_addr ) == ( bv_8_56_n181 )  ;
assign n11430 =  ( n11428 ) & (n11429 )  ;
assign n11431 =  ( n11430 ) & (wr )  ;
assign n11432 =  ( n11431 ) ? ( n5165 ) : ( iram_56 ) ;
assign n11433 = wr_addr[7:7] ;
assign n11434 =  ( n11433 ) == ( bv_1_0_n53 )  ;
assign n11435 =  ( wr_addr ) == ( bv_8_56_n181 )  ;
assign n11436 =  ( n11434 ) & (n11435 )  ;
assign n11437 =  ( n11436 ) & (wr )  ;
assign n11438 =  ( n11437 ) ? ( n5204 ) : ( iram_56 ) ;
assign n11439 = wr_addr[7:7] ;
assign n11440 =  ( n11439 ) == ( bv_1_0_n53 )  ;
assign n11441 =  ( wr_addr ) == ( bv_8_56_n181 )  ;
assign n11442 =  ( n11440 ) & (n11441 )  ;
assign n11443 =  ( n11442 ) & (wr )  ;
assign n11444 =  ( n11443 ) ? ( n5262 ) : ( iram_56 ) ;
assign n11445 = wr_addr[7:7] ;
assign n11446 =  ( n11445 ) == ( bv_1_0_n53 )  ;
assign n11447 =  ( wr_addr ) == ( bv_8_56_n181 )  ;
assign n11448 =  ( n11446 ) & (n11447 )  ;
assign n11449 =  ( n11448 ) & (wr )  ;
assign n11450 =  ( n11449 ) ? ( n5298 ) : ( iram_56 ) ;
assign n11451 = wr_addr[7:7] ;
assign n11452 =  ( n11451 ) == ( bv_1_0_n53 )  ;
assign n11453 =  ( wr_addr ) == ( bv_8_56_n181 )  ;
assign n11454 =  ( n11452 ) & (n11453 )  ;
assign n11455 =  ( n11454 ) & (wr )  ;
assign n11456 =  ( n11455 ) ? ( n5325 ) : ( iram_56 ) ;
assign n11457 = wr_addr[7:7] ;
assign n11458 =  ( n11457 ) == ( bv_1_0_n53 )  ;
assign n11459 =  ( wr_addr ) == ( bv_8_57_n183 )  ;
assign n11460 =  ( n11458 ) & (n11459 )  ;
assign n11461 =  ( n11460 ) & (wr )  ;
assign n11462 =  ( n11461 ) ? ( n4782 ) : ( iram_57 ) ;
assign n11463 = wr_addr[7:7] ;
assign n11464 =  ( n11463 ) == ( bv_1_0_n53 )  ;
assign n11465 =  ( wr_addr ) == ( bv_8_57_n183 )  ;
assign n11466 =  ( n11464 ) & (n11465 )  ;
assign n11467 =  ( n11466 ) & (wr )  ;
assign n11468 =  ( n11467 ) ? ( n4841 ) : ( iram_57 ) ;
assign n11469 = wr_addr[7:7] ;
assign n11470 =  ( n11469 ) == ( bv_1_0_n53 )  ;
assign n11471 =  ( wr_addr ) == ( bv_8_57_n183 )  ;
assign n11472 =  ( n11470 ) & (n11471 )  ;
assign n11473 =  ( n11472 ) & (wr )  ;
assign n11474 =  ( n11473 ) ? ( n5449 ) : ( iram_57 ) ;
assign n11475 = wr_addr[7:7] ;
assign n11476 =  ( n11475 ) == ( bv_1_0_n53 )  ;
assign n11477 =  ( wr_addr ) == ( bv_8_57_n183 )  ;
assign n11478 =  ( n11476 ) & (n11477 )  ;
assign n11479 =  ( n11478 ) & (wr )  ;
assign n11480 =  ( n11479 ) ? ( n4906 ) : ( iram_57 ) ;
assign n11481 = wr_addr[7:7] ;
assign n11482 =  ( n11481 ) == ( bv_1_0_n53 )  ;
assign n11483 =  ( wr_addr ) == ( bv_8_57_n183 )  ;
assign n11484 =  ( n11482 ) & (n11483 )  ;
assign n11485 =  ( n11484 ) & (wr )  ;
assign n11486 =  ( n11485 ) ? ( n5485 ) : ( iram_57 ) ;
assign n11487 = wr_addr[7:7] ;
assign n11488 =  ( n11487 ) == ( bv_1_0_n53 )  ;
assign n11489 =  ( wr_addr ) == ( bv_8_57_n183 )  ;
assign n11490 =  ( n11488 ) & (n11489 )  ;
assign n11491 =  ( n11490 ) & (wr )  ;
assign n11492 =  ( n11491 ) ? ( n5512 ) : ( iram_57 ) ;
assign n11493 = wr_addr[7:7] ;
assign n11494 =  ( n11493 ) == ( bv_1_0_n53 )  ;
assign n11495 =  ( wr_addr ) == ( bv_8_57_n183 )  ;
assign n11496 =  ( n11494 ) & (n11495 )  ;
assign n11497 =  ( n11496 ) & (wr )  ;
assign n11498 =  ( n11497 ) ? ( bv_8_0_n69 ) : ( iram_57 ) ;
assign n11499 = wr_addr[7:7] ;
assign n11500 =  ( n11499 ) == ( bv_1_0_n53 )  ;
assign n11501 =  ( wr_addr ) == ( bv_8_57_n183 )  ;
assign n11502 =  ( n11500 ) & (n11501 )  ;
assign n11503 =  ( n11502 ) & (wr )  ;
assign n11504 =  ( n11503 ) ? ( n5071 ) : ( iram_57 ) ;
assign n11505 = wr_addr[7:7] ;
assign n11506 =  ( n11505 ) == ( bv_1_0_n53 )  ;
assign n11507 =  ( wr_addr ) == ( bv_8_57_n183 )  ;
assign n11508 =  ( n11506 ) & (n11507 )  ;
assign n11509 =  ( n11508 ) & (wr )  ;
assign n11510 =  ( n11509 ) ? ( n5096 ) : ( iram_57 ) ;
assign n11511 = wr_addr[7:7] ;
assign n11512 =  ( n11511 ) == ( bv_1_0_n53 )  ;
assign n11513 =  ( wr_addr ) == ( bv_8_57_n183 )  ;
assign n11514 =  ( n11512 ) & (n11513 )  ;
assign n11515 =  ( n11514 ) & (wr )  ;
assign n11516 =  ( n11515 ) ? ( n5123 ) : ( iram_57 ) ;
assign n11517 = wr_addr[7:7] ;
assign n11518 =  ( n11517 ) == ( bv_1_0_n53 )  ;
assign n11519 =  ( wr_addr ) == ( bv_8_57_n183 )  ;
assign n11520 =  ( n11518 ) & (n11519 )  ;
assign n11521 =  ( n11520 ) & (wr )  ;
assign n11522 =  ( n11521 ) ? ( n5165 ) : ( iram_57 ) ;
assign n11523 = wr_addr[7:7] ;
assign n11524 =  ( n11523 ) == ( bv_1_0_n53 )  ;
assign n11525 =  ( wr_addr ) == ( bv_8_57_n183 )  ;
assign n11526 =  ( n11524 ) & (n11525 )  ;
assign n11527 =  ( n11526 ) & (wr )  ;
assign n11528 =  ( n11527 ) ? ( n5204 ) : ( iram_57 ) ;
assign n11529 = wr_addr[7:7] ;
assign n11530 =  ( n11529 ) == ( bv_1_0_n53 )  ;
assign n11531 =  ( wr_addr ) == ( bv_8_57_n183 )  ;
assign n11532 =  ( n11530 ) & (n11531 )  ;
assign n11533 =  ( n11532 ) & (wr )  ;
assign n11534 =  ( n11533 ) ? ( n5262 ) : ( iram_57 ) ;
assign n11535 = wr_addr[7:7] ;
assign n11536 =  ( n11535 ) == ( bv_1_0_n53 )  ;
assign n11537 =  ( wr_addr ) == ( bv_8_57_n183 )  ;
assign n11538 =  ( n11536 ) & (n11537 )  ;
assign n11539 =  ( n11538 ) & (wr )  ;
assign n11540 =  ( n11539 ) ? ( n5298 ) : ( iram_57 ) ;
assign n11541 = wr_addr[7:7] ;
assign n11542 =  ( n11541 ) == ( bv_1_0_n53 )  ;
assign n11543 =  ( wr_addr ) == ( bv_8_57_n183 )  ;
assign n11544 =  ( n11542 ) & (n11543 )  ;
assign n11545 =  ( n11544 ) & (wr )  ;
assign n11546 =  ( n11545 ) ? ( n5325 ) : ( iram_57 ) ;
assign n11547 = wr_addr[7:7] ;
assign n11548 =  ( n11547 ) == ( bv_1_0_n53 )  ;
assign n11549 =  ( wr_addr ) == ( bv_8_58_n185 )  ;
assign n11550 =  ( n11548 ) & (n11549 )  ;
assign n11551 =  ( n11550 ) & (wr )  ;
assign n11552 =  ( n11551 ) ? ( n4782 ) : ( iram_58 ) ;
assign n11553 = wr_addr[7:7] ;
assign n11554 =  ( n11553 ) == ( bv_1_0_n53 )  ;
assign n11555 =  ( wr_addr ) == ( bv_8_58_n185 )  ;
assign n11556 =  ( n11554 ) & (n11555 )  ;
assign n11557 =  ( n11556 ) & (wr )  ;
assign n11558 =  ( n11557 ) ? ( n4841 ) : ( iram_58 ) ;
assign n11559 = wr_addr[7:7] ;
assign n11560 =  ( n11559 ) == ( bv_1_0_n53 )  ;
assign n11561 =  ( wr_addr ) == ( bv_8_58_n185 )  ;
assign n11562 =  ( n11560 ) & (n11561 )  ;
assign n11563 =  ( n11562 ) & (wr )  ;
assign n11564 =  ( n11563 ) ? ( n5449 ) : ( iram_58 ) ;
assign n11565 = wr_addr[7:7] ;
assign n11566 =  ( n11565 ) == ( bv_1_0_n53 )  ;
assign n11567 =  ( wr_addr ) == ( bv_8_58_n185 )  ;
assign n11568 =  ( n11566 ) & (n11567 )  ;
assign n11569 =  ( n11568 ) & (wr )  ;
assign n11570 =  ( n11569 ) ? ( n4906 ) : ( iram_58 ) ;
assign n11571 = wr_addr[7:7] ;
assign n11572 =  ( n11571 ) == ( bv_1_0_n53 )  ;
assign n11573 =  ( wr_addr ) == ( bv_8_58_n185 )  ;
assign n11574 =  ( n11572 ) & (n11573 )  ;
assign n11575 =  ( n11574 ) & (wr )  ;
assign n11576 =  ( n11575 ) ? ( n5485 ) : ( iram_58 ) ;
assign n11577 = wr_addr[7:7] ;
assign n11578 =  ( n11577 ) == ( bv_1_0_n53 )  ;
assign n11579 =  ( wr_addr ) == ( bv_8_58_n185 )  ;
assign n11580 =  ( n11578 ) & (n11579 )  ;
assign n11581 =  ( n11580 ) & (wr )  ;
assign n11582 =  ( n11581 ) ? ( n5512 ) : ( iram_58 ) ;
assign n11583 = wr_addr[7:7] ;
assign n11584 =  ( n11583 ) == ( bv_1_0_n53 )  ;
assign n11585 =  ( wr_addr ) == ( bv_8_58_n185 )  ;
assign n11586 =  ( n11584 ) & (n11585 )  ;
assign n11587 =  ( n11586 ) & (wr )  ;
assign n11588 =  ( n11587 ) ? ( bv_8_0_n69 ) : ( iram_58 ) ;
assign n11589 = wr_addr[7:7] ;
assign n11590 =  ( n11589 ) == ( bv_1_0_n53 )  ;
assign n11591 =  ( wr_addr ) == ( bv_8_58_n185 )  ;
assign n11592 =  ( n11590 ) & (n11591 )  ;
assign n11593 =  ( n11592 ) & (wr )  ;
assign n11594 =  ( n11593 ) ? ( n5071 ) : ( iram_58 ) ;
assign n11595 = wr_addr[7:7] ;
assign n11596 =  ( n11595 ) == ( bv_1_0_n53 )  ;
assign n11597 =  ( wr_addr ) == ( bv_8_58_n185 )  ;
assign n11598 =  ( n11596 ) & (n11597 )  ;
assign n11599 =  ( n11598 ) & (wr )  ;
assign n11600 =  ( n11599 ) ? ( n5096 ) : ( iram_58 ) ;
assign n11601 = wr_addr[7:7] ;
assign n11602 =  ( n11601 ) == ( bv_1_0_n53 )  ;
assign n11603 =  ( wr_addr ) == ( bv_8_58_n185 )  ;
assign n11604 =  ( n11602 ) & (n11603 )  ;
assign n11605 =  ( n11604 ) & (wr )  ;
assign n11606 =  ( n11605 ) ? ( n5123 ) : ( iram_58 ) ;
assign n11607 = wr_addr[7:7] ;
assign n11608 =  ( n11607 ) == ( bv_1_0_n53 )  ;
assign n11609 =  ( wr_addr ) == ( bv_8_58_n185 )  ;
assign n11610 =  ( n11608 ) & (n11609 )  ;
assign n11611 =  ( n11610 ) & (wr )  ;
assign n11612 =  ( n11611 ) ? ( n5165 ) : ( iram_58 ) ;
assign n11613 = wr_addr[7:7] ;
assign n11614 =  ( n11613 ) == ( bv_1_0_n53 )  ;
assign n11615 =  ( wr_addr ) == ( bv_8_58_n185 )  ;
assign n11616 =  ( n11614 ) & (n11615 )  ;
assign n11617 =  ( n11616 ) & (wr )  ;
assign n11618 =  ( n11617 ) ? ( n5204 ) : ( iram_58 ) ;
assign n11619 = wr_addr[7:7] ;
assign n11620 =  ( n11619 ) == ( bv_1_0_n53 )  ;
assign n11621 =  ( wr_addr ) == ( bv_8_58_n185 )  ;
assign n11622 =  ( n11620 ) & (n11621 )  ;
assign n11623 =  ( n11622 ) & (wr )  ;
assign n11624 =  ( n11623 ) ? ( n5262 ) : ( iram_58 ) ;
assign n11625 = wr_addr[7:7] ;
assign n11626 =  ( n11625 ) == ( bv_1_0_n53 )  ;
assign n11627 =  ( wr_addr ) == ( bv_8_58_n185 )  ;
assign n11628 =  ( n11626 ) & (n11627 )  ;
assign n11629 =  ( n11628 ) & (wr )  ;
assign n11630 =  ( n11629 ) ? ( n5298 ) : ( iram_58 ) ;
assign n11631 = wr_addr[7:7] ;
assign n11632 =  ( n11631 ) == ( bv_1_0_n53 )  ;
assign n11633 =  ( wr_addr ) == ( bv_8_58_n185 )  ;
assign n11634 =  ( n11632 ) & (n11633 )  ;
assign n11635 =  ( n11634 ) & (wr )  ;
assign n11636 =  ( n11635 ) ? ( n5325 ) : ( iram_58 ) ;
assign n11637 = wr_addr[7:7] ;
assign n11638 =  ( n11637 ) == ( bv_1_0_n53 )  ;
assign n11639 =  ( wr_addr ) == ( bv_8_59_n187 )  ;
assign n11640 =  ( n11638 ) & (n11639 )  ;
assign n11641 =  ( n11640 ) & (wr )  ;
assign n11642 =  ( n11641 ) ? ( n4782 ) : ( iram_59 ) ;
assign n11643 = wr_addr[7:7] ;
assign n11644 =  ( n11643 ) == ( bv_1_0_n53 )  ;
assign n11645 =  ( wr_addr ) == ( bv_8_59_n187 )  ;
assign n11646 =  ( n11644 ) & (n11645 )  ;
assign n11647 =  ( n11646 ) & (wr )  ;
assign n11648 =  ( n11647 ) ? ( n4841 ) : ( iram_59 ) ;
assign n11649 = wr_addr[7:7] ;
assign n11650 =  ( n11649 ) == ( bv_1_0_n53 )  ;
assign n11651 =  ( wr_addr ) == ( bv_8_59_n187 )  ;
assign n11652 =  ( n11650 ) & (n11651 )  ;
assign n11653 =  ( n11652 ) & (wr )  ;
assign n11654 =  ( n11653 ) ? ( n5449 ) : ( iram_59 ) ;
assign n11655 = wr_addr[7:7] ;
assign n11656 =  ( n11655 ) == ( bv_1_0_n53 )  ;
assign n11657 =  ( wr_addr ) == ( bv_8_59_n187 )  ;
assign n11658 =  ( n11656 ) & (n11657 )  ;
assign n11659 =  ( n11658 ) & (wr )  ;
assign n11660 =  ( n11659 ) ? ( n4906 ) : ( iram_59 ) ;
assign n11661 = wr_addr[7:7] ;
assign n11662 =  ( n11661 ) == ( bv_1_0_n53 )  ;
assign n11663 =  ( wr_addr ) == ( bv_8_59_n187 )  ;
assign n11664 =  ( n11662 ) & (n11663 )  ;
assign n11665 =  ( n11664 ) & (wr )  ;
assign n11666 =  ( n11665 ) ? ( n5485 ) : ( iram_59 ) ;
assign n11667 = wr_addr[7:7] ;
assign n11668 =  ( n11667 ) == ( bv_1_0_n53 )  ;
assign n11669 =  ( wr_addr ) == ( bv_8_59_n187 )  ;
assign n11670 =  ( n11668 ) & (n11669 )  ;
assign n11671 =  ( n11670 ) & (wr )  ;
assign n11672 =  ( n11671 ) ? ( n5512 ) : ( iram_59 ) ;
assign n11673 = wr_addr[7:7] ;
assign n11674 =  ( n11673 ) == ( bv_1_0_n53 )  ;
assign n11675 =  ( wr_addr ) == ( bv_8_59_n187 )  ;
assign n11676 =  ( n11674 ) & (n11675 )  ;
assign n11677 =  ( n11676 ) & (wr )  ;
assign n11678 =  ( n11677 ) ? ( bv_8_0_n69 ) : ( iram_59 ) ;
assign n11679 = wr_addr[7:7] ;
assign n11680 =  ( n11679 ) == ( bv_1_0_n53 )  ;
assign n11681 =  ( wr_addr ) == ( bv_8_59_n187 )  ;
assign n11682 =  ( n11680 ) & (n11681 )  ;
assign n11683 =  ( n11682 ) & (wr )  ;
assign n11684 =  ( n11683 ) ? ( n5071 ) : ( iram_59 ) ;
assign n11685 = wr_addr[7:7] ;
assign n11686 =  ( n11685 ) == ( bv_1_0_n53 )  ;
assign n11687 =  ( wr_addr ) == ( bv_8_59_n187 )  ;
assign n11688 =  ( n11686 ) & (n11687 )  ;
assign n11689 =  ( n11688 ) & (wr )  ;
assign n11690 =  ( n11689 ) ? ( n5096 ) : ( iram_59 ) ;
assign n11691 = wr_addr[7:7] ;
assign n11692 =  ( n11691 ) == ( bv_1_0_n53 )  ;
assign n11693 =  ( wr_addr ) == ( bv_8_59_n187 )  ;
assign n11694 =  ( n11692 ) & (n11693 )  ;
assign n11695 =  ( n11694 ) & (wr )  ;
assign n11696 =  ( n11695 ) ? ( n5123 ) : ( iram_59 ) ;
assign n11697 = wr_addr[7:7] ;
assign n11698 =  ( n11697 ) == ( bv_1_0_n53 )  ;
assign n11699 =  ( wr_addr ) == ( bv_8_59_n187 )  ;
assign n11700 =  ( n11698 ) & (n11699 )  ;
assign n11701 =  ( n11700 ) & (wr )  ;
assign n11702 =  ( n11701 ) ? ( n5165 ) : ( iram_59 ) ;
assign n11703 = wr_addr[7:7] ;
assign n11704 =  ( n11703 ) == ( bv_1_0_n53 )  ;
assign n11705 =  ( wr_addr ) == ( bv_8_59_n187 )  ;
assign n11706 =  ( n11704 ) & (n11705 )  ;
assign n11707 =  ( n11706 ) & (wr )  ;
assign n11708 =  ( n11707 ) ? ( n5204 ) : ( iram_59 ) ;
assign n11709 = wr_addr[7:7] ;
assign n11710 =  ( n11709 ) == ( bv_1_0_n53 )  ;
assign n11711 =  ( wr_addr ) == ( bv_8_59_n187 )  ;
assign n11712 =  ( n11710 ) & (n11711 )  ;
assign n11713 =  ( n11712 ) & (wr )  ;
assign n11714 =  ( n11713 ) ? ( n5262 ) : ( iram_59 ) ;
assign n11715 = wr_addr[7:7] ;
assign n11716 =  ( n11715 ) == ( bv_1_0_n53 )  ;
assign n11717 =  ( wr_addr ) == ( bv_8_59_n187 )  ;
assign n11718 =  ( n11716 ) & (n11717 )  ;
assign n11719 =  ( n11718 ) & (wr )  ;
assign n11720 =  ( n11719 ) ? ( n5298 ) : ( iram_59 ) ;
assign n11721 = wr_addr[7:7] ;
assign n11722 =  ( n11721 ) == ( bv_1_0_n53 )  ;
assign n11723 =  ( wr_addr ) == ( bv_8_59_n187 )  ;
assign n11724 =  ( n11722 ) & (n11723 )  ;
assign n11725 =  ( n11724 ) & (wr )  ;
assign n11726 =  ( n11725 ) ? ( n5325 ) : ( iram_59 ) ;
assign n11727 = wr_addr[7:7] ;
assign n11728 =  ( n11727 ) == ( bv_1_0_n53 )  ;
assign n11729 =  ( wr_addr ) == ( bv_8_60_n189 )  ;
assign n11730 =  ( n11728 ) & (n11729 )  ;
assign n11731 =  ( n11730 ) & (wr )  ;
assign n11732 =  ( n11731 ) ? ( n4782 ) : ( iram_60 ) ;
assign n11733 = wr_addr[7:7] ;
assign n11734 =  ( n11733 ) == ( bv_1_0_n53 )  ;
assign n11735 =  ( wr_addr ) == ( bv_8_60_n189 )  ;
assign n11736 =  ( n11734 ) & (n11735 )  ;
assign n11737 =  ( n11736 ) & (wr )  ;
assign n11738 =  ( n11737 ) ? ( n4841 ) : ( iram_60 ) ;
assign n11739 = wr_addr[7:7] ;
assign n11740 =  ( n11739 ) == ( bv_1_0_n53 )  ;
assign n11741 =  ( wr_addr ) == ( bv_8_60_n189 )  ;
assign n11742 =  ( n11740 ) & (n11741 )  ;
assign n11743 =  ( n11742 ) & (wr )  ;
assign n11744 =  ( n11743 ) ? ( n5449 ) : ( iram_60 ) ;
assign n11745 = wr_addr[7:7] ;
assign n11746 =  ( n11745 ) == ( bv_1_0_n53 )  ;
assign n11747 =  ( wr_addr ) == ( bv_8_60_n189 )  ;
assign n11748 =  ( n11746 ) & (n11747 )  ;
assign n11749 =  ( n11748 ) & (wr )  ;
assign n11750 =  ( n11749 ) ? ( n4906 ) : ( iram_60 ) ;
assign n11751 = wr_addr[7:7] ;
assign n11752 =  ( n11751 ) == ( bv_1_0_n53 )  ;
assign n11753 =  ( wr_addr ) == ( bv_8_60_n189 )  ;
assign n11754 =  ( n11752 ) & (n11753 )  ;
assign n11755 =  ( n11754 ) & (wr )  ;
assign n11756 =  ( n11755 ) ? ( n5485 ) : ( iram_60 ) ;
assign n11757 = wr_addr[7:7] ;
assign n11758 =  ( n11757 ) == ( bv_1_0_n53 )  ;
assign n11759 =  ( wr_addr ) == ( bv_8_60_n189 )  ;
assign n11760 =  ( n11758 ) & (n11759 )  ;
assign n11761 =  ( n11760 ) & (wr )  ;
assign n11762 =  ( n11761 ) ? ( n5512 ) : ( iram_60 ) ;
assign n11763 = wr_addr[7:7] ;
assign n11764 =  ( n11763 ) == ( bv_1_0_n53 )  ;
assign n11765 =  ( wr_addr ) == ( bv_8_60_n189 )  ;
assign n11766 =  ( n11764 ) & (n11765 )  ;
assign n11767 =  ( n11766 ) & (wr )  ;
assign n11768 =  ( n11767 ) ? ( bv_8_0_n69 ) : ( iram_60 ) ;
assign n11769 = wr_addr[7:7] ;
assign n11770 =  ( n11769 ) == ( bv_1_0_n53 )  ;
assign n11771 =  ( wr_addr ) == ( bv_8_60_n189 )  ;
assign n11772 =  ( n11770 ) & (n11771 )  ;
assign n11773 =  ( n11772 ) & (wr )  ;
assign n11774 =  ( n11773 ) ? ( n5071 ) : ( iram_60 ) ;
assign n11775 = wr_addr[7:7] ;
assign n11776 =  ( n11775 ) == ( bv_1_0_n53 )  ;
assign n11777 =  ( wr_addr ) == ( bv_8_60_n189 )  ;
assign n11778 =  ( n11776 ) & (n11777 )  ;
assign n11779 =  ( n11778 ) & (wr )  ;
assign n11780 =  ( n11779 ) ? ( n5096 ) : ( iram_60 ) ;
assign n11781 = wr_addr[7:7] ;
assign n11782 =  ( n11781 ) == ( bv_1_0_n53 )  ;
assign n11783 =  ( wr_addr ) == ( bv_8_60_n189 )  ;
assign n11784 =  ( n11782 ) & (n11783 )  ;
assign n11785 =  ( n11784 ) & (wr )  ;
assign n11786 =  ( n11785 ) ? ( n5123 ) : ( iram_60 ) ;
assign n11787 = wr_addr[7:7] ;
assign n11788 =  ( n11787 ) == ( bv_1_0_n53 )  ;
assign n11789 =  ( wr_addr ) == ( bv_8_60_n189 )  ;
assign n11790 =  ( n11788 ) & (n11789 )  ;
assign n11791 =  ( n11790 ) & (wr )  ;
assign n11792 =  ( n11791 ) ? ( n5165 ) : ( iram_60 ) ;
assign n11793 = wr_addr[7:7] ;
assign n11794 =  ( n11793 ) == ( bv_1_0_n53 )  ;
assign n11795 =  ( wr_addr ) == ( bv_8_60_n189 )  ;
assign n11796 =  ( n11794 ) & (n11795 )  ;
assign n11797 =  ( n11796 ) & (wr )  ;
assign n11798 =  ( n11797 ) ? ( n5204 ) : ( iram_60 ) ;
assign n11799 = wr_addr[7:7] ;
assign n11800 =  ( n11799 ) == ( bv_1_0_n53 )  ;
assign n11801 =  ( wr_addr ) == ( bv_8_60_n189 )  ;
assign n11802 =  ( n11800 ) & (n11801 )  ;
assign n11803 =  ( n11802 ) & (wr )  ;
assign n11804 =  ( n11803 ) ? ( n5262 ) : ( iram_60 ) ;
assign n11805 = wr_addr[7:7] ;
assign n11806 =  ( n11805 ) == ( bv_1_0_n53 )  ;
assign n11807 =  ( wr_addr ) == ( bv_8_60_n189 )  ;
assign n11808 =  ( n11806 ) & (n11807 )  ;
assign n11809 =  ( n11808 ) & (wr )  ;
assign n11810 =  ( n11809 ) ? ( n5298 ) : ( iram_60 ) ;
assign n11811 = wr_addr[7:7] ;
assign n11812 =  ( n11811 ) == ( bv_1_0_n53 )  ;
assign n11813 =  ( wr_addr ) == ( bv_8_60_n189 )  ;
assign n11814 =  ( n11812 ) & (n11813 )  ;
assign n11815 =  ( n11814 ) & (wr )  ;
assign n11816 =  ( n11815 ) ? ( n5325 ) : ( iram_60 ) ;
assign n11817 = wr_addr[7:7] ;
assign n11818 =  ( n11817 ) == ( bv_1_0_n53 )  ;
assign n11819 =  ( wr_addr ) == ( bv_8_61_n191 )  ;
assign n11820 =  ( n11818 ) & (n11819 )  ;
assign n11821 =  ( n11820 ) & (wr )  ;
assign n11822 =  ( n11821 ) ? ( n4782 ) : ( iram_61 ) ;
assign n11823 = wr_addr[7:7] ;
assign n11824 =  ( n11823 ) == ( bv_1_0_n53 )  ;
assign n11825 =  ( wr_addr ) == ( bv_8_61_n191 )  ;
assign n11826 =  ( n11824 ) & (n11825 )  ;
assign n11827 =  ( n11826 ) & (wr )  ;
assign n11828 =  ( n11827 ) ? ( n4841 ) : ( iram_61 ) ;
assign n11829 = wr_addr[7:7] ;
assign n11830 =  ( n11829 ) == ( bv_1_0_n53 )  ;
assign n11831 =  ( wr_addr ) == ( bv_8_61_n191 )  ;
assign n11832 =  ( n11830 ) & (n11831 )  ;
assign n11833 =  ( n11832 ) & (wr )  ;
assign n11834 =  ( n11833 ) ? ( n5449 ) : ( iram_61 ) ;
assign n11835 = wr_addr[7:7] ;
assign n11836 =  ( n11835 ) == ( bv_1_0_n53 )  ;
assign n11837 =  ( wr_addr ) == ( bv_8_61_n191 )  ;
assign n11838 =  ( n11836 ) & (n11837 )  ;
assign n11839 =  ( n11838 ) & (wr )  ;
assign n11840 =  ( n11839 ) ? ( n4906 ) : ( iram_61 ) ;
assign n11841 = wr_addr[7:7] ;
assign n11842 =  ( n11841 ) == ( bv_1_0_n53 )  ;
assign n11843 =  ( wr_addr ) == ( bv_8_61_n191 )  ;
assign n11844 =  ( n11842 ) & (n11843 )  ;
assign n11845 =  ( n11844 ) & (wr )  ;
assign n11846 =  ( n11845 ) ? ( n5485 ) : ( iram_61 ) ;
assign n11847 = wr_addr[7:7] ;
assign n11848 =  ( n11847 ) == ( bv_1_0_n53 )  ;
assign n11849 =  ( wr_addr ) == ( bv_8_61_n191 )  ;
assign n11850 =  ( n11848 ) & (n11849 )  ;
assign n11851 =  ( n11850 ) & (wr )  ;
assign n11852 =  ( n11851 ) ? ( n5512 ) : ( iram_61 ) ;
assign n11853 = wr_addr[7:7] ;
assign n11854 =  ( n11853 ) == ( bv_1_0_n53 )  ;
assign n11855 =  ( wr_addr ) == ( bv_8_61_n191 )  ;
assign n11856 =  ( n11854 ) & (n11855 )  ;
assign n11857 =  ( n11856 ) & (wr )  ;
assign n11858 =  ( n11857 ) ? ( bv_8_0_n69 ) : ( iram_61 ) ;
assign n11859 = wr_addr[7:7] ;
assign n11860 =  ( n11859 ) == ( bv_1_0_n53 )  ;
assign n11861 =  ( wr_addr ) == ( bv_8_61_n191 )  ;
assign n11862 =  ( n11860 ) & (n11861 )  ;
assign n11863 =  ( n11862 ) & (wr )  ;
assign n11864 =  ( n11863 ) ? ( n5071 ) : ( iram_61 ) ;
assign n11865 = wr_addr[7:7] ;
assign n11866 =  ( n11865 ) == ( bv_1_0_n53 )  ;
assign n11867 =  ( wr_addr ) == ( bv_8_61_n191 )  ;
assign n11868 =  ( n11866 ) & (n11867 )  ;
assign n11869 =  ( n11868 ) & (wr )  ;
assign n11870 =  ( n11869 ) ? ( n5096 ) : ( iram_61 ) ;
assign n11871 = wr_addr[7:7] ;
assign n11872 =  ( n11871 ) == ( bv_1_0_n53 )  ;
assign n11873 =  ( wr_addr ) == ( bv_8_61_n191 )  ;
assign n11874 =  ( n11872 ) & (n11873 )  ;
assign n11875 =  ( n11874 ) & (wr )  ;
assign n11876 =  ( n11875 ) ? ( n5123 ) : ( iram_61 ) ;
assign n11877 = wr_addr[7:7] ;
assign n11878 =  ( n11877 ) == ( bv_1_0_n53 )  ;
assign n11879 =  ( wr_addr ) == ( bv_8_61_n191 )  ;
assign n11880 =  ( n11878 ) & (n11879 )  ;
assign n11881 =  ( n11880 ) & (wr )  ;
assign n11882 =  ( n11881 ) ? ( n5165 ) : ( iram_61 ) ;
assign n11883 = wr_addr[7:7] ;
assign n11884 =  ( n11883 ) == ( bv_1_0_n53 )  ;
assign n11885 =  ( wr_addr ) == ( bv_8_61_n191 )  ;
assign n11886 =  ( n11884 ) & (n11885 )  ;
assign n11887 =  ( n11886 ) & (wr )  ;
assign n11888 =  ( n11887 ) ? ( n5204 ) : ( iram_61 ) ;
assign n11889 = wr_addr[7:7] ;
assign n11890 =  ( n11889 ) == ( bv_1_0_n53 )  ;
assign n11891 =  ( wr_addr ) == ( bv_8_61_n191 )  ;
assign n11892 =  ( n11890 ) & (n11891 )  ;
assign n11893 =  ( n11892 ) & (wr )  ;
assign n11894 =  ( n11893 ) ? ( n5262 ) : ( iram_61 ) ;
assign n11895 = wr_addr[7:7] ;
assign n11896 =  ( n11895 ) == ( bv_1_0_n53 )  ;
assign n11897 =  ( wr_addr ) == ( bv_8_61_n191 )  ;
assign n11898 =  ( n11896 ) & (n11897 )  ;
assign n11899 =  ( n11898 ) & (wr )  ;
assign n11900 =  ( n11899 ) ? ( n5298 ) : ( iram_61 ) ;
assign n11901 = wr_addr[7:7] ;
assign n11902 =  ( n11901 ) == ( bv_1_0_n53 )  ;
assign n11903 =  ( wr_addr ) == ( bv_8_61_n191 )  ;
assign n11904 =  ( n11902 ) & (n11903 )  ;
assign n11905 =  ( n11904 ) & (wr )  ;
assign n11906 =  ( n11905 ) ? ( n5325 ) : ( iram_61 ) ;
assign n11907 = wr_addr[7:7] ;
assign n11908 =  ( n11907 ) == ( bv_1_0_n53 )  ;
assign n11909 =  ( wr_addr ) == ( bv_8_62_n193 )  ;
assign n11910 =  ( n11908 ) & (n11909 )  ;
assign n11911 =  ( n11910 ) & (wr )  ;
assign n11912 =  ( n11911 ) ? ( n4782 ) : ( iram_62 ) ;
assign n11913 = wr_addr[7:7] ;
assign n11914 =  ( n11913 ) == ( bv_1_0_n53 )  ;
assign n11915 =  ( wr_addr ) == ( bv_8_62_n193 )  ;
assign n11916 =  ( n11914 ) & (n11915 )  ;
assign n11917 =  ( n11916 ) & (wr )  ;
assign n11918 =  ( n11917 ) ? ( n4841 ) : ( iram_62 ) ;
assign n11919 = wr_addr[7:7] ;
assign n11920 =  ( n11919 ) == ( bv_1_0_n53 )  ;
assign n11921 =  ( wr_addr ) == ( bv_8_62_n193 )  ;
assign n11922 =  ( n11920 ) & (n11921 )  ;
assign n11923 =  ( n11922 ) & (wr )  ;
assign n11924 =  ( n11923 ) ? ( n5449 ) : ( iram_62 ) ;
assign n11925 = wr_addr[7:7] ;
assign n11926 =  ( n11925 ) == ( bv_1_0_n53 )  ;
assign n11927 =  ( wr_addr ) == ( bv_8_62_n193 )  ;
assign n11928 =  ( n11926 ) & (n11927 )  ;
assign n11929 =  ( n11928 ) & (wr )  ;
assign n11930 =  ( n11929 ) ? ( n4906 ) : ( iram_62 ) ;
assign n11931 = wr_addr[7:7] ;
assign n11932 =  ( n11931 ) == ( bv_1_0_n53 )  ;
assign n11933 =  ( wr_addr ) == ( bv_8_62_n193 )  ;
assign n11934 =  ( n11932 ) & (n11933 )  ;
assign n11935 =  ( n11934 ) & (wr )  ;
assign n11936 =  ( n11935 ) ? ( n5485 ) : ( iram_62 ) ;
assign n11937 = wr_addr[7:7] ;
assign n11938 =  ( n11937 ) == ( bv_1_0_n53 )  ;
assign n11939 =  ( wr_addr ) == ( bv_8_62_n193 )  ;
assign n11940 =  ( n11938 ) & (n11939 )  ;
assign n11941 =  ( n11940 ) & (wr )  ;
assign n11942 =  ( n11941 ) ? ( n5512 ) : ( iram_62 ) ;
assign n11943 = wr_addr[7:7] ;
assign n11944 =  ( n11943 ) == ( bv_1_0_n53 )  ;
assign n11945 =  ( wr_addr ) == ( bv_8_62_n193 )  ;
assign n11946 =  ( n11944 ) & (n11945 )  ;
assign n11947 =  ( n11946 ) & (wr )  ;
assign n11948 =  ( n11947 ) ? ( bv_8_0_n69 ) : ( iram_62 ) ;
assign n11949 = wr_addr[7:7] ;
assign n11950 =  ( n11949 ) == ( bv_1_0_n53 )  ;
assign n11951 =  ( wr_addr ) == ( bv_8_62_n193 )  ;
assign n11952 =  ( n11950 ) & (n11951 )  ;
assign n11953 =  ( n11952 ) & (wr )  ;
assign n11954 =  ( n11953 ) ? ( n5071 ) : ( iram_62 ) ;
assign n11955 = wr_addr[7:7] ;
assign n11956 =  ( n11955 ) == ( bv_1_0_n53 )  ;
assign n11957 =  ( wr_addr ) == ( bv_8_62_n193 )  ;
assign n11958 =  ( n11956 ) & (n11957 )  ;
assign n11959 =  ( n11958 ) & (wr )  ;
assign n11960 =  ( n11959 ) ? ( n5096 ) : ( iram_62 ) ;
assign n11961 = wr_addr[7:7] ;
assign n11962 =  ( n11961 ) == ( bv_1_0_n53 )  ;
assign n11963 =  ( wr_addr ) == ( bv_8_62_n193 )  ;
assign n11964 =  ( n11962 ) & (n11963 )  ;
assign n11965 =  ( n11964 ) & (wr )  ;
assign n11966 =  ( n11965 ) ? ( n5123 ) : ( iram_62 ) ;
assign n11967 = wr_addr[7:7] ;
assign n11968 =  ( n11967 ) == ( bv_1_0_n53 )  ;
assign n11969 =  ( wr_addr ) == ( bv_8_62_n193 )  ;
assign n11970 =  ( n11968 ) & (n11969 )  ;
assign n11971 =  ( n11970 ) & (wr )  ;
assign n11972 =  ( n11971 ) ? ( n5165 ) : ( iram_62 ) ;
assign n11973 = wr_addr[7:7] ;
assign n11974 =  ( n11973 ) == ( bv_1_0_n53 )  ;
assign n11975 =  ( wr_addr ) == ( bv_8_62_n193 )  ;
assign n11976 =  ( n11974 ) & (n11975 )  ;
assign n11977 =  ( n11976 ) & (wr )  ;
assign n11978 =  ( n11977 ) ? ( n5204 ) : ( iram_62 ) ;
assign n11979 = wr_addr[7:7] ;
assign n11980 =  ( n11979 ) == ( bv_1_0_n53 )  ;
assign n11981 =  ( wr_addr ) == ( bv_8_62_n193 )  ;
assign n11982 =  ( n11980 ) & (n11981 )  ;
assign n11983 =  ( n11982 ) & (wr )  ;
assign n11984 =  ( n11983 ) ? ( n5262 ) : ( iram_62 ) ;
assign n11985 = wr_addr[7:7] ;
assign n11986 =  ( n11985 ) == ( bv_1_0_n53 )  ;
assign n11987 =  ( wr_addr ) == ( bv_8_62_n193 )  ;
assign n11988 =  ( n11986 ) & (n11987 )  ;
assign n11989 =  ( n11988 ) & (wr )  ;
assign n11990 =  ( n11989 ) ? ( n5298 ) : ( iram_62 ) ;
assign n11991 = wr_addr[7:7] ;
assign n11992 =  ( n11991 ) == ( bv_1_0_n53 )  ;
assign n11993 =  ( wr_addr ) == ( bv_8_62_n193 )  ;
assign n11994 =  ( n11992 ) & (n11993 )  ;
assign n11995 =  ( n11994 ) & (wr )  ;
assign n11996 =  ( n11995 ) ? ( n5325 ) : ( iram_62 ) ;
assign n11997 = wr_addr[7:7] ;
assign n11998 =  ( n11997 ) == ( bv_1_0_n53 )  ;
assign n11999 =  ( wr_addr ) == ( bv_8_63_n195 )  ;
assign n12000 =  ( n11998 ) & (n11999 )  ;
assign n12001 =  ( n12000 ) & (wr )  ;
assign n12002 =  ( n12001 ) ? ( n4782 ) : ( iram_63 ) ;
assign n12003 = wr_addr[7:7] ;
assign n12004 =  ( n12003 ) == ( bv_1_0_n53 )  ;
assign n12005 =  ( wr_addr ) == ( bv_8_63_n195 )  ;
assign n12006 =  ( n12004 ) & (n12005 )  ;
assign n12007 =  ( n12006 ) & (wr )  ;
assign n12008 =  ( n12007 ) ? ( n4841 ) : ( iram_63 ) ;
assign n12009 = wr_addr[7:7] ;
assign n12010 =  ( n12009 ) == ( bv_1_0_n53 )  ;
assign n12011 =  ( wr_addr ) == ( bv_8_63_n195 )  ;
assign n12012 =  ( n12010 ) & (n12011 )  ;
assign n12013 =  ( n12012 ) & (wr )  ;
assign n12014 =  ( n12013 ) ? ( n5449 ) : ( iram_63 ) ;
assign n12015 = wr_addr[7:7] ;
assign n12016 =  ( n12015 ) == ( bv_1_0_n53 )  ;
assign n12017 =  ( wr_addr ) == ( bv_8_63_n195 )  ;
assign n12018 =  ( n12016 ) & (n12017 )  ;
assign n12019 =  ( n12018 ) & (wr )  ;
assign n12020 =  ( n12019 ) ? ( n4906 ) : ( iram_63 ) ;
assign n12021 = wr_addr[7:7] ;
assign n12022 =  ( n12021 ) == ( bv_1_0_n53 )  ;
assign n12023 =  ( wr_addr ) == ( bv_8_63_n195 )  ;
assign n12024 =  ( n12022 ) & (n12023 )  ;
assign n12025 =  ( n12024 ) & (wr )  ;
assign n12026 =  ( n12025 ) ? ( n5485 ) : ( iram_63 ) ;
assign n12027 = wr_addr[7:7] ;
assign n12028 =  ( n12027 ) == ( bv_1_0_n53 )  ;
assign n12029 =  ( wr_addr ) == ( bv_8_63_n195 )  ;
assign n12030 =  ( n12028 ) & (n12029 )  ;
assign n12031 =  ( n12030 ) & (wr )  ;
assign n12032 =  ( n12031 ) ? ( n5512 ) : ( iram_63 ) ;
assign n12033 = wr_addr[7:7] ;
assign n12034 =  ( n12033 ) == ( bv_1_0_n53 )  ;
assign n12035 =  ( wr_addr ) == ( bv_8_63_n195 )  ;
assign n12036 =  ( n12034 ) & (n12035 )  ;
assign n12037 =  ( n12036 ) & (wr )  ;
assign n12038 =  ( n12037 ) ? ( bv_8_0_n69 ) : ( iram_63 ) ;
assign n12039 = wr_addr[7:7] ;
assign n12040 =  ( n12039 ) == ( bv_1_0_n53 )  ;
assign n12041 =  ( wr_addr ) == ( bv_8_63_n195 )  ;
assign n12042 =  ( n12040 ) & (n12041 )  ;
assign n12043 =  ( n12042 ) & (wr )  ;
assign n12044 =  ( n12043 ) ? ( n5071 ) : ( iram_63 ) ;
assign n12045 = wr_addr[7:7] ;
assign n12046 =  ( n12045 ) == ( bv_1_0_n53 )  ;
assign n12047 =  ( wr_addr ) == ( bv_8_63_n195 )  ;
assign n12048 =  ( n12046 ) & (n12047 )  ;
assign n12049 =  ( n12048 ) & (wr )  ;
assign n12050 =  ( n12049 ) ? ( n5096 ) : ( iram_63 ) ;
assign n12051 = wr_addr[7:7] ;
assign n12052 =  ( n12051 ) == ( bv_1_0_n53 )  ;
assign n12053 =  ( wr_addr ) == ( bv_8_63_n195 )  ;
assign n12054 =  ( n12052 ) & (n12053 )  ;
assign n12055 =  ( n12054 ) & (wr )  ;
assign n12056 =  ( n12055 ) ? ( n5123 ) : ( iram_63 ) ;
assign n12057 = wr_addr[7:7] ;
assign n12058 =  ( n12057 ) == ( bv_1_0_n53 )  ;
assign n12059 =  ( wr_addr ) == ( bv_8_63_n195 )  ;
assign n12060 =  ( n12058 ) & (n12059 )  ;
assign n12061 =  ( n12060 ) & (wr )  ;
assign n12062 =  ( n12061 ) ? ( n5165 ) : ( iram_63 ) ;
assign n12063 = wr_addr[7:7] ;
assign n12064 =  ( n12063 ) == ( bv_1_0_n53 )  ;
assign n12065 =  ( wr_addr ) == ( bv_8_63_n195 )  ;
assign n12066 =  ( n12064 ) & (n12065 )  ;
assign n12067 =  ( n12066 ) & (wr )  ;
assign n12068 =  ( n12067 ) ? ( n5204 ) : ( iram_63 ) ;
assign n12069 = wr_addr[7:7] ;
assign n12070 =  ( n12069 ) == ( bv_1_0_n53 )  ;
assign n12071 =  ( wr_addr ) == ( bv_8_63_n195 )  ;
assign n12072 =  ( n12070 ) & (n12071 )  ;
assign n12073 =  ( n12072 ) & (wr )  ;
assign n12074 =  ( n12073 ) ? ( n5262 ) : ( iram_63 ) ;
assign n12075 = wr_addr[7:7] ;
assign n12076 =  ( n12075 ) == ( bv_1_0_n53 )  ;
assign n12077 =  ( wr_addr ) == ( bv_8_63_n195 )  ;
assign n12078 =  ( n12076 ) & (n12077 )  ;
assign n12079 =  ( n12078 ) & (wr )  ;
assign n12080 =  ( n12079 ) ? ( n5298 ) : ( iram_63 ) ;
assign n12081 = wr_addr[7:7] ;
assign n12082 =  ( n12081 ) == ( bv_1_0_n53 )  ;
assign n12083 =  ( wr_addr ) == ( bv_8_63_n195 )  ;
assign n12084 =  ( n12082 ) & (n12083 )  ;
assign n12085 =  ( n12084 ) & (wr )  ;
assign n12086 =  ( n12085 ) ? ( n5325 ) : ( iram_63 ) ;
assign n12087 = wr_addr[7:7] ;
assign n12088 =  ( n12087 ) == ( bv_1_0_n53 )  ;
assign n12089 =  ( wr_addr ) == ( bv_8_64_n197 )  ;
assign n12090 =  ( n12088 ) & (n12089 )  ;
assign n12091 =  ( n12090 ) & (wr )  ;
assign n12092 =  ( n12091 ) ? ( n4782 ) : ( iram_64 ) ;
assign n12093 = wr_addr[7:7] ;
assign n12094 =  ( n12093 ) == ( bv_1_0_n53 )  ;
assign n12095 =  ( wr_addr ) == ( bv_8_64_n197 )  ;
assign n12096 =  ( n12094 ) & (n12095 )  ;
assign n12097 =  ( n12096 ) & (wr )  ;
assign n12098 =  ( n12097 ) ? ( n4841 ) : ( iram_64 ) ;
assign n12099 = wr_addr[7:7] ;
assign n12100 =  ( n12099 ) == ( bv_1_0_n53 )  ;
assign n12101 =  ( wr_addr ) == ( bv_8_64_n197 )  ;
assign n12102 =  ( n12100 ) & (n12101 )  ;
assign n12103 =  ( n12102 ) & (wr )  ;
assign n12104 =  ( n12103 ) ? ( n5449 ) : ( iram_64 ) ;
assign n12105 = wr_addr[7:7] ;
assign n12106 =  ( n12105 ) == ( bv_1_0_n53 )  ;
assign n12107 =  ( wr_addr ) == ( bv_8_64_n197 )  ;
assign n12108 =  ( n12106 ) & (n12107 )  ;
assign n12109 =  ( n12108 ) & (wr )  ;
assign n12110 =  ( n12109 ) ? ( n4906 ) : ( iram_64 ) ;
assign n12111 = wr_addr[7:7] ;
assign n12112 =  ( n12111 ) == ( bv_1_0_n53 )  ;
assign n12113 =  ( wr_addr ) == ( bv_8_64_n197 )  ;
assign n12114 =  ( n12112 ) & (n12113 )  ;
assign n12115 =  ( n12114 ) & (wr )  ;
assign n12116 =  ( n12115 ) ? ( n5485 ) : ( iram_64 ) ;
assign n12117 = wr_addr[7:7] ;
assign n12118 =  ( n12117 ) == ( bv_1_0_n53 )  ;
assign n12119 =  ( wr_addr ) == ( bv_8_64_n197 )  ;
assign n12120 =  ( n12118 ) & (n12119 )  ;
assign n12121 =  ( n12120 ) & (wr )  ;
assign n12122 =  ( n12121 ) ? ( n5512 ) : ( iram_64 ) ;
assign n12123 = wr_addr[7:7] ;
assign n12124 =  ( n12123 ) == ( bv_1_0_n53 )  ;
assign n12125 =  ( wr_addr ) == ( bv_8_64_n197 )  ;
assign n12126 =  ( n12124 ) & (n12125 )  ;
assign n12127 =  ( n12126 ) & (wr )  ;
assign n12128 =  ( n12127 ) ? ( bv_8_0_n69 ) : ( iram_64 ) ;
assign n12129 = wr_addr[7:7] ;
assign n12130 =  ( n12129 ) == ( bv_1_0_n53 )  ;
assign n12131 =  ( wr_addr ) == ( bv_8_64_n197 )  ;
assign n12132 =  ( n12130 ) & (n12131 )  ;
assign n12133 =  ( n12132 ) & (wr )  ;
assign n12134 =  ( n12133 ) ? ( n5071 ) : ( iram_64 ) ;
assign n12135 = wr_addr[7:7] ;
assign n12136 =  ( n12135 ) == ( bv_1_0_n53 )  ;
assign n12137 =  ( wr_addr ) == ( bv_8_64_n197 )  ;
assign n12138 =  ( n12136 ) & (n12137 )  ;
assign n12139 =  ( n12138 ) & (wr )  ;
assign n12140 =  ( n12139 ) ? ( n5096 ) : ( iram_64 ) ;
assign n12141 = wr_addr[7:7] ;
assign n12142 =  ( n12141 ) == ( bv_1_0_n53 )  ;
assign n12143 =  ( wr_addr ) == ( bv_8_64_n197 )  ;
assign n12144 =  ( n12142 ) & (n12143 )  ;
assign n12145 =  ( n12144 ) & (wr )  ;
assign n12146 =  ( n12145 ) ? ( n5123 ) : ( iram_64 ) ;
assign n12147 = wr_addr[7:7] ;
assign n12148 =  ( n12147 ) == ( bv_1_0_n53 )  ;
assign n12149 =  ( wr_addr ) == ( bv_8_64_n197 )  ;
assign n12150 =  ( n12148 ) & (n12149 )  ;
assign n12151 =  ( n12150 ) & (wr )  ;
assign n12152 =  ( n12151 ) ? ( n5165 ) : ( iram_64 ) ;
assign n12153 = wr_addr[7:7] ;
assign n12154 =  ( n12153 ) == ( bv_1_0_n53 )  ;
assign n12155 =  ( wr_addr ) == ( bv_8_64_n197 )  ;
assign n12156 =  ( n12154 ) & (n12155 )  ;
assign n12157 =  ( n12156 ) & (wr )  ;
assign n12158 =  ( n12157 ) ? ( n5204 ) : ( iram_64 ) ;
assign n12159 = wr_addr[7:7] ;
assign n12160 =  ( n12159 ) == ( bv_1_0_n53 )  ;
assign n12161 =  ( wr_addr ) == ( bv_8_64_n197 )  ;
assign n12162 =  ( n12160 ) & (n12161 )  ;
assign n12163 =  ( n12162 ) & (wr )  ;
assign n12164 =  ( n12163 ) ? ( n5262 ) : ( iram_64 ) ;
assign n12165 = wr_addr[7:7] ;
assign n12166 =  ( n12165 ) == ( bv_1_0_n53 )  ;
assign n12167 =  ( wr_addr ) == ( bv_8_64_n197 )  ;
assign n12168 =  ( n12166 ) & (n12167 )  ;
assign n12169 =  ( n12168 ) & (wr )  ;
assign n12170 =  ( n12169 ) ? ( n5298 ) : ( iram_64 ) ;
assign n12171 = wr_addr[7:7] ;
assign n12172 =  ( n12171 ) == ( bv_1_0_n53 )  ;
assign n12173 =  ( wr_addr ) == ( bv_8_64_n197 )  ;
assign n12174 =  ( n12172 ) & (n12173 )  ;
assign n12175 =  ( n12174 ) & (wr )  ;
assign n12176 =  ( n12175 ) ? ( n5325 ) : ( iram_64 ) ;
assign n12177 = wr_addr[7:7] ;
assign n12178 =  ( n12177 ) == ( bv_1_0_n53 )  ;
assign n12179 =  ( wr_addr ) == ( bv_8_65_n199 )  ;
assign n12180 =  ( n12178 ) & (n12179 )  ;
assign n12181 =  ( n12180 ) & (wr )  ;
assign n12182 =  ( n12181 ) ? ( n4782 ) : ( iram_65 ) ;
assign n12183 = wr_addr[7:7] ;
assign n12184 =  ( n12183 ) == ( bv_1_0_n53 )  ;
assign n12185 =  ( wr_addr ) == ( bv_8_65_n199 )  ;
assign n12186 =  ( n12184 ) & (n12185 )  ;
assign n12187 =  ( n12186 ) & (wr )  ;
assign n12188 =  ( n12187 ) ? ( n4841 ) : ( iram_65 ) ;
assign n12189 = wr_addr[7:7] ;
assign n12190 =  ( n12189 ) == ( bv_1_0_n53 )  ;
assign n12191 =  ( wr_addr ) == ( bv_8_65_n199 )  ;
assign n12192 =  ( n12190 ) & (n12191 )  ;
assign n12193 =  ( n12192 ) & (wr )  ;
assign n12194 =  ( n12193 ) ? ( n5449 ) : ( iram_65 ) ;
assign n12195 = wr_addr[7:7] ;
assign n12196 =  ( n12195 ) == ( bv_1_0_n53 )  ;
assign n12197 =  ( wr_addr ) == ( bv_8_65_n199 )  ;
assign n12198 =  ( n12196 ) & (n12197 )  ;
assign n12199 =  ( n12198 ) & (wr )  ;
assign n12200 =  ( n12199 ) ? ( n4906 ) : ( iram_65 ) ;
assign n12201 = wr_addr[7:7] ;
assign n12202 =  ( n12201 ) == ( bv_1_0_n53 )  ;
assign n12203 =  ( wr_addr ) == ( bv_8_65_n199 )  ;
assign n12204 =  ( n12202 ) & (n12203 )  ;
assign n12205 =  ( n12204 ) & (wr )  ;
assign n12206 =  ( n12205 ) ? ( n5485 ) : ( iram_65 ) ;
assign n12207 = wr_addr[7:7] ;
assign n12208 =  ( n12207 ) == ( bv_1_0_n53 )  ;
assign n12209 =  ( wr_addr ) == ( bv_8_65_n199 )  ;
assign n12210 =  ( n12208 ) & (n12209 )  ;
assign n12211 =  ( n12210 ) & (wr )  ;
assign n12212 =  ( n12211 ) ? ( n5512 ) : ( iram_65 ) ;
assign n12213 = wr_addr[7:7] ;
assign n12214 =  ( n12213 ) == ( bv_1_0_n53 )  ;
assign n12215 =  ( wr_addr ) == ( bv_8_65_n199 )  ;
assign n12216 =  ( n12214 ) & (n12215 )  ;
assign n12217 =  ( n12216 ) & (wr )  ;
assign n12218 =  ( n12217 ) ? ( bv_8_0_n69 ) : ( iram_65 ) ;
assign n12219 = wr_addr[7:7] ;
assign n12220 =  ( n12219 ) == ( bv_1_0_n53 )  ;
assign n12221 =  ( wr_addr ) == ( bv_8_65_n199 )  ;
assign n12222 =  ( n12220 ) & (n12221 )  ;
assign n12223 =  ( n12222 ) & (wr )  ;
assign n12224 =  ( n12223 ) ? ( n5071 ) : ( iram_65 ) ;
assign n12225 = wr_addr[7:7] ;
assign n12226 =  ( n12225 ) == ( bv_1_0_n53 )  ;
assign n12227 =  ( wr_addr ) == ( bv_8_65_n199 )  ;
assign n12228 =  ( n12226 ) & (n12227 )  ;
assign n12229 =  ( n12228 ) & (wr )  ;
assign n12230 =  ( n12229 ) ? ( n5096 ) : ( iram_65 ) ;
assign n12231 = wr_addr[7:7] ;
assign n12232 =  ( n12231 ) == ( bv_1_0_n53 )  ;
assign n12233 =  ( wr_addr ) == ( bv_8_65_n199 )  ;
assign n12234 =  ( n12232 ) & (n12233 )  ;
assign n12235 =  ( n12234 ) & (wr )  ;
assign n12236 =  ( n12235 ) ? ( n5123 ) : ( iram_65 ) ;
assign n12237 = wr_addr[7:7] ;
assign n12238 =  ( n12237 ) == ( bv_1_0_n53 )  ;
assign n12239 =  ( wr_addr ) == ( bv_8_65_n199 )  ;
assign n12240 =  ( n12238 ) & (n12239 )  ;
assign n12241 =  ( n12240 ) & (wr )  ;
assign n12242 =  ( n12241 ) ? ( n5165 ) : ( iram_65 ) ;
assign n12243 = wr_addr[7:7] ;
assign n12244 =  ( n12243 ) == ( bv_1_0_n53 )  ;
assign n12245 =  ( wr_addr ) == ( bv_8_65_n199 )  ;
assign n12246 =  ( n12244 ) & (n12245 )  ;
assign n12247 =  ( n12246 ) & (wr )  ;
assign n12248 =  ( n12247 ) ? ( n5204 ) : ( iram_65 ) ;
assign n12249 = wr_addr[7:7] ;
assign n12250 =  ( n12249 ) == ( bv_1_0_n53 )  ;
assign n12251 =  ( wr_addr ) == ( bv_8_65_n199 )  ;
assign n12252 =  ( n12250 ) & (n12251 )  ;
assign n12253 =  ( n12252 ) & (wr )  ;
assign n12254 =  ( n12253 ) ? ( n5262 ) : ( iram_65 ) ;
assign n12255 = wr_addr[7:7] ;
assign n12256 =  ( n12255 ) == ( bv_1_0_n53 )  ;
assign n12257 =  ( wr_addr ) == ( bv_8_65_n199 )  ;
assign n12258 =  ( n12256 ) & (n12257 )  ;
assign n12259 =  ( n12258 ) & (wr )  ;
assign n12260 =  ( n12259 ) ? ( n5298 ) : ( iram_65 ) ;
assign n12261 = wr_addr[7:7] ;
assign n12262 =  ( n12261 ) == ( bv_1_0_n53 )  ;
assign n12263 =  ( wr_addr ) == ( bv_8_65_n199 )  ;
assign n12264 =  ( n12262 ) & (n12263 )  ;
assign n12265 =  ( n12264 ) & (wr )  ;
assign n12266 =  ( n12265 ) ? ( n5325 ) : ( iram_65 ) ;
assign n12267 = wr_addr[7:7] ;
assign n12268 =  ( n12267 ) == ( bv_1_0_n53 )  ;
assign n12269 =  ( wr_addr ) == ( bv_8_66_n201 )  ;
assign n12270 =  ( n12268 ) & (n12269 )  ;
assign n12271 =  ( n12270 ) & (wr )  ;
assign n12272 =  ( n12271 ) ? ( n4782 ) : ( iram_66 ) ;
assign n12273 = wr_addr[7:7] ;
assign n12274 =  ( n12273 ) == ( bv_1_0_n53 )  ;
assign n12275 =  ( wr_addr ) == ( bv_8_66_n201 )  ;
assign n12276 =  ( n12274 ) & (n12275 )  ;
assign n12277 =  ( n12276 ) & (wr )  ;
assign n12278 =  ( n12277 ) ? ( n4841 ) : ( iram_66 ) ;
assign n12279 = wr_addr[7:7] ;
assign n12280 =  ( n12279 ) == ( bv_1_0_n53 )  ;
assign n12281 =  ( wr_addr ) == ( bv_8_66_n201 )  ;
assign n12282 =  ( n12280 ) & (n12281 )  ;
assign n12283 =  ( n12282 ) & (wr )  ;
assign n12284 =  ( n12283 ) ? ( n5449 ) : ( iram_66 ) ;
assign n12285 = wr_addr[7:7] ;
assign n12286 =  ( n12285 ) == ( bv_1_0_n53 )  ;
assign n12287 =  ( wr_addr ) == ( bv_8_66_n201 )  ;
assign n12288 =  ( n12286 ) & (n12287 )  ;
assign n12289 =  ( n12288 ) & (wr )  ;
assign n12290 =  ( n12289 ) ? ( n4906 ) : ( iram_66 ) ;
assign n12291 = wr_addr[7:7] ;
assign n12292 =  ( n12291 ) == ( bv_1_0_n53 )  ;
assign n12293 =  ( wr_addr ) == ( bv_8_66_n201 )  ;
assign n12294 =  ( n12292 ) & (n12293 )  ;
assign n12295 =  ( n12294 ) & (wr )  ;
assign n12296 =  ( n12295 ) ? ( n5485 ) : ( iram_66 ) ;
assign n12297 = wr_addr[7:7] ;
assign n12298 =  ( n12297 ) == ( bv_1_0_n53 )  ;
assign n12299 =  ( wr_addr ) == ( bv_8_66_n201 )  ;
assign n12300 =  ( n12298 ) & (n12299 )  ;
assign n12301 =  ( n12300 ) & (wr )  ;
assign n12302 =  ( n12301 ) ? ( n5512 ) : ( iram_66 ) ;
assign n12303 = wr_addr[7:7] ;
assign n12304 =  ( n12303 ) == ( bv_1_0_n53 )  ;
assign n12305 =  ( wr_addr ) == ( bv_8_66_n201 )  ;
assign n12306 =  ( n12304 ) & (n12305 )  ;
assign n12307 =  ( n12306 ) & (wr )  ;
assign n12308 =  ( n12307 ) ? ( bv_8_0_n69 ) : ( iram_66 ) ;
assign n12309 = wr_addr[7:7] ;
assign n12310 =  ( n12309 ) == ( bv_1_0_n53 )  ;
assign n12311 =  ( wr_addr ) == ( bv_8_66_n201 )  ;
assign n12312 =  ( n12310 ) & (n12311 )  ;
assign n12313 =  ( n12312 ) & (wr )  ;
assign n12314 =  ( n12313 ) ? ( n5071 ) : ( iram_66 ) ;
assign n12315 = wr_addr[7:7] ;
assign n12316 =  ( n12315 ) == ( bv_1_0_n53 )  ;
assign n12317 =  ( wr_addr ) == ( bv_8_66_n201 )  ;
assign n12318 =  ( n12316 ) & (n12317 )  ;
assign n12319 =  ( n12318 ) & (wr )  ;
assign n12320 =  ( n12319 ) ? ( n5096 ) : ( iram_66 ) ;
assign n12321 = wr_addr[7:7] ;
assign n12322 =  ( n12321 ) == ( bv_1_0_n53 )  ;
assign n12323 =  ( wr_addr ) == ( bv_8_66_n201 )  ;
assign n12324 =  ( n12322 ) & (n12323 )  ;
assign n12325 =  ( n12324 ) & (wr )  ;
assign n12326 =  ( n12325 ) ? ( n5123 ) : ( iram_66 ) ;
assign n12327 = wr_addr[7:7] ;
assign n12328 =  ( n12327 ) == ( bv_1_0_n53 )  ;
assign n12329 =  ( wr_addr ) == ( bv_8_66_n201 )  ;
assign n12330 =  ( n12328 ) & (n12329 )  ;
assign n12331 =  ( n12330 ) & (wr )  ;
assign n12332 =  ( n12331 ) ? ( n5165 ) : ( iram_66 ) ;
assign n12333 = wr_addr[7:7] ;
assign n12334 =  ( n12333 ) == ( bv_1_0_n53 )  ;
assign n12335 =  ( wr_addr ) == ( bv_8_66_n201 )  ;
assign n12336 =  ( n12334 ) & (n12335 )  ;
assign n12337 =  ( n12336 ) & (wr )  ;
assign n12338 =  ( n12337 ) ? ( n5204 ) : ( iram_66 ) ;
assign n12339 = wr_addr[7:7] ;
assign n12340 =  ( n12339 ) == ( bv_1_0_n53 )  ;
assign n12341 =  ( wr_addr ) == ( bv_8_66_n201 )  ;
assign n12342 =  ( n12340 ) & (n12341 )  ;
assign n12343 =  ( n12342 ) & (wr )  ;
assign n12344 =  ( n12343 ) ? ( n5262 ) : ( iram_66 ) ;
assign n12345 = wr_addr[7:7] ;
assign n12346 =  ( n12345 ) == ( bv_1_0_n53 )  ;
assign n12347 =  ( wr_addr ) == ( bv_8_66_n201 )  ;
assign n12348 =  ( n12346 ) & (n12347 )  ;
assign n12349 =  ( n12348 ) & (wr )  ;
assign n12350 =  ( n12349 ) ? ( n5298 ) : ( iram_66 ) ;
assign n12351 = wr_addr[7:7] ;
assign n12352 =  ( n12351 ) == ( bv_1_0_n53 )  ;
assign n12353 =  ( wr_addr ) == ( bv_8_66_n201 )  ;
assign n12354 =  ( n12352 ) & (n12353 )  ;
assign n12355 =  ( n12354 ) & (wr )  ;
assign n12356 =  ( n12355 ) ? ( n5325 ) : ( iram_66 ) ;
assign n12357 = wr_addr[7:7] ;
assign n12358 =  ( n12357 ) == ( bv_1_0_n53 )  ;
assign n12359 =  ( wr_addr ) == ( bv_8_67_n203 )  ;
assign n12360 =  ( n12358 ) & (n12359 )  ;
assign n12361 =  ( n12360 ) & (wr )  ;
assign n12362 =  ( n12361 ) ? ( n4782 ) : ( iram_67 ) ;
assign n12363 = wr_addr[7:7] ;
assign n12364 =  ( n12363 ) == ( bv_1_0_n53 )  ;
assign n12365 =  ( wr_addr ) == ( bv_8_67_n203 )  ;
assign n12366 =  ( n12364 ) & (n12365 )  ;
assign n12367 =  ( n12366 ) & (wr )  ;
assign n12368 =  ( n12367 ) ? ( n4841 ) : ( iram_67 ) ;
assign n12369 = wr_addr[7:7] ;
assign n12370 =  ( n12369 ) == ( bv_1_0_n53 )  ;
assign n12371 =  ( wr_addr ) == ( bv_8_67_n203 )  ;
assign n12372 =  ( n12370 ) & (n12371 )  ;
assign n12373 =  ( n12372 ) & (wr )  ;
assign n12374 =  ( n12373 ) ? ( n5449 ) : ( iram_67 ) ;
assign n12375 = wr_addr[7:7] ;
assign n12376 =  ( n12375 ) == ( bv_1_0_n53 )  ;
assign n12377 =  ( wr_addr ) == ( bv_8_67_n203 )  ;
assign n12378 =  ( n12376 ) & (n12377 )  ;
assign n12379 =  ( n12378 ) & (wr )  ;
assign n12380 =  ( n12379 ) ? ( n4906 ) : ( iram_67 ) ;
assign n12381 = wr_addr[7:7] ;
assign n12382 =  ( n12381 ) == ( bv_1_0_n53 )  ;
assign n12383 =  ( wr_addr ) == ( bv_8_67_n203 )  ;
assign n12384 =  ( n12382 ) & (n12383 )  ;
assign n12385 =  ( n12384 ) & (wr )  ;
assign n12386 =  ( n12385 ) ? ( n5485 ) : ( iram_67 ) ;
assign n12387 = wr_addr[7:7] ;
assign n12388 =  ( n12387 ) == ( bv_1_0_n53 )  ;
assign n12389 =  ( wr_addr ) == ( bv_8_67_n203 )  ;
assign n12390 =  ( n12388 ) & (n12389 )  ;
assign n12391 =  ( n12390 ) & (wr )  ;
assign n12392 =  ( n12391 ) ? ( n5512 ) : ( iram_67 ) ;
assign n12393 = wr_addr[7:7] ;
assign n12394 =  ( n12393 ) == ( bv_1_0_n53 )  ;
assign n12395 =  ( wr_addr ) == ( bv_8_67_n203 )  ;
assign n12396 =  ( n12394 ) & (n12395 )  ;
assign n12397 =  ( n12396 ) & (wr )  ;
assign n12398 =  ( n12397 ) ? ( bv_8_0_n69 ) : ( iram_67 ) ;
assign n12399 = wr_addr[7:7] ;
assign n12400 =  ( n12399 ) == ( bv_1_0_n53 )  ;
assign n12401 =  ( wr_addr ) == ( bv_8_67_n203 )  ;
assign n12402 =  ( n12400 ) & (n12401 )  ;
assign n12403 =  ( n12402 ) & (wr )  ;
assign n12404 =  ( n12403 ) ? ( n5071 ) : ( iram_67 ) ;
assign n12405 = wr_addr[7:7] ;
assign n12406 =  ( n12405 ) == ( bv_1_0_n53 )  ;
assign n12407 =  ( wr_addr ) == ( bv_8_67_n203 )  ;
assign n12408 =  ( n12406 ) & (n12407 )  ;
assign n12409 =  ( n12408 ) & (wr )  ;
assign n12410 =  ( n12409 ) ? ( n5096 ) : ( iram_67 ) ;
assign n12411 = wr_addr[7:7] ;
assign n12412 =  ( n12411 ) == ( bv_1_0_n53 )  ;
assign n12413 =  ( wr_addr ) == ( bv_8_67_n203 )  ;
assign n12414 =  ( n12412 ) & (n12413 )  ;
assign n12415 =  ( n12414 ) & (wr )  ;
assign n12416 =  ( n12415 ) ? ( n5123 ) : ( iram_67 ) ;
assign n12417 = wr_addr[7:7] ;
assign n12418 =  ( n12417 ) == ( bv_1_0_n53 )  ;
assign n12419 =  ( wr_addr ) == ( bv_8_67_n203 )  ;
assign n12420 =  ( n12418 ) & (n12419 )  ;
assign n12421 =  ( n12420 ) & (wr )  ;
assign n12422 =  ( n12421 ) ? ( n5165 ) : ( iram_67 ) ;
assign n12423 = wr_addr[7:7] ;
assign n12424 =  ( n12423 ) == ( bv_1_0_n53 )  ;
assign n12425 =  ( wr_addr ) == ( bv_8_67_n203 )  ;
assign n12426 =  ( n12424 ) & (n12425 )  ;
assign n12427 =  ( n12426 ) & (wr )  ;
assign n12428 =  ( n12427 ) ? ( n5204 ) : ( iram_67 ) ;
assign n12429 = wr_addr[7:7] ;
assign n12430 =  ( n12429 ) == ( bv_1_0_n53 )  ;
assign n12431 =  ( wr_addr ) == ( bv_8_67_n203 )  ;
assign n12432 =  ( n12430 ) & (n12431 )  ;
assign n12433 =  ( n12432 ) & (wr )  ;
assign n12434 =  ( n12433 ) ? ( n5262 ) : ( iram_67 ) ;
assign n12435 = wr_addr[7:7] ;
assign n12436 =  ( n12435 ) == ( bv_1_0_n53 )  ;
assign n12437 =  ( wr_addr ) == ( bv_8_67_n203 )  ;
assign n12438 =  ( n12436 ) & (n12437 )  ;
assign n12439 =  ( n12438 ) & (wr )  ;
assign n12440 =  ( n12439 ) ? ( n5298 ) : ( iram_67 ) ;
assign n12441 = wr_addr[7:7] ;
assign n12442 =  ( n12441 ) == ( bv_1_0_n53 )  ;
assign n12443 =  ( wr_addr ) == ( bv_8_67_n203 )  ;
assign n12444 =  ( n12442 ) & (n12443 )  ;
assign n12445 =  ( n12444 ) & (wr )  ;
assign n12446 =  ( n12445 ) ? ( n5325 ) : ( iram_67 ) ;
assign n12447 = wr_addr[7:7] ;
assign n12448 =  ( n12447 ) == ( bv_1_0_n53 )  ;
assign n12449 =  ( wr_addr ) == ( bv_8_68_n205 )  ;
assign n12450 =  ( n12448 ) & (n12449 )  ;
assign n12451 =  ( n12450 ) & (wr )  ;
assign n12452 =  ( n12451 ) ? ( n4782 ) : ( iram_68 ) ;
assign n12453 = wr_addr[7:7] ;
assign n12454 =  ( n12453 ) == ( bv_1_0_n53 )  ;
assign n12455 =  ( wr_addr ) == ( bv_8_68_n205 )  ;
assign n12456 =  ( n12454 ) & (n12455 )  ;
assign n12457 =  ( n12456 ) & (wr )  ;
assign n12458 =  ( n12457 ) ? ( n4841 ) : ( iram_68 ) ;
assign n12459 = wr_addr[7:7] ;
assign n12460 =  ( n12459 ) == ( bv_1_0_n53 )  ;
assign n12461 =  ( wr_addr ) == ( bv_8_68_n205 )  ;
assign n12462 =  ( n12460 ) & (n12461 )  ;
assign n12463 =  ( n12462 ) & (wr )  ;
assign n12464 =  ( n12463 ) ? ( n5449 ) : ( iram_68 ) ;
assign n12465 = wr_addr[7:7] ;
assign n12466 =  ( n12465 ) == ( bv_1_0_n53 )  ;
assign n12467 =  ( wr_addr ) == ( bv_8_68_n205 )  ;
assign n12468 =  ( n12466 ) & (n12467 )  ;
assign n12469 =  ( n12468 ) & (wr )  ;
assign n12470 =  ( n12469 ) ? ( n4906 ) : ( iram_68 ) ;
assign n12471 = wr_addr[7:7] ;
assign n12472 =  ( n12471 ) == ( bv_1_0_n53 )  ;
assign n12473 =  ( wr_addr ) == ( bv_8_68_n205 )  ;
assign n12474 =  ( n12472 ) & (n12473 )  ;
assign n12475 =  ( n12474 ) & (wr )  ;
assign n12476 =  ( n12475 ) ? ( n5485 ) : ( iram_68 ) ;
assign n12477 = wr_addr[7:7] ;
assign n12478 =  ( n12477 ) == ( bv_1_0_n53 )  ;
assign n12479 =  ( wr_addr ) == ( bv_8_68_n205 )  ;
assign n12480 =  ( n12478 ) & (n12479 )  ;
assign n12481 =  ( n12480 ) & (wr )  ;
assign n12482 =  ( n12481 ) ? ( n5512 ) : ( iram_68 ) ;
assign n12483 = wr_addr[7:7] ;
assign n12484 =  ( n12483 ) == ( bv_1_0_n53 )  ;
assign n12485 =  ( wr_addr ) == ( bv_8_68_n205 )  ;
assign n12486 =  ( n12484 ) & (n12485 )  ;
assign n12487 =  ( n12486 ) & (wr )  ;
assign n12488 =  ( n12487 ) ? ( bv_8_0_n69 ) : ( iram_68 ) ;
assign n12489 = wr_addr[7:7] ;
assign n12490 =  ( n12489 ) == ( bv_1_0_n53 )  ;
assign n12491 =  ( wr_addr ) == ( bv_8_68_n205 )  ;
assign n12492 =  ( n12490 ) & (n12491 )  ;
assign n12493 =  ( n12492 ) & (wr )  ;
assign n12494 =  ( n12493 ) ? ( n5071 ) : ( iram_68 ) ;
assign n12495 = wr_addr[7:7] ;
assign n12496 =  ( n12495 ) == ( bv_1_0_n53 )  ;
assign n12497 =  ( wr_addr ) == ( bv_8_68_n205 )  ;
assign n12498 =  ( n12496 ) & (n12497 )  ;
assign n12499 =  ( n12498 ) & (wr )  ;
assign n12500 =  ( n12499 ) ? ( n5096 ) : ( iram_68 ) ;
assign n12501 = wr_addr[7:7] ;
assign n12502 =  ( n12501 ) == ( bv_1_0_n53 )  ;
assign n12503 =  ( wr_addr ) == ( bv_8_68_n205 )  ;
assign n12504 =  ( n12502 ) & (n12503 )  ;
assign n12505 =  ( n12504 ) & (wr )  ;
assign n12506 =  ( n12505 ) ? ( n5123 ) : ( iram_68 ) ;
assign n12507 = wr_addr[7:7] ;
assign n12508 =  ( n12507 ) == ( bv_1_0_n53 )  ;
assign n12509 =  ( wr_addr ) == ( bv_8_68_n205 )  ;
assign n12510 =  ( n12508 ) & (n12509 )  ;
assign n12511 =  ( n12510 ) & (wr )  ;
assign n12512 =  ( n12511 ) ? ( n5165 ) : ( iram_68 ) ;
assign n12513 = wr_addr[7:7] ;
assign n12514 =  ( n12513 ) == ( bv_1_0_n53 )  ;
assign n12515 =  ( wr_addr ) == ( bv_8_68_n205 )  ;
assign n12516 =  ( n12514 ) & (n12515 )  ;
assign n12517 =  ( n12516 ) & (wr )  ;
assign n12518 =  ( n12517 ) ? ( n5204 ) : ( iram_68 ) ;
assign n12519 = wr_addr[7:7] ;
assign n12520 =  ( n12519 ) == ( bv_1_0_n53 )  ;
assign n12521 =  ( wr_addr ) == ( bv_8_68_n205 )  ;
assign n12522 =  ( n12520 ) & (n12521 )  ;
assign n12523 =  ( n12522 ) & (wr )  ;
assign n12524 =  ( n12523 ) ? ( n5262 ) : ( iram_68 ) ;
assign n12525 = wr_addr[7:7] ;
assign n12526 =  ( n12525 ) == ( bv_1_0_n53 )  ;
assign n12527 =  ( wr_addr ) == ( bv_8_68_n205 )  ;
assign n12528 =  ( n12526 ) & (n12527 )  ;
assign n12529 =  ( n12528 ) & (wr )  ;
assign n12530 =  ( n12529 ) ? ( n5298 ) : ( iram_68 ) ;
assign n12531 = wr_addr[7:7] ;
assign n12532 =  ( n12531 ) == ( bv_1_0_n53 )  ;
assign n12533 =  ( wr_addr ) == ( bv_8_68_n205 )  ;
assign n12534 =  ( n12532 ) & (n12533 )  ;
assign n12535 =  ( n12534 ) & (wr )  ;
assign n12536 =  ( n12535 ) ? ( n5325 ) : ( iram_68 ) ;
assign n12537 = wr_addr[7:7] ;
assign n12538 =  ( n12537 ) == ( bv_1_0_n53 )  ;
assign n12539 =  ( wr_addr ) == ( bv_8_69_n207 )  ;
assign n12540 =  ( n12538 ) & (n12539 )  ;
assign n12541 =  ( n12540 ) & (wr )  ;
assign n12542 =  ( n12541 ) ? ( n4782 ) : ( iram_69 ) ;
assign n12543 = wr_addr[7:7] ;
assign n12544 =  ( n12543 ) == ( bv_1_0_n53 )  ;
assign n12545 =  ( wr_addr ) == ( bv_8_69_n207 )  ;
assign n12546 =  ( n12544 ) & (n12545 )  ;
assign n12547 =  ( n12546 ) & (wr )  ;
assign n12548 =  ( n12547 ) ? ( n4841 ) : ( iram_69 ) ;
assign n12549 = wr_addr[7:7] ;
assign n12550 =  ( n12549 ) == ( bv_1_0_n53 )  ;
assign n12551 =  ( wr_addr ) == ( bv_8_69_n207 )  ;
assign n12552 =  ( n12550 ) & (n12551 )  ;
assign n12553 =  ( n12552 ) & (wr )  ;
assign n12554 =  ( n12553 ) ? ( n5449 ) : ( iram_69 ) ;
assign n12555 = wr_addr[7:7] ;
assign n12556 =  ( n12555 ) == ( bv_1_0_n53 )  ;
assign n12557 =  ( wr_addr ) == ( bv_8_69_n207 )  ;
assign n12558 =  ( n12556 ) & (n12557 )  ;
assign n12559 =  ( n12558 ) & (wr )  ;
assign n12560 =  ( n12559 ) ? ( n4906 ) : ( iram_69 ) ;
assign n12561 = wr_addr[7:7] ;
assign n12562 =  ( n12561 ) == ( bv_1_0_n53 )  ;
assign n12563 =  ( wr_addr ) == ( bv_8_69_n207 )  ;
assign n12564 =  ( n12562 ) & (n12563 )  ;
assign n12565 =  ( n12564 ) & (wr )  ;
assign n12566 =  ( n12565 ) ? ( n5485 ) : ( iram_69 ) ;
assign n12567 = wr_addr[7:7] ;
assign n12568 =  ( n12567 ) == ( bv_1_0_n53 )  ;
assign n12569 =  ( wr_addr ) == ( bv_8_69_n207 )  ;
assign n12570 =  ( n12568 ) & (n12569 )  ;
assign n12571 =  ( n12570 ) & (wr )  ;
assign n12572 =  ( n12571 ) ? ( n5512 ) : ( iram_69 ) ;
assign n12573 = wr_addr[7:7] ;
assign n12574 =  ( n12573 ) == ( bv_1_0_n53 )  ;
assign n12575 =  ( wr_addr ) == ( bv_8_69_n207 )  ;
assign n12576 =  ( n12574 ) & (n12575 )  ;
assign n12577 =  ( n12576 ) & (wr )  ;
assign n12578 =  ( n12577 ) ? ( bv_8_0_n69 ) : ( iram_69 ) ;
assign n12579 = wr_addr[7:7] ;
assign n12580 =  ( n12579 ) == ( bv_1_0_n53 )  ;
assign n12581 =  ( wr_addr ) == ( bv_8_69_n207 )  ;
assign n12582 =  ( n12580 ) & (n12581 )  ;
assign n12583 =  ( n12582 ) & (wr )  ;
assign n12584 =  ( n12583 ) ? ( n5071 ) : ( iram_69 ) ;
assign n12585 = wr_addr[7:7] ;
assign n12586 =  ( n12585 ) == ( bv_1_0_n53 )  ;
assign n12587 =  ( wr_addr ) == ( bv_8_69_n207 )  ;
assign n12588 =  ( n12586 ) & (n12587 )  ;
assign n12589 =  ( n12588 ) & (wr )  ;
assign n12590 =  ( n12589 ) ? ( n5096 ) : ( iram_69 ) ;
assign n12591 = wr_addr[7:7] ;
assign n12592 =  ( n12591 ) == ( bv_1_0_n53 )  ;
assign n12593 =  ( wr_addr ) == ( bv_8_69_n207 )  ;
assign n12594 =  ( n12592 ) & (n12593 )  ;
assign n12595 =  ( n12594 ) & (wr )  ;
assign n12596 =  ( n12595 ) ? ( n5123 ) : ( iram_69 ) ;
assign n12597 = wr_addr[7:7] ;
assign n12598 =  ( n12597 ) == ( bv_1_0_n53 )  ;
assign n12599 =  ( wr_addr ) == ( bv_8_69_n207 )  ;
assign n12600 =  ( n12598 ) & (n12599 )  ;
assign n12601 =  ( n12600 ) & (wr )  ;
assign n12602 =  ( n12601 ) ? ( n5165 ) : ( iram_69 ) ;
assign n12603 = wr_addr[7:7] ;
assign n12604 =  ( n12603 ) == ( bv_1_0_n53 )  ;
assign n12605 =  ( wr_addr ) == ( bv_8_69_n207 )  ;
assign n12606 =  ( n12604 ) & (n12605 )  ;
assign n12607 =  ( n12606 ) & (wr )  ;
assign n12608 =  ( n12607 ) ? ( n5204 ) : ( iram_69 ) ;
assign n12609 = wr_addr[7:7] ;
assign n12610 =  ( n12609 ) == ( bv_1_0_n53 )  ;
assign n12611 =  ( wr_addr ) == ( bv_8_69_n207 )  ;
assign n12612 =  ( n12610 ) & (n12611 )  ;
assign n12613 =  ( n12612 ) & (wr )  ;
assign n12614 =  ( n12613 ) ? ( n5262 ) : ( iram_69 ) ;
assign n12615 = wr_addr[7:7] ;
assign n12616 =  ( n12615 ) == ( bv_1_0_n53 )  ;
assign n12617 =  ( wr_addr ) == ( bv_8_69_n207 )  ;
assign n12618 =  ( n12616 ) & (n12617 )  ;
assign n12619 =  ( n12618 ) & (wr )  ;
assign n12620 =  ( n12619 ) ? ( n5298 ) : ( iram_69 ) ;
assign n12621 = wr_addr[7:7] ;
assign n12622 =  ( n12621 ) == ( bv_1_0_n53 )  ;
assign n12623 =  ( wr_addr ) == ( bv_8_69_n207 )  ;
assign n12624 =  ( n12622 ) & (n12623 )  ;
assign n12625 =  ( n12624 ) & (wr )  ;
assign n12626 =  ( n12625 ) ? ( n5325 ) : ( iram_69 ) ;
assign n12627 = wr_addr[7:7] ;
assign n12628 =  ( n12627 ) == ( bv_1_0_n53 )  ;
assign n12629 =  ( wr_addr ) == ( bv_8_70_n209 )  ;
assign n12630 =  ( n12628 ) & (n12629 )  ;
assign n12631 =  ( n12630 ) & (wr )  ;
assign n12632 =  ( n12631 ) ? ( n4782 ) : ( iram_70 ) ;
assign n12633 = wr_addr[7:7] ;
assign n12634 =  ( n12633 ) == ( bv_1_0_n53 )  ;
assign n12635 =  ( wr_addr ) == ( bv_8_70_n209 )  ;
assign n12636 =  ( n12634 ) & (n12635 )  ;
assign n12637 =  ( n12636 ) & (wr )  ;
assign n12638 =  ( n12637 ) ? ( n4841 ) : ( iram_70 ) ;
assign n12639 = wr_addr[7:7] ;
assign n12640 =  ( n12639 ) == ( bv_1_0_n53 )  ;
assign n12641 =  ( wr_addr ) == ( bv_8_70_n209 )  ;
assign n12642 =  ( n12640 ) & (n12641 )  ;
assign n12643 =  ( n12642 ) & (wr )  ;
assign n12644 =  ( n12643 ) ? ( n5449 ) : ( iram_70 ) ;
assign n12645 = wr_addr[7:7] ;
assign n12646 =  ( n12645 ) == ( bv_1_0_n53 )  ;
assign n12647 =  ( wr_addr ) == ( bv_8_70_n209 )  ;
assign n12648 =  ( n12646 ) & (n12647 )  ;
assign n12649 =  ( n12648 ) & (wr )  ;
assign n12650 =  ( n12649 ) ? ( n4906 ) : ( iram_70 ) ;
assign n12651 = wr_addr[7:7] ;
assign n12652 =  ( n12651 ) == ( bv_1_0_n53 )  ;
assign n12653 =  ( wr_addr ) == ( bv_8_70_n209 )  ;
assign n12654 =  ( n12652 ) & (n12653 )  ;
assign n12655 =  ( n12654 ) & (wr )  ;
assign n12656 =  ( n12655 ) ? ( n5485 ) : ( iram_70 ) ;
assign n12657 = wr_addr[7:7] ;
assign n12658 =  ( n12657 ) == ( bv_1_0_n53 )  ;
assign n12659 =  ( wr_addr ) == ( bv_8_70_n209 )  ;
assign n12660 =  ( n12658 ) & (n12659 )  ;
assign n12661 =  ( n12660 ) & (wr )  ;
assign n12662 =  ( n12661 ) ? ( n5512 ) : ( iram_70 ) ;
assign n12663 = wr_addr[7:7] ;
assign n12664 =  ( n12663 ) == ( bv_1_0_n53 )  ;
assign n12665 =  ( wr_addr ) == ( bv_8_70_n209 )  ;
assign n12666 =  ( n12664 ) & (n12665 )  ;
assign n12667 =  ( n12666 ) & (wr )  ;
assign n12668 =  ( n12667 ) ? ( bv_8_0_n69 ) : ( iram_70 ) ;
assign n12669 = wr_addr[7:7] ;
assign n12670 =  ( n12669 ) == ( bv_1_0_n53 )  ;
assign n12671 =  ( wr_addr ) == ( bv_8_70_n209 )  ;
assign n12672 =  ( n12670 ) & (n12671 )  ;
assign n12673 =  ( n12672 ) & (wr )  ;
assign n12674 =  ( n12673 ) ? ( n5071 ) : ( iram_70 ) ;
assign n12675 = wr_addr[7:7] ;
assign n12676 =  ( n12675 ) == ( bv_1_0_n53 )  ;
assign n12677 =  ( wr_addr ) == ( bv_8_70_n209 )  ;
assign n12678 =  ( n12676 ) & (n12677 )  ;
assign n12679 =  ( n12678 ) & (wr )  ;
assign n12680 =  ( n12679 ) ? ( n5096 ) : ( iram_70 ) ;
assign n12681 = wr_addr[7:7] ;
assign n12682 =  ( n12681 ) == ( bv_1_0_n53 )  ;
assign n12683 =  ( wr_addr ) == ( bv_8_70_n209 )  ;
assign n12684 =  ( n12682 ) & (n12683 )  ;
assign n12685 =  ( n12684 ) & (wr )  ;
assign n12686 =  ( n12685 ) ? ( n5123 ) : ( iram_70 ) ;
assign n12687 = wr_addr[7:7] ;
assign n12688 =  ( n12687 ) == ( bv_1_0_n53 )  ;
assign n12689 =  ( wr_addr ) == ( bv_8_70_n209 )  ;
assign n12690 =  ( n12688 ) & (n12689 )  ;
assign n12691 =  ( n12690 ) & (wr )  ;
assign n12692 =  ( n12691 ) ? ( n5165 ) : ( iram_70 ) ;
assign n12693 = wr_addr[7:7] ;
assign n12694 =  ( n12693 ) == ( bv_1_0_n53 )  ;
assign n12695 =  ( wr_addr ) == ( bv_8_70_n209 )  ;
assign n12696 =  ( n12694 ) & (n12695 )  ;
assign n12697 =  ( n12696 ) & (wr )  ;
assign n12698 =  ( n12697 ) ? ( n5204 ) : ( iram_70 ) ;
assign n12699 = wr_addr[7:7] ;
assign n12700 =  ( n12699 ) == ( bv_1_0_n53 )  ;
assign n12701 =  ( wr_addr ) == ( bv_8_70_n209 )  ;
assign n12702 =  ( n12700 ) & (n12701 )  ;
assign n12703 =  ( n12702 ) & (wr )  ;
assign n12704 =  ( n12703 ) ? ( n5262 ) : ( iram_70 ) ;
assign n12705 = wr_addr[7:7] ;
assign n12706 =  ( n12705 ) == ( bv_1_0_n53 )  ;
assign n12707 =  ( wr_addr ) == ( bv_8_70_n209 )  ;
assign n12708 =  ( n12706 ) & (n12707 )  ;
assign n12709 =  ( n12708 ) & (wr )  ;
assign n12710 =  ( n12709 ) ? ( n5298 ) : ( iram_70 ) ;
assign n12711 = wr_addr[7:7] ;
assign n12712 =  ( n12711 ) == ( bv_1_0_n53 )  ;
assign n12713 =  ( wr_addr ) == ( bv_8_70_n209 )  ;
assign n12714 =  ( n12712 ) & (n12713 )  ;
assign n12715 =  ( n12714 ) & (wr )  ;
assign n12716 =  ( n12715 ) ? ( n5325 ) : ( iram_70 ) ;
assign n12717 = wr_addr[7:7] ;
assign n12718 =  ( n12717 ) == ( bv_1_0_n53 )  ;
assign n12719 =  ( wr_addr ) == ( bv_8_71_n211 )  ;
assign n12720 =  ( n12718 ) & (n12719 )  ;
assign n12721 =  ( n12720 ) & (wr )  ;
assign n12722 =  ( n12721 ) ? ( n4782 ) : ( iram_71 ) ;
assign n12723 = wr_addr[7:7] ;
assign n12724 =  ( n12723 ) == ( bv_1_0_n53 )  ;
assign n12725 =  ( wr_addr ) == ( bv_8_71_n211 )  ;
assign n12726 =  ( n12724 ) & (n12725 )  ;
assign n12727 =  ( n12726 ) & (wr )  ;
assign n12728 =  ( n12727 ) ? ( n4841 ) : ( iram_71 ) ;
assign n12729 = wr_addr[7:7] ;
assign n12730 =  ( n12729 ) == ( bv_1_0_n53 )  ;
assign n12731 =  ( wr_addr ) == ( bv_8_71_n211 )  ;
assign n12732 =  ( n12730 ) & (n12731 )  ;
assign n12733 =  ( n12732 ) & (wr )  ;
assign n12734 =  ( n12733 ) ? ( n5449 ) : ( iram_71 ) ;
assign n12735 = wr_addr[7:7] ;
assign n12736 =  ( n12735 ) == ( bv_1_0_n53 )  ;
assign n12737 =  ( wr_addr ) == ( bv_8_71_n211 )  ;
assign n12738 =  ( n12736 ) & (n12737 )  ;
assign n12739 =  ( n12738 ) & (wr )  ;
assign n12740 =  ( n12739 ) ? ( n4906 ) : ( iram_71 ) ;
assign n12741 = wr_addr[7:7] ;
assign n12742 =  ( n12741 ) == ( bv_1_0_n53 )  ;
assign n12743 =  ( wr_addr ) == ( bv_8_71_n211 )  ;
assign n12744 =  ( n12742 ) & (n12743 )  ;
assign n12745 =  ( n12744 ) & (wr )  ;
assign n12746 =  ( n12745 ) ? ( n5485 ) : ( iram_71 ) ;
assign n12747 = wr_addr[7:7] ;
assign n12748 =  ( n12747 ) == ( bv_1_0_n53 )  ;
assign n12749 =  ( wr_addr ) == ( bv_8_71_n211 )  ;
assign n12750 =  ( n12748 ) & (n12749 )  ;
assign n12751 =  ( n12750 ) & (wr )  ;
assign n12752 =  ( n12751 ) ? ( n5512 ) : ( iram_71 ) ;
assign n12753 = wr_addr[7:7] ;
assign n12754 =  ( n12753 ) == ( bv_1_0_n53 )  ;
assign n12755 =  ( wr_addr ) == ( bv_8_71_n211 )  ;
assign n12756 =  ( n12754 ) & (n12755 )  ;
assign n12757 =  ( n12756 ) & (wr )  ;
assign n12758 =  ( n12757 ) ? ( bv_8_0_n69 ) : ( iram_71 ) ;
assign n12759 = wr_addr[7:7] ;
assign n12760 =  ( n12759 ) == ( bv_1_0_n53 )  ;
assign n12761 =  ( wr_addr ) == ( bv_8_71_n211 )  ;
assign n12762 =  ( n12760 ) & (n12761 )  ;
assign n12763 =  ( n12762 ) & (wr )  ;
assign n12764 =  ( n12763 ) ? ( n5071 ) : ( iram_71 ) ;
assign n12765 = wr_addr[7:7] ;
assign n12766 =  ( n12765 ) == ( bv_1_0_n53 )  ;
assign n12767 =  ( wr_addr ) == ( bv_8_71_n211 )  ;
assign n12768 =  ( n12766 ) & (n12767 )  ;
assign n12769 =  ( n12768 ) & (wr )  ;
assign n12770 =  ( n12769 ) ? ( n5096 ) : ( iram_71 ) ;
assign n12771 = wr_addr[7:7] ;
assign n12772 =  ( n12771 ) == ( bv_1_0_n53 )  ;
assign n12773 =  ( wr_addr ) == ( bv_8_71_n211 )  ;
assign n12774 =  ( n12772 ) & (n12773 )  ;
assign n12775 =  ( n12774 ) & (wr )  ;
assign n12776 =  ( n12775 ) ? ( n5123 ) : ( iram_71 ) ;
assign n12777 = wr_addr[7:7] ;
assign n12778 =  ( n12777 ) == ( bv_1_0_n53 )  ;
assign n12779 =  ( wr_addr ) == ( bv_8_71_n211 )  ;
assign n12780 =  ( n12778 ) & (n12779 )  ;
assign n12781 =  ( n12780 ) & (wr )  ;
assign n12782 =  ( n12781 ) ? ( n5165 ) : ( iram_71 ) ;
assign n12783 = wr_addr[7:7] ;
assign n12784 =  ( n12783 ) == ( bv_1_0_n53 )  ;
assign n12785 =  ( wr_addr ) == ( bv_8_71_n211 )  ;
assign n12786 =  ( n12784 ) & (n12785 )  ;
assign n12787 =  ( n12786 ) & (wr )  ;
assign n12788 =  ( n12787 ) ? ( n5204 ) : ( iram_71 ) ;
assign n12789 = wr_addr[7:7] ;
assign n12790 =  ( n12789 ) == ( bv_1_0_n53 )  ;
assign n12791 =  ( wr_addr ) == ( bv_8_71_n211 )  ;
assign n12792 =  ( n12790 ) & (n12791 )  ;
assign n12793 =  ( n12792 ) & (wr )  ;
assign n12794 =  ( n12793 ) ? ( n5262 ) : ( iram_71 ) ;
assign n12795 = wr_addr[7:7] ;
assign n12796 =  ( n12795 ) == ( bv_1_0_n53 )  ;
assign n12797 =  ( wr_addr ) == ( bv_8_71_n211 )  ;
assign n12798 =  ( n12796 ) & (n12797 )  ;
assign n12799 =  ( n12798 ) & (wr )  ;
assign n12800 =  ( n12799 ) ? ( n5298 ) : ( iram_71 ) ;
assign n12801 = wr_addr[7:7] ;
assign n12802 =  ( n12801 ) == ( bv_1_0_n53 )  ;
assign n12803 =  ( wr_addr ) == ( bv_8_71_n211 )  ;
assign n12804 =  ( n12802 ) & (n12803 )  ;
assign n12805 =  ( n12804 ) & (wr )  ;
assign n12806 =  ( n12805 ) ? ( n5325 ) : ( iram_71 ) ;
assign n12807 = wr_addr[7:7] ;
assign n12808 =  ( n12807 ) == ( bv_1_0_n53 )  ;
assign n12809 =  ( wr_addr ) == ( bv_8_72_n213 )  ;
assign n12810 =  ( n12808 ) & (n12809 )  ;
assign n12811 =  ( n12810 ) & (wr )  ;
assign n12812 =  ( n12811 ) ? ( n4782 ) : ( iram_72 ) ;
assign n12813 = wr_addr[7:7] ;
assign n12814 =  ( n12813 ) == ( bv_1_0_n53 )  ;
assign n12815 =  ( wr_addr ) == ( bv_8_72_n213 )  ;
assign n12816 =  ( n12814 ) & (n12815 )  ;
assign n12817 =  ( n12816 ) & (wr )  ;
assign n12818 =  ( n12817 ) ? ( n4841 ) : ( iram_72 ) ;
assign n12819 = wr_addr[7:7] ;
assign n12820 =  ( n12819 ) == ( bv_1_0_n53 )  ;
assign n12821 =  ( wr_addr ) == ( bv_8_72_n213 )  ;
assign n12822 =  ( n12820 ) & (n12821 )  ;
assign n12823 =  ( n12822 ) & (wr )  ;
assign n12824 =  ( n12823 ) ? ( n5449 ) : ( iram_72 ) ;
assign n12825 = wr_addr[7:7] ;
assign n12826 =  ( n12825 ) == ( bv_1_0_n53 )  ;
assign n12827 =  ( wr_addr ) == ( bv_8_72_n213 )  ;
assign n12828 =  ( n12826 ) & (n12827 )  ;
assign n12829 =  ( n12828 ) & (wr )  ;
assign n12830 =  ( n12829 ) ? ( n4906 ) : ( iram_72 ) ;
assign n12831 = wr_addr[7:7] ;
assign n12832 =  ( n12831 ) == ( bv_1_0_n53 )  ;
assign n12833 =  ( wr_addr ) == ( bv_8_72_n213 )  ;
assign n12834 =  ( n12832 ) & (n12833 )  ;
assign n12835 =  ( n12834 ) & (wr )  ;
assign n12836 =  ( n12835 ) ? ( n5485 ) : ( iram_72 ) ;
assign n12837 = wr_addr[7:7] ;
assign n12838 =  ( n12837 ) == ( bv_1_0_n53 )  ;
assign n12839 =  ( wr_addr ) == ( bv_8_72_n213 )  ;
assign n12840 =  ( n12838 ) & (n12839 )  ;
assign n12841 =  ( n12840 ) & (wr )  ;
assign n12842 =  ( n12841 ) ? ( n5512 ) : ( iram_72 ) ;
assign n12843 = wr_addr[7:7] ;
assign n12844 =  ( n12843 ) == ( bv_1_0_n53 )  ;
assign n12845 =  ( wr_addr ) == ( bv_8_72_n213 )  ;
assign n12846 =  ( n12844 ) & (n12845 )  ;
assign n12847 =  ( n12846 ) & (wr )  ;
assign n12848 =  ( n12847 ) ? ( bv_8_0_n69 ) : ( iram_72 ) ;
assign n12849 = wr_addr[7:7] ;
assign n12850 =  ( n12849 ) == ( bv_1_0_n53 )  ;
assign n12851 =  ( wr_addr ) == ( bv_8_72_n213 )  ;
assign n12852 =  ( n12850 ) & (n12851 )  ;
assign n12853 =  ( n12852 ) & (wr )  ;
assign n12854 =  ( n12853 ) ? ( n5071 ) : ( iram_72 ) ;
assign n12855 = wr_addr[7:7] ;
assign n12856 =  ( n12855 ) == ( bv_1_0_n53 )  ;
assign n12857 =  ( wr_addr ) == ( bv_8_72_n213 )  ;
assign n12858 =  ( n12856 ) & (n12857 )  ;
assign n12859 =  ( n12858 ) & (wr )  ;
assign n12860 =  ( n12859 ) ? ( n5096 ) : ( iram_72 ) ;
assign n12861 = wr_addr[7:7] ;
assign n12862 =  ( n12861 ) == ( bv_1_0_n53 )  ;
assign n12863 =  ( wr_addr ) == ( bv_8_72_n213 )  ;
assign n12864 =  ( n12862 ) & (n12863 )  ;
assign n12865 =  ( n12864 ) & (wr )  ;
assign n12866 =  ( n12865 ) ? ( n5123 ) : ( iram_72 ) ;
assign n12867 = wr_addr[7:7] ;
assign n12868 =  ( n12867 ) == ( bv_1_0_n53 )  ;
assign n12869 =  ( wr_addr ) == ( bv_8_72_n213 )  ;
assign n12870 =  ( n12868 ) & (n12869 )  ;
assign n12871 =  ( n12870 ) & (wr )  ;
assign n12872 =  ( n12871 ) ? ( n5165 ) : ( iram_72 ) ;
assign n12873 = wr_addr[7:7] ;
assign n12874 =  ( n12873 ) == ( bv_1_0_n53 )  ;
assign n12875 =  ( wr_addr ) == ( bv_8_72_n213 )  ;
assign n12876 =  ( n12874 ) & (n12875 )  ;
assign n12877 =  ( n12876 ) & (wr )  ;
assign n12878 =  ( n12877 ) ? ( n5204 ) : ( iram_72 ) ;
assign n12879 = wr_addr[7:7] ;
assign n12880 =  ( n12879 ) == ( bv_1_0_n53 )  ;
assign n12881 =  ( wr_addr ) == ( bv_8_72_n213 )  ;
assign n12882 =  ( n12880 ) & (n12881 )  ;
assign n12883 =  ( n12882 ) & (wr )  ;
assign n12884 =  ( n12883 ) ? ( n5262 ) : ( iram_72 ) ;
assign n12885 = wr_addr[7:7] ;
assign n12886 =  ( n12885 ) == ( bv_1_0_n53 )  ;
assign n12887 =  ( wr_addr ) == ( bv_8_72_n213 )  ;
assign n12888 =  ( n12886 ) & (n12887 )  ;
assign n12889 =  ( n12888 ) & (wr )  ;
assign n12890 =  ( n12889 ) ? ( n5298 ) : ( iram_72 ) ;
assign n12891 = wr_addr[7:7] ;
assign n12892 =  ( n12891 ) == ( bv_1_0_n53 )  ;
assign n12893 =  ( wr_addr ) == ( bv_8_72_n213 )  ;
assign n12894 =  ( n12892 ) & (n12893 )  ;
assign n12895 =  ( n12894 ) & (wr )  ;
assign n12896 =  ( n12895 ) ? ( n5325 ) : ( iram_72 ) ;
assign n12897 = wr_addr[7:7] ;
assign n12898 =  ( n12897 ) == ( bv_1_0_n53 )  ;
assign n12899 =  ( wr_addr ) == ( bv_8_73_n215 )  ;
assign n12900 =  ( n12898 ) & (n12899 )  ;
assign n12901 =  ( n12900 ) & (wr )  ;
assign n12902 =  ( n12901 ) ? ( n4782 ) : ( iram_73 ) ;
assign n12903 = wr_addr[7:7] ;
assign n12904 =  ( n12903 ) == ( bv_1_0_n53 )  ;
assign n12905 =  ( wr_addr ) == ( bv_8_73_n215 )  ;
assign n12906 =  ( n12904 ) & (n12905 )  ;
assign n12907 =  ( n12906 ) & (wr )  ;
assign n12908 =  ( n12907 ) ? ( n4841 ) : ( iram_73 ) ;
assign n12909 = wr_addr[7:7] ;
assign n12910 =  ( n12909 ) == ( bv_1_0_n53 )  ;
assign n12911 =  ( wr_addr ) == ( bv_8_73_n215 )  ;
assign n12912 =  ( n12910 ) & (n12911 )  ;
assign n12913 =  ( n12912 ) & (wr )  ;
assign n12914 =  ( n12913 ) ? ( n5449 ) : ( iram_73 ) ;
assign n12915 = wr_addr[7:7] ;
assign n12916 =  ( n12915 ) == ( bv_1_0_n53 )  ;
assign n12917 =  ( wr_addr ) == ( bv_8_73_n215 )  ;
assign n12918 =  ( n12916 ) & (n12917 )  ;
assign n12919 =  ( n12918 ) & (wr )  ;
assign n12920 =  ( n12919 ) ? ( n4906 ) : ( iram_73 ) ;
assign n12921 = wr_addr[7:7] ;
assign n12922 =  ( n12921 ) == ( bv_1_0_n53 )  ;
assign n12923 =  ( wr_addr ) == ( bv_8_73_n215 )  ;
assign n12924 =  ( n12922 ) & (n12923 )  ;
assign n12925 =  ( n12924 ) & (wr )  ;
assign n12926 =  ( n12925 ) ? ( n5485 ) : ( iram_73 ) ;
assign n12927 = wr_addr[7:7] ;
assign n12928 =  ( n12927 ) == ( bv_1_0_n53 )  ;
assign n12929 =  ( wr_addr ) == ( bv_8_73_n215 )  ;
assign n12930 =  ( n12928 ) & (n12929 )  ;
assign n12931 =  ( n12930 ) & (wr )  ;
assign n12932 =  ( n12931 ) ? ( n5512 ) : ( iram_73 ) ;
assign n12933 = wr_addr[7:7] ;
assign n12934 =  ( n12933 ) == ( bv_1_0_n53 )  ;
assign n12935 =  ( wr_addr ) == ( bv_8_73_n215 )  ;
assign n12936 =  ( n12934 ) & (n12935 )  ;
assign n12937 =  ( n12936 ) & (wr )  ;
assign n12938 =  ( n12937 ) ? ( bv_8_0_n69 ) : ( iram_73 ) ;
assign n12939 = wr_addr[7:7] ;
assign n12940 =  ( n12939 ) == ( bv_1_0_n53 )  ;
assign n12941 =  ( wr_addr ) == ( bv_8_73_n215 )  ;
assign n12942 =  ( n12940 ) & (n12941 )  ;
assign n12943 =  ( n12942 ) & (wr )  ;
assign n12944 =  ( n12943 ) ? ( n5071 ) : ( iram_73 ) ;
assign n12945 = wr_addr[7:7] ;
assign n12946 =  ( n12945 ) == ( bv_1_0_n53 )  ;
assign n12947 =  ( wr_addr ) == ( bv_8_73_n215 )  ;
assign n12948 =  ( n12946 ) & (n12947 )  ;
assign n12949 =  ( n12948 ) & (wr )  ;
assign n12950 =  ( n12949 ) ? ( n5096 ) : ( iram_73 ) ;
assign n12951 = wr_addr[7:7] ;
assign n12952 =  ( n12951 ) == ( bv_1_0_n53 )  ;
assign n12953 =  ( wr_addr ) == ( bv_8_73_n215 )  ;
assign n12954 =  ( n12952 ) & (n12953 )  ;
assign n12955 =  ( n12954 ) & (wr )  ;
assign n12956 =  ( n12955 ) ? ( n5123 ) : ( iram_73 ) ;
assign n12957 = wr_addr[7:7] ;
assign n12958 =  ( n12957 ) == ( bv_1_0_n53 )  ;
assign n12959 =  ( wr_addr ) == ( bv_8_73_n215 )  ;
assign n12960 =  ( n12958 ) & (n12959 )  ;
assign n12961 =  ( n12960 ) & (wr )  ;
assign n12962 =  ( n12961 ) ? ( n5165 ) : ( iram_73 ) ;
assign n12963 = wr_addr[7:7] ;
assign n12964 =  ( n12963 ) == ( bv_1_0_n53 )  ;
assign n12965 =  ( wr_addr ) == ( bv_8_73_n215 )  ;
assign n12966 =  ( n12964 ) & (n12965 )  ;
assign n12967 =  ( n12966 ) & (wr )  ;
assign n12968 =  ( n12967 ) ? ( n5204 ) : ( iram_73 ) ;
assign n12969 = wr_addr[7:7] ;
assign n12970 =  ( n12969 ) == ( bv_1_0_n53 )  ;
assign n12971 =  ( wr_addr ) == ( bv_8_73_n215 )  ;
assign n12972 =  ( n12970 ) & (n12971 )  ;
assign n12973 =  ( n12972 ) & (wr )  ;
assign n12974 =  ( n12973 ) ? ( n5262 ) : ( iram_73 ) ;
assign n12975 = wr_addr[7:7] ;
assign n12976 =  ( n12975 ) == ( bv_1_0_n53 )  ;
assign n12977 =  ( wr_addr ) == ( bv_8_73_n215 )  ;
assign n12978 =  ( n12976 ) & (n12977 )  ;
assign n12979 =  ( n12978 ) & (wr )  ;
assign n12980 =  ( n12979 ) ? ( n5298 ) : ( iram_73 ) ;
assign n12981 = wr_addr[7:7] ;
assign n12982 =  ( n12981 ) == ( bv_1_0_n53 )  ;
assign n12983 =  ( wr_addr ) == ( bv_8_73_n215 )  ;
assign n12984 =  ( n12982 ) & (n12983 )  ;
assign n12985 =  ( n12984 ) & (wr )  ;
assign n12986 =  ( n12985 ) ? ( n5325 ) : ( iram_73 ) ;
assign n12987 = wr_addr[7:7] ;
assign n12988 =  ( n12987 ) == ( bv_1_0_n53 )  ;
assign n12989 =  ( wr_addr ) == ( bv_8_74_n217 )  ;
assign n12990 =  ( n12988 ) & (n12989 )  ;
assign n12991 =  ( n12990 ) & (wr )  ;
assign n12992 =  ( n12991 ) ? ( n4782 ) : ( iram_74 ) ;
assign n12993 = wr_addr[7:7] ;
assign n12994 =  ( n12993 ) == ( bv_1_0_n53 )  ;
assign n12995 =  ( wr_addr ) == ( bv_8_74_n217 )  ;
assign n12996 =  ( n12994 ) & (n12995 )  ;
assign n12997 =  ( n12996 ) & (wr )  ;
assign n12998 =  ( n12997 ) ? ( n4841 ) : ( iram_74 ) ;
assign n12999 = wr_addr[7:7] ;
assign n13000 =  ( n12999 ) == ( bv_1_0_n53 )  ;
assign n13001 =  ( wr_addr ) == ( bv_8_74_n217 )  ;
assign n13002 =  ( n13000 ) & (n13001 )  ;
assign n13003 =  ( n13002 ) & (wr )  ;
assign n13004 =  ( n13003 ) ? ( n5449 ) : ( iram_74 ) ;
assign n13005 = wr_addr[7:7] ;
assign n13006 =  ( n13005 ) == ( bv_1_0_n53 )  ;
assign n13007 =  ( wr_addr ) == ( bv_8_74_n217 )  ;
assign n13008 =  ( n13006 ) & (n13007 )  ;
assign n13009 =  ( n13008 ) & (wr )  ;
assign n13010 =  ( n13009 ) ? ( n4906 ) : ( iram_74 ) ;
assign n13011 = wr_addr[7:7] ;
assign n13012 =  ( n13011 ) == ( bv_1_0_n53 )  ;
assign n13013 =  ( wr_addr ) == ( bv_8_74_n217 )  ;
assign n13014 =  ( n13012 ) & (n13013 )  ;
assign n13015 =  ( n13014 ) & (wr )  ;
assign n13016 =  ( n13015 ) ? ( n5485 ) : ( iram_74 ) ;
assign n13017 = wr_addr[7:7] ;
assign n13018 =  ( n13017 ) == ( bv_1_0_n53 )  ;
assign n13019 =  ( wr_addr ) == ( bv_8_74_n217 )  ;
assign n13020 =  ( n13018 ) & (n13019 )  ;
assign n13021 =  ( n13020 ) & (wr )  ;
assign n13022 =  ( n13021 ) ? ( n5512 ) : ( iram_74 ) ;
assign n13023 = wr_addr[7:7] ;
assign n13024 =  ( n13023 ) == ( bv_1_0_n53 )  ;
assign n13025 =  ( wr_addr ) == ( bv_8_74_n217 )  ;
assign n13026 =  ( n13024 ) & (n13025 )  ;
assign n13027 =  ( n13026 ) & (wr )  ;
assign n13028 =  ( n13027 ) ? ( bv_8_0_n69 ) : ( iram_74 ) ;
assign n13029 = wr_addr[7:7] ;
assign n13030 =  ( n13029 ) == ( bv_1_0_n53 )  ;
assign n13031 =  ( wr_addr ) == ( bv_8_74_n217 )  ;
assign n13032 =  ( n13030 ) & (n13031 )  ;
assign n13033 =  ( n13032 ) & (wr )  ;
assign n13034 =  ( n13033 ) ? ( n5071 ) : ( iram_74 ) ;
assign n13035 = wr_addr[7:7] ;
assign n13036 =  ( n13035 ) == ( bv_1_0_n53 )  ;
assign n13037 =  ( wr_addr ) == ( bv_8_74_n217 )  ;
assign n13038 =  ( n13036 ) & (n13037 )  ;
assign n13039 =  ( n13038 ) & (wr )  ;
assign n13040 =  ( n13039 ) ? ( n5096 ) : ( iram_74 ) ;
assign n13041 = wr_addr[7:7] ;
assign n13042 =  ( n13041 ) == ( bv_1_0_n53 )  ;
assign n13043 =  ( wr_addr ) == ( bv_8_74_n217 )  ;
assign n13044 =  ( n13042 ) & (n13043 )  ;
assign n13045 =  ( n13044 ) & (wr )  ;
assign n13046 =  ( n13045 ) ? ( n5123 ) : ( iram_74 ) ;
assign n13047 = wr_addr[7:7] ;
assign n13048 =  ( n13047 ) == ( bv_1_0_n53 )  ;
assign n13049 =  ( wr_addr ) == ( bv_8_74_n217 )  ;
assign n13050 =  ( n13048 ) & (n13049 )  ;
assign n13051 =  ( n13050 ) & (wr )  ;
assign n13052 =  ( n13051 ) ? ( n5165 ) : ( iram_74 ) ;
assign n13053 = wr_addr[7:7] ;
assign n13054 =  ( n13053 ) == ( bv_1_0_n53 )  ;
assign n13055 =  ( wr_addr ) == ( bv_8_74_n217 )  ;
assign n13056 =  ( n13054 ) & (n13055 )  ;
assign n13057 =  ( n13056 ) & (wr )  ;
assign n13058 =  ( n13057 ) ? ( n5204 ) : ( iram_74 ) ;
assign n13059 = wr_addr[7:7] ;
assign n13060 =  ( n13059 ) == ( bv_1_0_n53 )  ;
assign n13061 =  ( wr_addr ) == ( bv_8_74_n217 )  ;
assign n13062 =  ( n13060 ) & (n13061 )  ;
assign n13063 =  ( n13062 ) & (wr )  ;
assign n13064 =  ( n13063 ) ? ( n5262 ) : ( iram_74 ) ;
assign n13065 = wr_addr[7:7] ;
assign n13066 =  ( n13065 ) == ( bv_1_0_n53 )  ;
assign n13067 =  ( wr_addr ) == ( bv_8_74_n217 )  ;
assign n13068 =  ( n13066 ) & (n13067 )  ;
assign n13069 =  ( n13068 ) & (wr )  ;
assign n13070 =  ( n13069 ) ? ( n5298 ) : ( iram_74 ) ;
assign n13071 = wr_addr[7:7] ;
assign n13072 =  ( n13071 ) == ( bv_1_0_n53 )  ;
assign n13073 =  ( wr_addr ) == ( bv_8_74_n217 )  ;
assign n13074 =  ( n13072 ) & (n13073 )  ;
assign n13075 =  ( n13074 ) & (wr )  ;
assign n13076 =  ( n13075 ) ? ( n5325 ) : ( iram_74 ) ;
assign n13077 = wr_addr[7:7] ;
assign n13078 =  ( n13077 ) == ( bv_1_0_n53 )  ;
assign n13079 =  ( wr_addr ) == ( bv_8_75_n219 )  ;
assign n13080 =  ( n13078 ) & (n13079 )  ;
assign n13081 =  ( n13080 ) & (wr )  ;
assign n13082 =  ( n13081 ) ? ( n4782 ) : ( iram_75 ) ;
assign n13083 = wr_addr[7:7] ;
assign n13084 =  ( n13083 ) == ( bv_1_0_n53 )  ;
assign n13085 =  ( wr_addr ) == ( bv_8_75_n219 )  ;
assign n13086 =  ( n13084 ) & (n13085 )  ;
assign n13087 =  ( n13086 ) & (wr )  ;
assign n13088 =  ( n13087 ) ? ( n4841 ) : ( iram_75 ) ;
assign n13089 = wr_addr[7:7] ;
assign n13090 =  ( n13089 ) == ( bv_1_0_n53 )  ;
assign n13091 =  ( wr_addr ) == ( bv_8_75_n219 )  ;
assign n13092 =  ( n13090 ) & (n13091 )  ;
assign n13093 =  ( n13092 ) & (wr )  ;
assign n13094 =  ( n13093 ) ? ( n5449 ) : ( iram_75 ) ;
assign n13095 = wr_addr[7:7] ;
assign n13096 =  ( n13095 ) == ( bv_1_0_n53 )  ;
assign n13097 =  ( wr_addr ) == ( bv_8_75_n219 )  ;
assign n13098 =  ( n13096 ) & (n13097 )  ;
assign n13099 =  ( n13098 ) & (wr )  ;
assign n13100 =  ( n13099 ) ? ( n4906 ) : ( iram_75 ) ;
assign n13101 = wr_addr[7:7] ;
assign n13102 =  ( n13101 ) == ( bv_1_0_n53 )  ;
assign n13103 =  ( wr_addr ) == ( bv_8_75_n219 )  ;
assign n13104 =  ( n13102 ) & (n13103 )  ;
assign n13105 =  ( n13104 ) & (wr )  ;
assign n13106 =  ( n13105 ) ? ( n5485 ) : ( iram_75 ) ;
assign n13107 = wr_addr[7:7] ;
assign n13108 =  ( n13107 ) == ( bv_1_0_n53 )  ;
assign n13109 =  ( wr_addr ) == ( bv_8_75_n219 )  ;
assign n13110 =  ( n13108 ) & (n13109 )  ;
assign n13111 =  ( n13110 ) & (wr )  ;
assign n13112 =  ( n13111 ) ? ( n5512 ) : ( iram_75 ) ;
assign n13113 = wr_addr[7:7] ;
assign n13114 =  ( n13113 ) == ( bv_1_0_n53 )  ;
assign n13115 =  ( wr_addr ) == ( bv_8_75_n219 )  ;
assign n13116 =  ( n13114 ) & (n13115 )  ;
assign n13117 =  ( n13116 ) & (wr )  ;
assign n13118 =  ( n13117 ) ? ( bv_8_0_n69 ) : ( iram_75 ) ;
assign n13119 = wr_addr[7:7] ;
assign n13120 =  ( n13119 ) == ( bv_1_0_n53 )  ;
assign n13121 =  ( wr_addr ) == ( bv_8_75_n219 )  ;
assign n13122 =  ( n13120 ) & (n13121 )  ;
assign n13123 =  ( n13122 ) & (wr )  ;
assign n13124 =  ( n13123 ) ? ( n5071 ) : ( iram_75 ) ;
assign n13125 = wr_addr[7:7] ;
assign n13126 =  ( n13125 ) == ( bv_1_0_n53 )  ;
assign n13127 =  ( wr_addr ) == ( bv_8_75_n219 )  ;
assign n13128 =  ( n13126 ) & (n13127 )  ;
assign n13129 =  ( n13128 ) & (wr )  ;
assign n13130 =  ( n13129 ) ? ( n5096 ) : ( iram_75 ) ;
assign n13131 = wr_addr[7:7] ;
assign n13132 =  ( n13131 ) == ( bv_1_0_n53 )  ;
assign n13133 =  ( wr_addr ) == ( bv_8_75_n219 )  ;
assign n13134 =  ( n13132 ) & (n13133 )  ;
assign n13135 =  ( n13134 ) & (wr )  ;
assign n13136 =  ( n13135 ) ? ( n5123 ) : ( iram_75 ) ;
assign n13137 = wr_addr[7:7] ;
assign n13138 =  ( n13137 ) == ( bv_1_0_n53 )  ;
assign n13139 =  ( wr_addr ) == ( bv_8_75_n219 )  ;
assign n13140 =  ( n13138 ) & (n13139 )  ;
assign n13141 =  ( n13140 ) & (wr )  ;
assign n13142 =  ( n13141 ) ? ( n5165 ) : ( iram_75 ) ;
assign n13143 = wr_addr[7:7] ;
assign n13144 =  ( n13143 ) == ( bv_1_0_n53 )  ;
assign n13145 =  ( wr_addr ) == ( bv_8_75_n219 )  ;
assign n13146 =  ( n13144 ) & (n13145 )  ;
assign n13147 =  ( n13146 ) & (wr )  ;
assign n13148 =  ( n13147 ) ? ( n5204 ) : ( iram_75 ) ;
assign n13149 = wr_addr[7:7] ;
assign n13150 =  ( n13149 ) == ( bv_1_0_n53 )  ;
assign n13151 =  ( wr_addr ) == ( bv_8_75_n219 )  ;
assign n13152 =  ( n13150 ) & (n13151 )  ;
assign n13153 =  ( n13152 ) & (wr )  ;
assign n13154 =  ( n13153 ) ? ( n5262 ) : ( iram_75 ) ;
assign n13155 = wr_addr[7:7] ;
assign n13156 =  ( n13155 ) == ( bv_1_0_n53 )  ;
assign n13157 =  ( wr_addr ) == ( bv_8_75_n219 )  ;
assign n13158 =  ( n13156 ) & (n13157 )  ;
assign n13159 =  ( n13158 ) & (wr )  ;
assign n13160 =  ( n13159 ) ? ( n5298 ) : ( iram_75 ) ;
assign n13161 = wr_addr[7:7] ;
assign n13162 =  ( n13161 ) == ( bv_1_0_n53 )  ;
assign n13163 =  ( wr_addr ) == ( bv_8_75_n219 )  ;
assign n13164 =  ( n13162 ) & (n13163 )  ;
assign n13165 =  ( n13164 ) & (wr )  ;
assign n13166 =  ( n13165 ) ? ( n5325 ) : ( iram_75 ) ;
assign n13167 = wr_addr[7:7] ;
assign n13168 =  ( n13167 ) == ( bv_1_0_n53 )  ;
assign n13169 =  ( wr_addr ) == ( bv_8_76_n221 )  ;
assign n13170 =  ( n13168 ) & (n13169 )  ;
assign n13171 =  ( n13170 ) & (wr )  ;
assign n13172 =  ( n13171 ) ? ( n4782 ) : ( iram_76 ) ;
assign n13173 = wr_addr[7:7] ;
assign n13174 =  ( n13173 ) == ( bv_1_0_n53 )  ;
assign n13175 =  ( wr_addr ) == ( bv_8_76_n221 )  ;
assign n13176 =  ( n13174 ) & (n13175 )  ;
assign n13177 =  ( n13176 ) & (wr )  ;
assign n13178 =  ( n13177 ) ? ( n4841 ) : ( iram_76 ) ;
assign n13179 = wr_addr[7:7] ;
assign n13180 =  ( n13179 ) == ( bv_1_0_n53 )  ;
assign n13181 =  ( wr_addr ) == ( bv_8_76_n221 )  ;
assign n13182 =  ( n13180 ) & (n13181 )  ;
assign n13183 =  ( n13182 ) & (wr )  ;
assign n13184 =  ( n13183 ) ? ( n5449 ) : ( iram_76 ) ;
assign n13185 = wr_addr[7:7] ;
assign n13186 =  ( n13185 ) == ( bv_1_0_n53 )  ;
assign n13187 =  ( wr_addr ) == ( bv_8_76_n221 )  ;
assign n13188 =  ( n13186 ) & (n13187 )  ;
assign n13189 =  ( n13188 ) & (wr )  ;
assign n13190 =  ( n13189 ) ? ( n4906 ) : ( iram_76 ) ;
assign n13191 = wr_addr[7:7] ;
assign n13192 =  ( n13191 ) == ( bv_1_0_n53 )  ;
assign n13193 =  ( wr_addr ) == ( bv_8_76_n221 )  ;
assign n13194 =  ( n13192 ) & (n13193 )  ;
assign n13195 =  ( n13194 ) & (wr )  ;
assign n13196 =  ( n13195 ) ? ( n5485 ) : ( iram_76 ) ;
assign n13197 = wr_addr[7:7] ;
assign n13198 =  ( n13197 ) == ( bv_1_0_n53 )  ;
assign n13199 =  ( wr_addr ) == ( bv_8_76_n221 )  ;
assign n13200 =  ( n13198 ) & (n13199 )  ;
assign n13201 =  ( n13200 ) & (wr )  ;
assign n13202 =  ( n13201 ) ? ( n5512 ) : ( iram_76 ) ;
assign n13203 = wr_addr[7:7] ;
assign n13204 =  ( n13203 ) == ( bv_1_0_n53 )  ;
assign n13205 =  ( wr_addr ) == ( bv_8_76_n221 )  ;
assign n13206 =  ( n13204 ) & (n13205 )  ;
assign n13207 =  ( n13206 ) & (wr )  ;
assign n13208 =  ( n13207 ) ? ( bv_8_0_n69 ) : ( iram_76 ) ;
assign n13209 = wr_addr[7:7] ;
assign n13210 =  ( n13209 ) == ( bv_1_0_n53 )  ;
assign n13211 =  ( wr_addr ) == ( bv_8_76_n221 )  ;
assign n13212 =  ( n13210 ) & (n13211 )  ;
assign n13213 =  ( n13212 ) & (wr )  ;
assign n13214 =  ( n13213 ) ? ( n5071 ) : ( iram_76 ) ;
assign n13215 = wr_addr[7:7] ;
assign n13216 =  ( n13215 ) == ( bv_1_0_n53 )  ;
assign n13217 =  ( wr_addr ) == ( bv_8_76_n221 )  ;
assign n13218 =  ( n13216 ) & (n13217 )  ;
assign n13219 =  ( n13218 ) & (wr )  ;
assign n13220 =  ( n13219 ) ? ( n5096 ) : ( iram_76 ) ;
assign n13221 = wr_addr[7:7] ;
assign n13222 =  ( n13221 ) == ( bv_1_0_n53 )  ;
assign n13223 =  ( wr_addr ) == ( bv_8_76_n221 )  ;
assign n13224 =  ( n13222 ) & (n13223 )  ;
assign n13225 =  ( n13224 ) & (wr )  ;
assign n13226 =  ( n13225 ) ? ( n5123 ) : ( iram_76 ) ;
assign n13227 = wr_addr[7:7] ;
assign n13228 =  ( n13227 ) == ( bv_1_0_n53 )  ;
assign n13229 =  ( wr_addr ) == ( bv_8_76_n221 )  ;
assign n13230 =  ( n13228 ) & (n13229 )  ;
assign n13231 =  ( n13230 ) & (wr )  ;
assign n13232 =  ( n13231 ) ? ( n5165 ) : ( iram_76 ) ;
assign n13233 = wr_addr[7:7] ;
assign n13234 =  ( n13233 ) == ( bv_1_0_n53 )  ;
assign n13235 =  ( wr_addr ) == ( bv_8_76_n221 )  ;
assign n13236 =  ( n13234 ) & (n13235 )  ;
assign n13237 =  ( n13236 ) & (wr )  ;
assign n13238 =  ( n13237 ) ? ( n5204 ) : ( iram_76 ) ;
assign n13239 = wr_addr[7:7] ;
assign n13240 =  ( n13239 ) == ( bv_1_0_n53 )  ;
assign n13241 =  ( wr_addr ) == ( bv_8_76_n221 )  ;
assign n13242 =  ( n13240 ) & (n13241 )  ;
assign n13243 =  ( n13242 ) & (wr )  ;
assign n13244 =  ( n13243 ) ? ( n5262 ) : ( iram_76 ) ;
assign n13245 = wr_addr[7:7] ;
assign n13246 =  ( n13245 ) == ( bv_1_0_n53 )  ;
assign n13247 =  ( wr_addr ) == ( bv_8_76_n221 )  ;
assign n13248 =  ( n13246 ) & (n13247 )  ;
assign n13249 =  ( n13248 ) & (wr )  ;
assign n13250 =  ( n13249 ) ? ( n5298 ) : ( iram_76 ) ;
assign n13251 = wr_addr[7:7] ;
assign n13252 =  ( n13251 ) == ( bv_1_0_n53 )  ;
assign n13253 =  ( wr_addr ) == ( bv_8_76_n221 )  ;
assign n13254 =  ( n13252 ) & (n13253 )  ;
assign n13255 =  ( n13254 ) & (wr )  ;
assign n13256 =  ( n13255 ) ? ( n5325 ) : ( iram_76 ) ;
assign n13257 = wr_addr[7:7] ;
assign n13258 =  ( n13257 ) == ( bv_1_0_n53 )  ;
assign n13259 =  ( wr_addr ) == ( bv_8_77_n223 )  ;
assign n13260 =  ( n13258 ) & (n13259 )  ;
assign n13261 =  ( n13260 ) & (wr )  ;
assign n13262 =  ( n13261 ) ? ( n4782 ) : ( iram_77 ) ;
assign n13263 = wr_addr[7:7] ;
assign n13264 =  ( n13263 ) == ( bv_1_0_n53 )  ;
assign n13265 =  ( wr_addr ) == ( bv_8_77_n223 )  ;
assign n13266 =  ( n13264 ) & (n13265 )  ;
assign n13267 =  ( n13266 ) & (wr )  ;
assign n13268 =  ( n13267 ) ? ( n4841 ) : ( iram_77 ) ;
assign n13269 = wr_addr[7:7] ;
assign n13270 =  ( n13269 ) == ( bv_1_0_n53 )  ;
assign n13271 =  ( wr_addr ) == ( bv_8_77_n223 )  ;
assign n13272 =  ( n13270 ) & (n13271 )  ;
assign n13273 =  ( n13272 ) & (wr )  ;
assign n13274 =  ( n13273 ) ? ( n5449 ) : ( iram_77 ) ;
assign n13275 = wr_addr[7:7] ;
assign n13276 =  ( n13275 ) == ( bv_1_0_n53 )  ;
assign n13277 =  ( wr_addr ) == ( bv_8_77_n223 )  ;
assign n13278 =  ( n13276 ) & (n13277 )  ;
assign n13279 =  ( n13278 ) & (wr )  ;
assign n13280 =  ( n13279 ) ? ( n4906 ) : ( iram_77 ) ;
assign n13281 = wr_addr[7:7] ;
assign n13282 =  ( n13281 ) == ( bv_1_0_n53 )  ;
assign n13283 =  ( wr_addr ) == ( bv_8_77_n223 )  ;
assign n13284 =  ( n13282 ) & (n13283 )  ;
assign n13285 =  ( n13284 ) & (wr )  ;
assign n13286 =  ( n13285 ) ? ( n5485 ) : ( iram_77 ) ;
assign n13287 = wr_addr[7:7] ;
assign n13288 =  ( n13287 ) == ( bv_1_0_n53 )  ;
assign n13289 =  ( wr_addr ) == ( bv_8_77_n223 )  ;
assign n13290 =  ( n13288 ) & (n13289 )  ;
assign n13291 =  ( n13290 ) & (wr )  ;
assign n13292 =  ( n13291 ) ? ( n5512 ) : ( iram_77 ) ;
assign n13293 = wr_addr[7:7] ;
assign n13294 =  ( n13293 ) == ( bv_1_0_n53 )  ;
assign n13295 =  ( wr_addr ) == ( bv_8_77_n223 )  ;
assign n13296 =  ( n13294 ) & (n13295 )  ;
assign n13297 =  ( n13296 ) & (wr )  ;
assign n13298 =  ( n13297 ) ? ( bv_8_0_n69 ) : ( iram_77 ) ;
assign n13299 = wr_addr[7:7] ;
assign n13300 =  ( n13299 ) == ( bv_1_0_n53 )  ;
assign n13301 =  ( wr_addr ) == ( bv_8_77_n223 )  ;
assign n13302 =  ( n13300 ) & (n13301 )  ;
assign n13303 =  ( n13302 ) & (wr )  ;
assign n13304 =  ( n13303 ) ? ( n5071 ) : ( iram_77 ) ;
assign n13305 = wr_addr[7:7] ;
assign n13306 =  ( n13305 ) == ( bv_1_0_n53 )  ;
assign n13307 =  ( wr_addr ) == ( bv_8_77_n223 )  ;
assign n13308 =  ( n13306 ) & (n13307 )  ;
assign n13309 =  ( n13308 ) & (wr )  ;
assign n13310 =  ( n13309 ) ? ( n5096 ) : ( iram_77 ) ;
assign n13311 = wr_addr[7:7] ;
assign n13312 =  ( n13311 ) == ( bv_1_0_n53 )  ;
assign n13313 =  ( wr_addr ) == ( bv_8_77_n223 )  ;
assign n13314 =  ( n13312 ) & (n13313 )  ;
assign n13315 =  ( n13314 ) & (wr )  ;
assign n13316 =  ( n13315 ) ? ( n5123 ) : ( iram_77 ) ;
assign n13317 = wr_addr[7:7] ;
assign n13318 =  ( n13317 ) == ( bv_1_0_n53 )  ;
assign n13319 =  ( wr_addr ) == ( bv_8_77_n223 )  ;
assign n13320 =  ( n13318 ) & (n13319 )  ;
assign n13321 =  ( n13320 ) & (wr )  ;
assign n13322 =  ( n13321 ) ? ( n5165 ) : ( iram_77 ) ;
assign n13323 = wr_addr[7:7] ;
assign n13324 =  ( n13323 ) == ( bv_1_0_n53 )  ;
assign n13325 =  ( wr_addr ) == ( bv_8_77_n223 )  ;
assign n13326 =  ( n13324 ) & (n13325 )  ;
assign n13327 =  ( n13326 ) & (wr )  ;
assign n13328 =  ( n13327 ) ? ( n5204 ) : ( iram_77 ) ;
assign n13329 = wr_addr[7:7] ;
assign n13330 =  ( n13329 ) == ( bv_1_0_n53 )  ;
assign n13331 =  ( wr_addr ) == ( bv_8_77_n223 )  ;
assign n13332 =  ( n13330 ) & (n13331 )  ;
assign n13333 =  ( n13332 ) & (wr )  ;
assign n13334 =  ( n13333 ) ? ( n5262 ) : ( iram_77 ) ;
assign n13335 = wr_addr[7:7] ;
assign n13336 =  ( n13335 ) == ( bv_1_0_n53 )  ;
assign n13337 =  ( wr_addr ) == ( bv_8_77_n223 )  ;
assign n13338 =  ( n13336 ) & (n13337 )  ;
assign n13339 =  ( n13338 ) & (wr )  ;
assign n13340 =  ( n13339 ) ? ( n5298 ) : ( iram_77 ) ;
assign n13341 = wr_addr[7:7] ;
assign n13342 =  ( n13341 ) == ( bv_1_0_n53 )  ;
assign n13343 =  ( wr_addr ) == ( bv_8_77_n223 )  ;
assign n13344 =  ( n13342 ) & (n13343 )  ;
assign n13345 =  ( n13344 ) & (wr )  ;
assign n13346 =  ( n13345 ) ? ( n5325 ) : ( iram_77 ) ;
assign n13347 = wr_addr[7:7] ;
assign n13348 =  ( n13347 ) == ( bv_1_0_n53 )  ;
assign n13349 =  ( wr_addr ) == ( bv_8_78_n225 )  ;
assign n13350 =  ( n13348 ) & (n13349 )  ;
assign n13351 =  ( n13350 ) & (wr )  ;
assign n13352 =  ( n13351 ) ? ( n4782 ) : ( iram_78 ) ;
assign n13353 = wr_addr[7:7] ;
assign n13354 =  ( n13353 ) == ( bv_1_0_n53 )  ;
assign n13355 =  ( wr_addr ) == ( bv_8_78_n225 )  ;
assign n13356 =  ( n13354 ) & (n13355 )  ;
assign n13357 =  ( n13356 ) & (wr )  ;
assign n13358 =  ( n13357 ) ? ( n4841 ) : ( iram_78 ) ;
assign n13359 = wr_addr[7:7] ;
assign n13360 =  ( n13359 ) == ( bv_1_0_n53 )  ;
assign n13361 =  ( wr_addr ) == ( bv_8_78_n225 )  ;
assign n13362 =  ( n13360 ) & (n13361 )  ;
assign n13363 =  ( n13362 ) & (wr )  ;
assign n13364 =  ( n13363 ) ? ( n5449 ) : ( iram_78 ) ;
assign n13365 = wr_addr[7:7] ;
assign n13366 =  ( n13365 ) == ( bv_1_0_n53 )  ;
assign n13367 =  ( wr_addr ) == ( bv_8_78_n225 )  ;
assign n13368 =  ( n13366 ) & (n13367 )  ;
assign n13369 =  ( n13368 ) & (wr )  ;
assign n13370 =  ( n13369 ) ? ( n4906 ) : ( iram_78 ) ;
assign n13371 = wr_addr[7:7] ;
assign n13372 =  ( n13371 ) == ( bv_1_0_n53 )  ;
assign n13373 =  ( wr_addr ) == ( bv_8_78_n225 )  ;
assign n13374 =  ( n13372 ) & (n13373 )  ;
assign n13375 =  ( n13374 ) & (wr )  ;
assign n13376 =  ( n13375 ) ? ( n5485 ) : ( iram_78 ) ;
assign n13377 = wr_addr[7:7] ;
assign n13378 =  ( n13377 ) == ( bv_1_0_n53 )  ;
assign n13379 =  ( wr_addr ) == ( bv_8_78_n225 )  ;
assign n13380 =  ( n13378 ) & (n13379 )  ;
assign n13381 =  ( n13380 ) & (wr )  ;
assign n13382 =  ( n13381 ) ? ( n5512 ) : ( iram_78 ) ;
assign n13383 = wr_addr[7:7] ;
assign n13384 =  ( n13383 ) == ( bv_1_0_n53 )  ;
assign n13385 =  ( wr_addr ) == ( bv_8_78_n225 )  ;
assign n13386 =  ( n13384 ) & (n13385 )  ;
assign n13387 =  ( n13386 ) & (wr )  ;
assign n13388 =  ( n13387 ) ? ( bv_8_0_n69 ) : ( iram_78 ) ;
assign n13389 = wr_addr[7:7] ;
assign n13390 =  ( n13389 ) == ( bv_1_0_n53 )  ;
assign n13391 =  ( wr_addr ) == ( bv_8_78_n225 )  ;
assign n13392 =  ( n13390 ) & (n13391 )  ;
assign n13393 =  ( n13392 ) & (wr )  ;
assign n13394 =  ( n13393 ) ? ( n5071 ) : ( iram_78 ) ;
assign n13395 = wr_addr[7:7] ;
assign n13396 =  ( n13395 ) == ( bv_1_0_n53 )  ;
assign n13397 =  ( wr_addr ) == ( bv_8_78_n225 )  ;
assign n13398 =  ( n13396 ) & (n13397 )  ;
assign n13399 =  ( n13398 ) & (wr )  ;
assign n13400 =  ( n13399 ) ? ( n5096 ) : ( iram_78 ) ;
assign n13401 = wr_addr[7:7] ;
assign n13402 =  ( n13401 ) == ( bv_1_0_n53 )  ;
assign n13403 =  ( wr_addr ) == ( bv_8_78_n225 )  ;
assign n13404 =  ( n13402 ) & (n13403 )  ;
assign n13405 =  ( n13404 ) & (wr )  ;
assign n13406 =  ( n13405 ) ? ( n5123 ) : ( iram_78 ) ;
assign n13407 = wr_addr[7:7] ;
assign n13408 =  ( n13407 ) == ( bv_1_0_n53 )  ;
assign n13409 =  ( wr_addr ) == ( bv_8_78_n225 )  ;
assign n13410 =  ( n13408 ) & (n13409 )  ;
assign n13411 =  ( n13410 ) & (wr )  ;
assign n13412 =  ( n13411 ) ? ( n5165 ) : ( iram_78 ) ;
assign n13413 = wr_addr[7:7] ;
assign n13414 =  ( n13413 ) == ( bv_1_0_n53 )  ;
assign n13415 =  ( wr_addr ) == ( bv_8_78_n225 )  ;
assign n13416 =  ( n13414 ) & (n13415 )  ;
assign n13417 =  ( n13416 ) & (wr )  ;
assign n13418 =  ( n13417 ) ? ( n5204 ) : ( iram_78 ) ;
assign n13419 = wr_addr[7:7] ;
assign n13420 =  ( n13419 ) == ( bv_1_0_n53 )  ;
assign n13421 =  ( wr_addr ) == ( bv_8_78_n225 )  ;
assign n13422 =  ( n13420 ) & (n13421 )  ;
assign n13423 =  ( n13422 ) & (wr )  ;
assign n13424 =  ( n13423 ) ? ( n5262 ) : ( iram_78 ) ;
assign n13425 = wr_addr[7:7] ;
assign n13426 =  ( n13425 ) == ( bv_1_0_n53 )  ;
assign n13427 =  ( wr_addr ) == ( bv_8_78_n225 )  ;
assign n13428 =  ( n13426 ) & (n13427 )  ;
assign n13429 =  ( n13428 ) & (wr )  ;
assign n13430 =  ( n13429 ) ? ( n5298 ) : ( iram_78 ) ;
assign n13431 = wr_addr[7:7] ;
assign n13432 =  ( n13431 ) == ( bv_1_0_n53 )  ;
assign n13433 =  ( wr_addr ) == ( bv_8_78_n225 )  ;
assign n13434 =  ( n13432 ) & (n13433 )  ;
assign n13435 =  ( n13434 ) & (wr )  ;
assign n13436 =  ( n13435 ) ? ( n5325 ) : ( iram_78 ) ;
assign n13437 = wr_addr[7:7] ;
assign n13438 =  ( n13437 ) == ( bv_1_0_n53 )  ;
assign n13439 =  ( wr_addr ) == ( bv_8_79_n227 )  ;
assign n13440 =  ( n13438 ) & (n13439 )  ;
assign n13441 =  ( n13440 ) & (wr )  ;
assign n13442 =  ( n13441 ) ? ( n4782 ) : ( iram_79 ) ;
assign n13443 = wr_addr[7:7] ;
assign n13444 =  ( n13443 ) == ( bv_1_0_n53 )  ;
assign n13445 =  ( wr_addr ) == ( bv_8_79_n227 )  ;
assign n13446 =  ( n13444 ) & (n13445 )  ;
assign n13447 =  ( n13446 ) & (wr )  ;
assign n13448 =  ( n13447 ) ? ( n4841 ) : ( iram_79 ) ;
assign n13449 = wr_addr[7:7] ;
assign n13450 =  ( n13449 ) == ( bv_1_0_n53 )  ;
assign n13451 =  ( wr_addr ) == ( bv_8_79_n227 )  ;
assign n13452 =  ( n13450 ) & (n13451 )  ;
assign n13453 =  ( n13452 ) & (wr )  ;
assign n13454 =  ( n13453 ) ? ( n5449 ) : ( iram_79 ) ;
assign n13455 = wr_addr[7:7] ;
assign n13456 =  ( n13455 ) == ( bv_1_0_n53 )  ;
assign n13457 =  ( wr_addr ) == ( bv_8_79_n227 )  ;
assign n13458 =  ( n13456 ) & (n13457 )  ;
assign n13459 =  ( n13458 ) & (wr )  ;
assign n13460 =  ( n13459 ) ? ( n4906 ) : ( iram_79 ) ;
assign n13461 = wr_addr[7:7] ;
assign n13462 =  ( n13461 ) == ( bv_1_0_n53 )  ;
assign n13463 =  ( wr_addr ) == ( bv_8_79_n227 )  ;
assign n13464 =  ( n13462 ) & (n13463 )  ;
assign n13465 =  ( n13464 ) & (wr )  ;
assign n13466 =  ( n13465 ) ? ( n5485 ) : ( iram_79 ) ;
assign n13467 = wr_addr[7:7] ;
assign n13468 =  ( n13467 ) == ( bv_1_0_n53 )  ;
assign n13469 =  ( wr_addr ) == ( bv_8_79_n227 )  ;
assign n13470 =  ( n13468 ) & (n13469 )  ;
assign n13471 =  ( n13470 ) & (wr )  ;
assign n13472 =  ( n13471 ) ? ( n5512 ) : ( iram_79 ) ;
assign n13473 = wr_addr[7:7] ;
assign n13474 =  ( n13473 ) == ( bv_1_0_n53 )  ;
assign n13475 =  ( wr_addr ) == ( bv_8_79_n227 )  ;
assign n13476 =  ( n13474 ) & (n13475 )  ;
assign n13477 =  ( n13476 ) & (wr )  ;
assign n13478 =  ( n13477 ) ? ( bv_8_0_n69 ) : ( iram_79 ) ;
assign n13479 = wr_addr[7:7] ;
assign n13480 =  ( n13479 ) == ( bv_1_0_n53 )  ;
assign n13481 =  ( wr_addr ) == ( bv_8_79_n227 )  ;
assign n13482 =  ( n13480 ) & (n13481 )  ;
assign n13483 =  ( n13482 ) & (wr )  ;
assign n13484 =  ( n13483 ) ? ( n5071 ) : ( iram_79 ) ;
assign n13485 = wr_addr[7:7] ;
assign n13486 =  ( n13485 ) == ( bv_1_0_n53 )  ;
assign n13487 =  ( wr_addr ) == ( bv_8_79_n227 )  ;
assign n13488 =  ( n13486 ) & (n13487 )  ;
assign n13489 =  ( n13488 ) & (wr )  ;
assign n13490 =  ( n13489 ) ? ( n5096 ) : ( iram_79 ) ;
assign n13491 = wr_addr[7:7] ;
assign n13492 =  ( n13491 ) == ( bv_1_0_n53 )  ;
assign n13493 =  ( wr_addr ) == ( bv_8_79_n227 )  ;
assign n13494 =  ( n13492 ) & (n13493 )  ;
assign n13495 =  ( n13494 ) & (wr )  ;
assign n13496 =  ( n13495 ) ? ( n5123 ) : ( iram_79 ) ;
assign n13497 = wr_addr[7:7] ;
assign n13498 =  ( n13497 ) == ( bv_1_0_n53 )  ;
assign n13499 =  ( wr_addr ) == ( bv_8_79_n227 )  ;
assign n13500 =  ( n13498 ) & (n13499 )  ;
assign n13501 =  ( n13500 ) & (wr )  ;
assign n13502 =  ( n13501 ) ? ( n5165 ) : ( iram_79 ) ;
assign n13503 = wr_addr[7:7] ;
assign n13504 =  ( n13503 ) == ( bv_1_0_n53 )  ;
assign n13505 =  ( wr_addr ) == ( bv_8_79_n227 )  ;
assign n13506 =  ( n13504 ) & (n13505 )  ;
assign n13507 =  ( n13506 ) & (wr )  ;
assign n13508 =  ( n13507 ) ? ( n5204 ) : ( iram_79 ) ;
assign n13509 = wr_addr[7:7] ;
assign n13510 =  ( n13509 ) == ( bv_1_0_n53 )  ;
assign n13511 =  ( wr_addr ) == ( bv_8_79_n227 )  ;
assign n13512 =  ( n13510 ) & (n13511 )  ;
assign n13513 =  ( n13512 ) & (wr )  ;
assign n13514 =  ( n13513 ) ? ( n5262 ) : ( iram_79 ) ;
assign n13515 = wr_addr[7:7] ;
assign n13516 =  ( n13515 ) == ( bv_1_0_n53 )  ;
assign n13517 =  ( wr_addr ) == ( bv_8_79_n227 )  ;
assign n13518 =  ( n13516 ) & (n13517 )  ;
assign n13519 =  ( n13518 ) & (wr )  ;
assign n13520 =  ( n13519 ) ? ( n5298 ) : ( iram_79 ) ;
assign n13521 = wr_addr[7:7] ;
assign n13522 =  ( n13521 ) == ( bv_1_0_n53 )  ;
assign n13523 =  ( wr_addr ) == ( bv_8_79_n227 )  ;
assign n13524 =  ( n13522 ) & (n13523 )  ;
assign n13525 =  ( n13524 ) & (wr )  ;
assign n13526 =  ( n13525 ) ? ( n5325 ) : ( iram_79 ) ;
assign n13527 = wr_addr[7:7] ;
assign n13528 =  ( n13527 ) == ( bv_1_0_n53 )  ;
assign n13529 =  ( wr_addr ) == ( bv_8_80_n229 )  ;
assign n13530 =  ( n13528 ) & (n13529 )  ;
assign n13531 =  ( n13530 ) & (wr )  ;
assign n13532 =  ( n13531 ) ? ( n4782 ) : ( iram_80 ) ;
assign n13533 = wr_addr[7:7] ;
assign n13534 =  ( n13533 ) == ( bv_1_0_n53 )  ;
assign n13535 =  ( wr_addr ) == ( bv_8_80_n229 )  ;
assign n13536 =  ( n13534 ) & (n13535 )  ;
assign n13537 =  ( n13536 ) & (wr )  ;
assign n13538 =  ( n13537 ) ? ( n4841 ) : ( iram_80 ) ;
assign n13539 = wr_addr[7:7] ;
assign n13540 =  ( n13539 ) == ( bv_1_0_n53 )  ;
assign n13541 =  ( wr_addr ) == ( bv_8_80_n229 )  ;
assign n13542 =  ( n13540 ) & (n13541 )  ;
assign n13543 =  ( n13542 ) & (wr )  ;
assign n13544 =  ( n13543 ) ? ( n5449 ) : ( iram_80 ) ;
assign n13545 = wr_addr[7:7] ;
assign n13546 =  ( n13545 ) == ( bv_1_0_n53 )  ;
assign n13547 =  ( wr_addr ) == ( bv_8_80_n229 )  ;
assign n13548 =  ( n13546 ) & (n13547 )  ;
assign n13549 =  ( n13548 ) & (wr )  ;
assign n13550 =  ( n13549 ) ? ( n4906 ) : ( iram_80 ) ;
assign n13551 = wr_addr[7:7] ;
assign n13552 =  ( n13551 ) == ( bv_1_0_n53 )  ;
assign n13553 =  ( wr_addr ) == ( bv_8_80_n229 )  ;
assign n13554 =  ( n13552 ) & (n13553 )  ;
assign n13555 =  ( n13554 ) & (wr )  ;
assign n13556 =  ( n13555 ) ? ( n5485 ) : ( iram_80 ) ;
assign n13557 = wr_addr[7:7] ;
assign n13558 =  ( n13557 ) == ( bv_1_0_n53 )  ;
assign n13559 =  ( wr_addr ) == ( bv_8_80_n229 )  ;
assign n13560 =  ( n13558 ) & (n13559 )  ;
assign n13561 =  ( n13560 ) & (wr )  ;
assign n13562 =  ( n13561 ) ? ( n5512 ) : ( iram_80 ) ;
assign n13563 = wr_addr[7:7] ;
assign n13564 =  ( n13563 ) == ( bv_1_0_n53 )  ;
assign n13565 =  ( wr_addr ) == ( bv_8_80_n229 )  ;
assign n13566 =  ( n13564 ) & (n13565 )  ;
assign n13567 =  ( n13566 ) & (wr )  ;
assign n13568 =  ( n13567 ) ? ( bv_8_0_n69 ) : ( iram_80 ) ;
assign n13569 = wr_addr[7:7] ;
assign n13570 =  ( n13569 ) == ( bv_1_0_n53 )  ;
assign n13571 =  ( wr_addr ) == ( bv_8_80_n229 )  ;
assign n13572 =  ( n13570 ) & (n13571 )  ;
assign n13573 =  ( n13572 ) & (wr )  ;
assign n13574 =  ( n13573 ) ? ( n5071 ) : ( iram_80 ) ;
assign n13575 = wr_addr[7:7] ;
assign n13576 =  ( n13575 ) == ( bv_1_0_n53 )  ;
assign n13577 =  ( wr_addr ) == ( bv_8_80_n229 )  ;
assign n13578 =  ( n13576 ) & (n13577 )  ;
assign n13579 =  ( n13578 ) & (wr )  ;
assign n13580 =  ( n13579 ) ? ( n5096 ) : ( iram_80 ) ;
assign n13581 = wr_addr[7:7] ;
assign n13582 =  ( n13581 ) == ( bv_1_0_n53 )  ;
assign n13583 =  ( wr_addr ) == ( bv_8_80_n229 )  ;
assign n13584 =  ( n13582 ) & (n13583 )  ;
assign n13585 =  ( n13584 ) & (wr )  ;
assign n13586 =  ( n13585 ) ? ( n5123 ) : ( iram_80 ) ;
assign n13587 = wr_addr[7:7] ;
assign n13588 =  ( n13587 ) == ( bv_1_0_n53 )  ;
assign n13589 =  ( wr_addr ) == ( bv_8_80_n229 )  ;
assign n13590 =  ( n13588 ) & (n13589 )  ;
assign n13591 =  ( n13590 ) & (wr )  ;
assign n13592 =  ( n13591 ) ? ( n5165 ) : ( iram_80 ) ;
assign n13593 = wr_addr[7:7] ;
assign n13594 =  ( n13593 ) == ( bv_1_0_n53 )  ;
assign n13595 =  ( wr_addr ) == ( bv_8_80_n229 )  ;
assign n13596 =  ( n13594 ) & (n13595 )  ;
assign n13597 =  ( n13596 ) & (wr )  ;
assign n13598 =  ( n13597 ) ? ( n5204 ) : ( iram_80 ) ;
assign n13599 = wr_addr[7:7] ;
assign n13600 =  ( n13599 ) == ( bv_1_0_n53 )  ;
assign n13601 =  ( wr_addr ) == ( bv_8_80_n229 )  ;
assign n13602 =  ( n13600 ) & (n13601 )  ;
assign n13603 =  ( n13602 ) & (wr )  ;
assign n13604 =  ( n13603 ) ? ( n5262 ) : ( iram_80 ) ;
assign n13605 = wr_addr[7:7] ;
assign n13606 =  ( n13605 ) == ( bv_1_0_n53 )  ;
assign n13607 =  ( wr_addr ) == ( bv_8_80_n229 )  ;
assign n13608 =  ( n13606 ) & (n13607 )  ;
assign n13609 =  ( n13608 ) & (wr )  ;
assign n13610 =  ( n13609 ) ? ( n5298 ) : ( iram_80 ) ;
assign n13611 = wr_addr[7:7] ;
assign n13612 =  ( n13611 ) == ( bv_1_0_n53 )  ;
assign n13613 =  ( wr_addr ) == ( bv_8_80_n229 )  ;
assign n13614 =  ( n13612 ) & (n13613 )  ;
assign n13615 =  ( n13614 ) & (wr )  ;
assign n13616 =  ( n13615 ) ? ( n5325 ) : ( iram_80 ) ;
assign n13617 = wr_addr[7:7] ;
assign n13618 =  ( n13617 ) == ( bv_1_0_n53 )  ;
assign n13619 =  ( wr_addr ) == ( bv_8_81_n231 )  ;
assign n13620 =  ( n13618 ) & (n13619 )  ;
assign n13621 =  ( n13620 ) & (wr )  ;
assign n13622 =  ( n13621 ) ? ( n4782 ) : ( iram_81 ) ;
assign n13623 = wr_addr[7:7] ;
assign n13624 =  ( n13623 ) == ( bv_1_0_n53 )  ;
assign n13625 =  ( wr_addr ) == ( bv_8_81_n231 )  ;
assign n13626 =  ( n13624 ) & (n13625 )  ;
assign n13627 =  ( n13626 ) & (wr )  ;
assign n13628 =  ( n13627 ) ? ( n4841 ) : ( iram_81 ) ;
assign n13629 = wr_addr[7:7] ;
assign n13630 =  ( n13629 ) == ( bv_1_0_n53 )  ;
assign n13631 =  ( wr_addr ) == ( bv_8_81_n231 )  ;
assign n13632 =  ( n13630 ) & (n13631 )  ;
assign n13633 =  ( n13632 ) & (wr )  ;
assign n13634 =  ( n13633 ) ? ( n5449 ) : ( iram_81 ) ;
assign n13635 = wr_addr[7:7] ;
assign n13636 =  ( n13635 ) == ( bv_1_0_n53 )  ;
assign n13637 =  ( wr_addr ) == ( bv_8_81_n231 )  ;
assign n13638 =  ( n13636 ) & (n13637 )  ;
assign n13639 =  ( n13638 ) & (wr )  ;
assign n13640 =  ( n13639 ) ? ( n4906 ) : ( iram_81 ) ;
assign n13641 = wr_addr[7:7] ;
assign n13642 =  ( n13641 ) == ( bv_1_0_n53 )  ;
assign n13643 =  ( wr_addr ) == ( bv_8_81_n231 )  ;
assign n13644 =  ( n13642 ) & (n13643 )  ;
assign n13645 =  ( n13644 ) & (wr )  ;
assign n13646 =  ( n13645 ) ? ( n5485 ) : ( iram_81 ) ;
assign n13647 = wr_addr[7:7] ;
assign n13648 =  ( n13647 ) == ( bv_1_0_n53 )  ;
assign n13649 =  ( wr_addr ) == ( bv_8_81_n231 )  ;
assign n13650 =  ( n13648 ) & (n13649 )  ;
assign n13651 =  ( n13650 ) & (wr )  ;
assign n13652 =  ( n13651 ) ? ( n5512 ) : ( iram_81 ) ;
assign n13653 = wr_addr[7:7] ;
assign n13654 =  ( n13653 ) == ( bv_1_0_n53 )  ;
assign n13655 =  ( wr_addr ) == ( bv_8_81_n231 )  ;
assign n13656 =  ( n13654 ) & (n13655 )  ;
assign n13657 =  ( n13656 ) & (wr )  ;
assign n13658 =  ( n13657 ) ? ( bv_8_0_n69 ) : ( iram_81 ) ;
assign n13659 = wr_addr[7:7] ;
assign n13660 =  ( n13659 ) == ( bv_1_0_n53 )  ;
assign n13661 =  ( wr_addr ) == ( bv_8_81_n231 )  ;
assign n13662 =  ( n13660 ) & (n13661 )  ;
assign n13663 =  ( n13662 ) & (wr )  ;
assign n13664 =  ( n13663 ) ? ( n5071 ) : ( iram_81 ) ;
assign n13665 = wr_addr[7:7] ;
assign n13666 =  ( n13665 ) == ( bv_1_0_n53 )  ;
assign n13667 =  ( wr_addr ) == ( bv_8_81_n231 )  ;
assign n13668 =  ( n13666 ) & (n13667 )  ;
assign n13669 =  ( n13668 ) & (wr )  ;
assign n13670 =  ( n13669 ) ? ( n5096 ) : ( iram_81 ) ;
assign n13671 = wr_addr[7:7] ;
assign n13672 =  ( n13671 ) == ( bv_1_0_n53 )  ;
assign n13673 =  ( wr_addr ) == ( bv_8_81_n231 )  ;
assign n13674 =  ( n13672 ) & (n13673 )  ;
assign n13675 =  ( n13674 ) & (wr )  ;
assign n13676 =  ( n13675 ) ? ( n5123 ) : ( iram_81 ) ;
assign n13677 = wr_addr[7:7] ;
assign n13678 =  ( n13677 ) == ( bv_1_0_n53 )  ;
assign n13679 =  ( wr_addr ) == ( bv_8_81_n231 )  ;
assign n13680 =  ( n13678 ) & (n13679 )  ;
assign n13681 =  ( n13680 ) & (wr )  ;
assign n13682 =  ( n13681 ) ? ( n5165 ) : ( iram_81 ) ;
assign n13683 = wr_addr[7:7] ;
assign n13684 =  ( n13683 ) == ( bv_1_0_n53 )  ;
assign n13685 =  ( wr_addr ) == ( bv_8_81_n231 )  ;
assign n13686 =  ( n13684 ) & (n13685 )  ;
assign n13687 =  ( n13686 ) & (wr )  ;
assign n13688 =  ( n13687 ) ? ( n5204 ) : ( iram_81 ) ;
assign n13689 = wr_addr[7:7] ;
assign n13690 =  ( n13689 ) == ( bv_1_0_n53 )  ;
assign n13691 =  ( wr_addr ) == ( bv_8_81_n231 )  ;
assign n13692 =  ( n13690 ) & (n13691 )  ;
assign n13693 =  ( n13692 ) & (wr )  ;
assign n13694 =  ( n13693 ) ? ( n5262 ) : ( iram_81 ) ;
assign n13695 = wr_addr[7:7] ;
assign n13696 =  ( n13695 ) == ( bv_1_0_n53 )  ;
assign n13697 =  ( wr_addr ) == ( bv_8_81_n231 )  ;
assign n13698 =  ( n13696 ) & (n13697 )  ;
assign n13699 =  ( n13698 ) & (wr )  ;
assign n13700 =  ( n13699 ) ? ( n5298 ) : ( iram_81 ) ;
assign n13701 = wr_addr[7:7] ;
assign n13702 =  ( n13701 ) == ( bv_1_0_n53 )  ;
assign n13703 =  ( wr_addr ) == ( bv_8_81_n231 )  ;
assign n13704 =  ( n13702 ) & (n13703 )  ;
assign n13705 =  ( n13704 ) & (wr )  ;
assign n13706 =  ( n13705 ) ? ( n5325 ) : ( iram_81 ) ;
assign n13707 = wr_addr[7:7] ;
assign n13708 =  ( n13707 ) == ( bv_1_0_n53 )  ;
assign n13709 =  ( wr_addr ) == ( bv_8_82_n233 )  ;
assign n13710 =  ( n13708 ) & (n13709 )  ;
assign n13711 =  ( n13710 ) & (wr )  ;
assign n13712 =  ( n13711 ) ? ( n4782 ) : ( iram_82 ) ;
assign n13713 = wr_addr[7:7] ;
assign n13714 =  ( n13713 ) == ( bv_1_0_n53 )  ;
assign n13715 =  ( wr_addr ) == ( bv_8_82_n233 )  ;
assign n13716 =  ( n13714 ) & (n13715 )  ;
assign n13717 =  ( n13716 ) & (wr )  ;
assign n13718 =  ( n13717 ) ? ( n4841 ) : ( iram_82 ) ;
assign n13719 = wr_addr[7:7] ;
assign n13720 =  ( n13719 ) == ( bv_1_0_n53 )  ;
assign n13721 =  ( wr_addr ) == ( bv_8_82_n233 )  ;
assign n13722 =  ( n13720 ) & (n13721 )  ;
assign n13723 =  ( n13722 ) & (wr )  ;
assign n13724 =  ( n13723 ) ? ( n5449 ) : ( iram_82 ) ;
assign n13725 = wr_addr[7:7] ;
assign n13726 =  ( n13725 ) == ( bv_1_0_n53 )  ;
assign n13727 =  ( wr_addr ) == ( bv_8_82_n233 )  ;
assign n13728 =  ( n13726 ) & (n13727 )  ;
assign n13729 =  ( n13728 ) & (wr )  ;
assign n13730 =  ( n13729 ) ? ( n4906 ) : ( iram_82 ) ;
assign n13731 = wr_addr[7:7] ;
assign n13732 =  ( n13731 ) == ( bv_1_0_n53 )  ;
assign n13733 =  ( wr_addr ) == ( bv_8_82_n233 )  ;
assign n13734 =  ( n13732 ) & (n13733 )  ;
assign n13735 =  ( n13734 ) & (wr )  ;
assign n13736 =  ( n13735 ) ? ( n5485 ) : ( iram_82 ) ;
assign n13737 = wr_addr[7:7] ;
assign n13738 =  ( n13737 ) == ( bv_1_0_n53 )  ;
assign n13739 =  ( wr_addr ) == ( bv_8_82_n233 )  ;
assign n13740 =  ( n13738 ) & (n13739 )  ;
assign n13741 =  ( n13740 ) & (wr )  ;
assign n13742 =  ( n13741 ) ? ( n5512 ) : ( iram_82 ) ;
assign n13743 = wr_addr[7:7] ;
assign n13744 =  ( n13743 ) == ( bv_1_0_n53 )  ;
assign n13745 =  ( wr_addr ) == ( bv_8_82_n233 )  ;
assign n13746 =  ( n13744 ) & (n13745 )  ;
assign n13747 =  ( n13746 ) & (wr )  ;
assign n13748 =  ( n13747 ) ? ( bv_8_0_n69 ) : ( iram_82 ) ;
assign n13749 = wr_addr[7:7] ;
assign n13750 =  ( n13749 ) == ( bv_1_0_n53 )  ;
assign n13751 =  ( wr_addr ) == ( bv_8_82_n233 )  ;
assign n13752 =  ( n13750 ) & (n13751 )  ;
assign n13753 =  ( n13752 ) & (wr )  ;
assign n13754 =  ( n13753 ) ? ( n5071 ) : ( iram_82 ) ;
assign n13755 = wr_addr[7:7] ;
assign n13756 =  ( n13755 ) == ( bv_1_0_n53 )  ;
assign n13757 =  ( wr_addr ) == ( bv_8_82_n233 )  ;
assign n13758 =  ( n13756 ) & (n13757 )  ;
assign n13759 =  ( n13758 ) & (wr )  ;
assign n13760 =  ( n13759 ) ? ( n5096 ) : ( iram_82 ) ;
assign n13761 = wr_addr[7:7] ;
assign n13762 =  ( n13761 ) == ( bv_1_0_n53 )  ;
assign n13763 =  ( wr_addr ) == ( bv_8_82_n233 )  ;
assign n13764 =  ( n13762 ) & (n13763 )  ;
assign n13765 =  ( n13764 ) & (wr )  ;
assign n13766 =  ( n13765 ) ? ( n5123 ) : ( iram_82 ) ;
assign n13767 = wr_addr[7:7] ;
assign n13768 =  ( n13767 ) == ( bv_1_0_n53 )  ;
assign n13769 =  ( wr_addr ) == ( bv_8_82_n233 )  ;
assign n13770 =  ( n13768 ) & (n13769 )  ;
assign n13771 =  ( n13770 ) & (wr )  ;
assign n13772 =  ( n13771 ) ? ( n5165 ) : ( iram_82 ) ;
assign n13773 = wr_addr[7:7] ;
assign n13774 =  ( n13773 ) == ( bv_1_0_n53 )  ;
assign n13775 =  ( wr_addr ) == ( bv_8_82_n233 )  ;
assign n13776 =  ( n13774 ) & (n13775 )  ;
assign n13777 =  ( n13776 ) & (wr )  ;
assign n13778 =  ( n13777 ) ? ( n5204 ) : ( iram_82 ) ;
assign n13779 = wr_addr[7:7] ;
assign n13780 =  ( n13779 ) == ( bv_1_0_n53 )  ;
assign n13781 =  ( wr_addr ) == ( bv_8_82_n233 )  ;
assign n13782 =  ( n13780 ) & (n13781 )  ;
assign n13783 =  ( n13782 ) & (wr )  ;
assign n13784 =  ( n13783 ) ? ( n5262 ) : ( iram_82 ) ;
assign n13785 = wr_addr[7:7] ;
assign n13786 =  ( n13785 ) == ( bv_1_0_n53 )  ;
assign n13787 =  ( wr_addr ) == ( bv_8_82_n233 )  ;
assign n13788 =  ( n13786 ) & (n13787 )  ;
assign n13789 =  ( n13788 ) & (wr )  ;
assign n13790 =  ( n13789 ) ? ( n5298 ) : ( iram_82 ) ;
assign n13791 = wr_addr[7:7] ;
assign n13792 =  ( n13791 ) == ( bv_1_0_n53 )  ;
assign n13793 =  ( wr_addr ) == ( bv_8_82_n233 )  ;
assign n13794 =  ( n13792 ) & (n13793 )  ;
assign n13795 =  ( n13794 ) & (wr )  ;
assign n13796 =  ( n13795 ) ? ( n5325 ) : ( iram_82 ) ;
assign n13797 = wr_addr[7:7] ;
assign n13798 =  ( n13797 ) == ( bv_1_0_n53 )  ;
assign n13799 =  ( wr_addr ) == ( bv_8_83_n235 )  ;
assign n13800 =  ( n13798 ) & (n13799 )  ;
assign n13801 =  ( n13800 ) & (wr )  ;
assign n13802 =  ( n13801 ) ? ( n4782 ) : ( iram_83 ) ;
assign n13803 = wr_addr[7:7] ;
assign n13804 =  ( n13803 ) == ( bv_1_0_n53 )  ;
assign n13805 =  ( wr_addr ) == ( bv_8_83_n235 )  ;
assign n13806 =  ( n13804 ) & (n13805 )  ;
assign n13807 =  ( n13806 ) & (wr )  ;
assign n13808 =  ( n13807 ) ? ( n4841 ) : ( iram_83 ) ;
assign n13809 = wr_addr[7:7] ;
assign n13810 =  ( n13809 ) == ( bv_1_0_n53 )  ;
assign n13811 =  ( wr_addr ) == ( bv_8_83_n235 )  ;
assign n13812 =  ( n13810 ) & (n13811 )  ;
assign n13813 =  ( n13812 ) & (wr )  ;
assign n13814 =  ( n13813 ) ? ( n5449 ) : ( iram_83 ) ;
assign n13815 = wr_addr[7:7] ;
assign n13816 =  ( n13815 ) == ( bv_1_0_n53 )  ;
assign n13817 =  ( wr_addr ) == ( bv_8_83_n235 )  ;
assign n13818 =  ( n13816 ) & (n13817 )  ;
assign n13819 =  ( n13818 ) & (wr )  ;
assign n13820 =  ( n13819 ) ? ( n4906 ) : ( iram_83 ) ;
assign n13821 = wr_addr[7:7] ;
assign n13822 =  ( n13821 ) == ( bv_1_0_n53 )  ;
assign n13823 =  ( wr_addr ) == ( bv_8_83_n235 )  ;
assign n13824 =  ( n13822 ) & (n13823 )  ;
assign n13825 =  ( n13824 ) & (wr )  ;
assign n13826 =  ( n13825 ) ? ( n5485 ) : ( iram_83 ) ;
assign n13827 = wr_addr[7:7] ;
assign n13828 =  ( n13827 ) == ( bv_1_0_n53 )  ;
assign n13829 =  ( wr_addr ) == ( bv_8_83_n235 )  ;
assign n13830 =  ( n13828 ) & (n13829 )  ;
assign n13831 =  ( n13830 ) & (wr )  ;
assign n13832 =  ( n13831 ) ? ( n5512 ) : ( iram_83 ) ;
assign n13833 = wr_addr[7:7] ;
assign n13834 =  ( n13833 ) == ( bv_1_0_n53 )  ;
assign n13835 =  ( wr_addr ) == ( bv_8_83_n235 )  ;
assign n13836 =  ( n13834 ) & (n13835 )  ;
assign n13837 =  ( n13836 ) & (wr )  ;
assign n13838 =  ( n13837 ) ? ( bv_8_0_n69 ) : ( iram_83 ) ;
assign n13839 = wr_addr[7:7] ;
assign n13840 =  ( n13839 ) == ( bv_1_0_n53 )  ;
assign n13841 =  ( wr_addr ) == ( bv_8_83_n235 )  ;
assign n13842 =  ( n13840 ) & (n13841 )  ;
assign n13843 =  ( n13842 ) & (wr )  ;
assign n13844 =  ( n13843 ) ? ( n5071 ) : ( iram_83 ) ;
assign n13845 = wr_addr[7:7] ;
assign n13846 =  ( n13845 ) == ( bv_1_0_n53 )  ;
assign n13847 =  ( wr_addr ) == ( bv_8_83_n235 )  ;
assign n13848 =  ( n13846 ) & (n13847 )  ;
assign n13849 =  ( n13848 ) & (wr )  ;
assign n13850 =  ( n13849 ) ? ( n5096 ) : ( iram_83 ) ;
assign n13851 = wr_addr[7:7] ;
assign n13852 =  ( n13851 ) == ( bv_1_0_n53 )  ;
assign n13853 =  ( wr_addr ) == ( bv_8_83_n235 )  ;
assign n13854 =  ( n13852 ) & (n13853 )  ;
assign n13855 =  ( n13854 ) & (wr )  ;
assign n13856 =  ( n13855 ) ? ( n5123 ) : ( iram_83 ) ;
assign n13857 = wr_addr[7:7] ;
assign n13858 =  ( n13857 ) == ( bv_1_0_n53 )  ;
assign n13859 =  ( wr_addr ) == ( bv_8_83_n235 )  ;
assign n13860 =  ( n13858 ) & (n13859 )  ;
assign n13861 =  ( n13860 ) & (wr )  ;
assign n13862 =  ( n13861 ) ? ( n5165 ) : ( iram_83 ) ;
assign n13863 = wr_addr[7:7] ;
assign n13864 =  ( n13863 ) == ( bv_1_0_n53 )  ;
assign n13865 =  ( wr_addr ) == ( bv_8_83_n235 )  ;
assign n13866 =  ( n13864 ) & (n13865 )  ;
assign n13867 =  ( n13866 ) & (wr )  ;
assign n13868 =  ( n13867 ) ? ( n5204 ) : ( iram_83 ) ;
assign n13869 = wr_addr[7:7] ;
assign n13870 =  ( n13869 ) == ( bv_1_0_n53 )  ;
assign n13871 =  ( wr_addr ) == ( bv_8_83_n235 )  ;
assign n13872 =  ( n13870 ) & (n13871 )  ;
assign n13873 =  ( n13872 ) & (wr )  ;
assign n13874 =  ( n13873 ) ? ( n5262 ) : ( iram_83 ) ;
assign n13875 = wr_addr[7:7] ;
assign n13876 =  ( n13875 ) == ( bv_1_0_n53 )  ;
assign n13877 =  ( wr_addr ) == ( bv_8_83_n235 )  ;
assign n13878 =  ( n13876 ) & (n13877 )  ;
assign n13879 =  ( n13878 ) & (wr )  ;
assign n13880 =  ( n13879 ) ? ( n5298 ) : ( iram_83 ) ;
assign n13881 = wr_addr[7:7] ;
assign n13882 =  ( n13881 ) == ( bv_1_0_n53 )  ;
assign n13883 =  ( wr_addr ) == ( bv_8_83_n235 )  ;
assign n13884 =  ( n13882 ) & (n13883 )  ;
assign n13885 =  ( n13884 ) & (wr )  ;
assign n13886 =  ( n13885 ) ? ( n5325 ) : ( iram_83 ) ;
assign n13887 = wr_addr[7:7] ;
assign n13888 =  ( n13887 ) == ( bv_1_0_n53 )  ;
assign n13889 =  ( wr_addr ) == ( bv_8_84_n237 )  ;
assign n13890 =  ( n13888 ) & (n13889 )  ;
assign n13891 =  ( n13890 ) & (wr )  ;
assign n13892 =  ( n13891 ) ? ( n4782 ) : ( iram_84 ) ;
assign n13893 = wr_addr[7:7] ;
assign n13894 =  ( n13893 ) == ( bv_1_0_n53 )  ;
assign n13895 =  ( wr_addr ) == ( bv_8_84_n237 )  ;
assign n13896 =  ( n13894 ) & (n13895 )  ;
assign n13897 =  ( n13896 ) & (wr )  ;
assign n13898 =  ( n13897 ) ? ( n4841 ) : ( iram_84 ) ;
assign n13899 = wr_addr[7:7] ;
assign n13900 =  ( n13899 ) == ( bv_1_0_n53 )  ;
assign n13901 =  ( wr_addr ) == ( bv_8_84_n237 )  ;
assign n13902 =  ( n13900 ) & (n13901 )  ;
assign n13903 =  ( n13902 ) & (wr )  ;
assign n13904 =  ( n13903 ) ? ( n5449 ) : ( iram_84 ) ;
assign n13905 = wr_addr[7:7] ;
assign n13906 =  ( n13905 ) == ( bv_1_0_n53 )  ;
assign n13907 =  ( wr_addr ) == ( bv_8_84_n237 )  ;
assign n13908 =  ( n13906 ) & (n13907 )  ;
assign n13909 =  ( n13908 ) & (wr )  ;
assign n13910 =  ( n13909 ) ? ( n4906 ) : ( iram_84 ) ;
assign n13911 = wr_addr[7:7] ;
assign n13912 =  ( n13911 ) == ( bv_1_0_n53 )  ;
assign n13913 =  ( wr_addr ) == ( bv_8_84_n237 )  ;
assign n13914 =  ( n13912 ) & (n13913 )  ;
assign n13915 =  ( n13914 ) & (wr )  ;
assign n13916 =  ( n13915 ) ? ( n5485 ) : ( iram_84 ) ;
assign n13917 = wr_addr[7:7] ;
assign n13918 =  ( n13917 ) == ( bv_1_0_n53 )  ;
assign n13919 =  ( wr_addr ) == ( bv_8_84_n237 )  ;
assign n13920 =  ( n13918 ) & (n13919 )  ;
assign n13921 =  ( n13920 ) & (wr )  ;
assign n13922 =  ( n13921 ) ? ( n5512 ) : ( iram_84 ) ;
assign n13923 = wr_addr[7:7] ;
assign n13924 =  ( n13923 ) == ( bv_1_0_n53 )  ;
assign n13925 =  ( wr_addr ) == ( bv_8_84_n237 )  ;
assign n13926 =  ( n13924 ) & (n13925 )  ;
assign n13927 =  ( n13926 ) & (wr )  ;
assign n13928 =  ( n13927 ) ? ( bv_8_0_n69 ) : ( iram_84 ) ;
assign n13929 = wr_addr[7:7] ;
assign n13930 =  ( n13929 ) == ( bv_1_0_n53 )  ;
assign n13931 =  ( wr_addr ) == ( bv_8_84_n237 )  ;
assign n13932 =  ( n13930 ) & (n13931 )  ;
assign n13933 =  ( n13932 ) & (wr )  ;
assign n13934 =  ( n13933 ) ? ( n5071 ) : ( iram_84 ) ;
assign n13935 = wr_addr[7:7] ;
assign n13936 =  ( n13935 ) == ( bv_1_0_n53 )  ;
assign n13937 =  ( wr_addr ) == ( bv_8_84_n237 )  ;
assign n13938 =  ( n13936 ) & (n13937 )  ;
assign n13939 =  ( n13938 ) & (wr )  ;
assign n13940 =  ( n13939 ) ? ( n5096 ) : ( iram_84 ) ;
assign n13941 = wr_addr[7:7] ;
assign n13942 =  ( n13941 ) == ( bv_1_0_n53 )  ;
assign n13943 =  ( wr_addr ) == ( bv_8_84_n237 )  ;
assign n13944 =  ( n13942 ) & (n13943 )  ;
assign n13945 =  ( n13944 ) & (wr )  ;
assign n13946 =  ( n13945 ) ? ( n5123 ) : ( iram_84 ) ;
assign n13947 = wr_addr[7:7] ;
assign n13948 =  ( n13947 ) == ( bv_1_0_n53 )  ;
assign n13949 =  ( wr_addr ) == ( bv_8_84_n237 )  ;
assign n13950 =  ( n13948 ) & (n13949 )  ;
assign n13951 =  ( n13950 ) & (wr )  ;
assign n13952 =  ( n13951 ) ? ( n5165 ) : ( iram_84 ) ;
assign n13953 = wr_addr[7:7] ;
assign n13954 =  ( n13953 ) == ( bv_1_0_n53 )  ;
assign n13955 =  ( wr_addr ) == ( bv_8_84_n237 )  ;
assign n13956 =  ( n13954 ) & (n13955 )  ;
assign n13957 =  ( n13956 ) & (wr )  ;
assign n13958 =  ( n13957 ) ? ( n5204 ) : ( iram_84 ) ;
assign n13959 = wr_addr[7:7] ;
assign n13960 =  ( n13959 ) == ( bv_1_0_n53 )  ;
assign n13961 =  ( wr_addr ) == ( bv_8_84_n237 )  ;
assign n13962 =  ( n13960 ) & (n13961 )  ;
assign n13963 =  ( n13962 ) & (wr )  ;
assign n13964 =  ( n13963 ) ? ( n5262 ) : ( iram_84 ) ;
assign n13965 = wr_addr[7:7] ;
assign n13966 =  ( n13965 ) == ( bv_1_0_n53 )  ;
assign n13967 =  ( wr_addr ) == ( bv_8_84_n237 )  ;
assign n13968 =  ( n13966 ) & (n13967 )  ;
assign n13969 =  ( n13968 ) & (wr )  ;
assign n13970 =  ( n13969 ) ? ( n5298 ) : ( iram_84 ) ;
assign n13971 = wr_addr[7:7] ;
assign n13972 =  ( n13971 ) == ( bv_1_0_n53 )  ;
assign n13973 =  ( wr_addr ) == ( bv_8_84_n237 )  ;
assign n13974 =  ( n13972 ) & (n13973 )  ;
assign n13975 =  ( n13974 ) & (wr )  ;
assign n13976 =  ( n13975 ) ? ( n5325 ) : ( iram_84 ) ;
assign n13977 = wr_addr[7:7] ;
assign n13978 =  ( n13977 ) == ( bv_1_0_n53 )  ;
assign n13979 =  ( wr_addr ) == ( bv_8_85_n239 )  ;
assign n13980 =  ( n13978 ) & (n13979 )  ;
assign n13981 =  ( n13980 ) & (wr )  ;
assign n13982 =  ( n13981 ) ? ( n4782 ) : ( iram_85 ) ;
assign n13983 = wr_addr[7:7] ;
assign n13984 =  ( n13983 ) == ( bv_1_0_n53 )  ;
assign n13985 =  ( wr_addr ) == ( bv_8_85_n239 )  ;
assign n13986 =  ( n13984 ) & (n13985 )  ;
assign n13987 =  ( n13986 ) & (wr )  ;
assign n13988 =  ( n13987 ) ? ( n4841 ) : ( iram_85 ) ;
assign n13989 = wr_addr[7:7] ;
assign n13990 =  ( n13989 ) == ( bv_1_0_n53 )  ;
assign n13991 =  ( wr_addr ) == ( bv_8_85_n239 )  ;
assign n13992 =  ( n13990 ) & (n13991 )  ;
assign n13993 =  ( n13992 ) & (wr )  ;
assign n13994 =  ( n13993 ) ? ( n5449 ) : ( iram_85 ) ;
assign n13995 = wr_addr[7:7] ;
assign n13996 =  ( n13995 ) == ( bv_1_0_n53 )  ;
assign n13997 =  ( wr_addr ) == ( bv_8_85_n239 )  ;
assign n13998 =  ( n13996 ) & (n13997 )  ;
assign n13999 =  ( n13998 ) & (wr )  ;
assign n14000 =  ( n13999 ) ? ( n4906 ) : ( iram_85 ) ;
assign n14001 = wr_addr[7:7] ;
assign n14002 =  ( n14001 ) == ( bv_1_0_n53 )  ;
assign n14003 =  ( wr_addr ) == ( bv_8_85_n239 )  ;
assign n14004 =  ( n14002 ) & (n14003 )  ;
assign n14005 =  ( n14004 ) & (wr )  ;
assign n14006 =  ( n14005 ) ? ( n5485 ) : ( iram_85 ) ;
assign n14007 = wr_addr[7:7] ;
assign n14008 =  ( n14007 ) == ( bv_1_0_n53 )  ;
assign n14009 =  ( wr_addr ) == ( bv_8_85_n239 )  ;
assign n14010 =  ( n14008 ) & (n14009 )  ;
assign n14011 =  ( n14010 ) & (wr )  ;
assign n14012 =  ( n14011 ) ? ( n5512 ) : ( iram_85 ) ;
assign n14013 = wr_addr[7:7] ;
assign n14014 =  ( n14013 ) == ( bv_1_0_n53 )  ;
assign n14015 =  ( wr_addr ) == ( bv_8_85_n239 )  ;
assign n14016 =  ( n14014 ) & (n14015 )  ;
assign n14017 =  ( n14016 ) & (wr )  ;
assign n14018 =  ( n14017 ) ? ( bv_8_0_n69 ) : ( iram_85 ) ;
assign n14019 = wr_addr[7:7] ;
assign n14020 =  ( n14019 ) == ( bv_1_0_n53 )  ;
assign n14021 =  ( wr_addr ) == ( bv_8_85_n239 )  ;
assign n14022 =  ( n14020 ) & (n14021 )  ;
assign n14023 =  ( n14022 ) & (wr )  ;
assign n14024 =  ( n14023 ) ? ( n5071 ) : ( iram_85 ) ;
assign n14025 = wr_addr[7:7] ;
assign n14026 =  ( n14025 ) == ( bv_1_0_n53 )  ;
assign n14027 =  ( wr_addr ) == ( bv_8_85_n239 )  ;
assign n14028 =  ( n14026 ) & (n14027 )  ;
assign n14029 =  ( n14028 ) & (wr )  ;
assign n14030 =  ( n14029 ) ? ( n5096 ) : ( iram_85 ) ;
assign n14031 = wr_addr[7:7] ;
assign n14032 =  ( n14031 ) == ( bv_1_0_n53 )  ;
assign n14033 =  ( wr_addr ) == ( bv_8_85_n239 )  ;
assign n14034 =  ( n14032 ) & (n14033 )  ;
assign n14035 =  ( n14034 ) & (wr )  ;
assign n14036 =  ( n14035 ) ? ( n5123 ) : ( iram_85 ) ;
assign n14037 = wr_addr[7:7] ;
assign n14038 =  ( n14037 ) == ( bv_1_0_n53 )  ;
assign n14039 =  ( wr_addr ) == ( bv_8_85_n239 )  ;
assign n14040 =  ( n14038 ) & (n14039 )  ;
assign n14041 =  ( n14040 ) & (wr )  ;
assign n14042 =  ( n14041 ) ? ( n5165 ) : ( iram_85 ) ;
assign n14043 = wr_addr[7:7] ;
assign n14044 =  ( n14043 ) == ( bv_1_0_n53 )  ;
assign n14045 =  ( wr_addr ) == ( bv_8_85_n239 )  ;
assign n14046 =  ( n14044 ) & (n14045 )  ;
assign n14047 =  ( n14046 ) & (wr )  ;
assign n14048 =  ( n14047 ) ? ( n5204 ) : ( iram_85 ) ;
assign n14049 = wr_addr[7:7] ;
assign n14050 =  ( n14049 ) == ( bv_1_0_n53 )  ;
assign n14051 =  ( wr_addr ) == ( bv_8_85_n239 )  ;
assign n14052 =  ( n14050 ) & (n14051 )  ;
assign n14053 =  ( n14052 ) & (wr )  ;
assign n14054 =  ( n14053 ) ? ( n5262 ) : ( iram_85 ) ;
assign n14055 = wr_addr[7:7] ;
assign n14056 =  ( n14055 ) == ( bv_1_0_n53 )  ;
assign n14057 =  ( wr_addr ) == ( bv_8_85_n239 )  ;
assign n14058 =  ( n14056 ) & (n14057 )  ;
assign n14059 =  ( n14058 ) & (wr )  ;
assign n14060 =  ( n14059 ) ? ( n5298 ) : ( iram_85 ) ;
assign n14061 = wr_addr[7:7] ;
assign n14062 =  ( n14061 ) == ( bv_1_0_n53 )  ;
assign n14063 =  ( wr_addr ) == ( bv_8_85_n239 )  ;
assign n14064 =  ( n14062 ) & (n14063 )  ;
assign n14065 =  ( n14064 ) & (wr )  ;
assign n14066 =  ( n14065 ) ? ( n5325 ) : ( iram_85 ) ;
assign n14067 = wr_addr[7:7] ;
assign n14068 =  ( n14067 ) == ( bv_1_0_n53 )  ;
assign n14069 =  ( wr_addr ) == ( bv_8_86_n241 )  ;
assign n14070 =  ( n14068 ) & (n14069 )  ;
assign n14071 =  ( n14070 ) & (wr )  ;
assign n14072 =  ( n14071 ) ? ( n4782 ) : ( iram_86 ) ;
assign n14073 = wr_addr[7:7] ;
assign n14074 =  ( n14073 ) == ( bv_1_0_n53 )  ;
assign n14075 =  ( wr_addr ) == ( bv_8_86_n241 )  ;
assign n14076 =  ( n14074 ) & (n14075 )  ;
assign n14077 =  ( n14076 ) & (wr )  ;
assign n14078 =  ( n14077 ) ? ( n4841 ) : ( iram_86 ) ;
assign n14079 = wr_addr[7:7] ;
assign n14080 =  ( n14079 ) == ( bv_1_0_n53 )  ;
assign n14081 =  ( wr_addr ) == ( bv_8_86_n241 )  ;
assign n14082 =  ( n14080 ) & (n14081 )  ;
assign n14083 =  ( n14082 ) & (wr )  ;
assign n14084 =  ( n14083 ) ? ( n5449 ) : ( iram_86 ) ;
assign n14085 = wr_addr[7:7] ;
assign n14086 =  ( n14085 ) == ( bv_1_0_n53 )  ;
assign n14087 =  ( wr_addr ) == ( bv_8_86_n241 )  ;
assign n14088 =  ( n14086 ) & (n14087 )  ;
assign n14089 =  ( n14088 ) & (wr )  ;
assign n14090 =  ( n14089 ) ? ( n4906 ) : ( iram_86 ) ;
assign n14091 = wr_addr[7:7] ;
assign n14092 =  ( n14091 ) == ( bv_1_0_n53 )  ;
assign n14093 =  ( wr_addr ) == ( bv_8_86_n241 )  ;
assign n14094 =  ( n14092 ) & (n14093 )  ;
assign n14095 =  ( n14094 ) & (wr )  ;
assign n14096 =  ( n14095 ) ? ( n5485 ) : ( iram_86 ) ;
assign n14097 = wr_addr[7:7] ;
assign n14098 =  ( n14097 ) == ( bv_1_0_n53 )  ;
assign n14099 =  ( wr_addr ) == ( bv_8_86_n241 )  ;
assign n14100 =  ( n14098 ) & (n14099 )  ;
assign n14101 =  ( n14100 ) & (wr )  ;
assign n14102 =  ( n14101 ) ? ( n5512 ) : ( iram_86 ) ;
assign n14103 = wr_addr[7:7] ;
assign n14104 =  ( n14103 ) == ( bv_1_0_n53 )  ;
assign n14105 =  ( wr_addr ) == ( bv_8_86_n241 )  ;
assign n14106 =  ( n14104 ) & (n14105 )  ;
assign n14107 =  ( n14106 ) & (wr )  ;
assign n14108 =  ( n14107 ) ? ( bv_8_0_n69 ) : ( iram_86 ) ;
assign n14109 = wr_addr[7:7] ;
assign n14110 =  ( n14109 ) == ( bv_1_0_n53 )  ;
assign n14111 =  ( wr_addr ) == ( bv_8_86_n241 )  ;
assign n14112 =  ( n14110 ) & (n14111 )  ;
assign n14113 =  ( n14112 ) & (wr )  ;
assign n14114 =  ( n14113 ) ? ( n5071 ) : ( iram_86 ) ;
assign n14115 = wr_addr[7:7] ;
assign n14116 =  ( n14115 ) == ( bv_1_0_n53 )  ;
assign n14117 =  ( wr_addr ) == ( bv_8_86_n241 )  ;
assign n14118 =  ( n14116 ) & (n14117 )  ;
assign n14119 =  ( n14118 ) & (wr )  ;
assign n14120 =  ( n14119 ) ? ( n5096 ) : ( iram_86 ) ;
assign n14121 = wr_addr[7:7] ;
assign n14122 =  ( n14121 ) == ( bv_1_0_n53 )  ;
assign n14123 =  ( wr_addr ) == ( bv_8_86_n241 )  ;
assign n14124 =  ( n14122 ) & (n14123 )  ;
assign n14125 =  ( n14124 ) & (wr )  ;
assign n14126 =  ( n14125 ) ? ( n5123 ) : ( iram_86 ) ;
assign n14127 = wr_addr[7:7] ;
assign n14128 =  ( n14127 ) == ( bv_1_0_n53 )  ;
assign n14129 =  ( wr_addr ) == ( bv_8_86_n241 )  ;
assign n14130 =  ( n14128 ) & (n14129 )  ;
assign n14131 =  ( n14130 ) & (wr )  ;
assign n14132 =  ( n14131 ) ? ( n5165 ) : ( iram_86 ) ;
assign n14133 = wr_addr[7:7] ;
assign n14134 =  ( n14133 ) == ( bv_1_0_n53 )  ;
assign n14135 =  ( wr_addr ) == ( bv_8_86_n241 )  ;
assign n14136 =  ( n14134 ) & (n14135 )  ;
assign n14137 =  ( n14136 ) & (wr )  ;
assign n14138 =  ( n14137 ) ? ( n5204 ) : ( iram_86 ) ;
assign n14139 = wr_addr[7:7] ;
assign n14140 =  ( n14139 ) == ( bv_1_0_n53 )  ;
assign n14141 =  ( wr_addr ) == ( bv_8_86_n241 )  ;
assign n14142 =  ( n14140 ) & (n14141 )  ;
assign n14143 =  ( n14142 ) & (wr )  ;
assign n14144 =  ( n14143 ) ? ( n5262 ) : ( iram_86 ) ;
assign n14145 = wr_addr[7:7] ;
assign n14146 =  ( n14145 ) == ( bv_1_0_n53 )  ;
assign n14147 =  ( wr_addr ) == ( bv_8_86_n241 )  ;
assign n14148 =  ( n14146 ) & (n14147 )  ;
assign n14149 =  ( n14148 ) & (wr )  ;
assign n14150 =  ( n14149 ) ? ( n5298 ) : ( iram_86 ) ;
assign n14151 = wr_addr[7:7] ;
assign n14152 =  ( n14151 ) == ( bv_1_0_n53 )  ;
assign n14153 =  ( wr_addr ) == ( bv_8_86_n241 )  ;
assign n14154 =  ( n14152 ) & (n14153 )  ;
assign n14155 =  ( n14154 ) & (wr )  ;
assign n14156 =  ( n14155 ) ? ( n5325 ) : ( iram_86 ) ;
assign n14157 = wr_addr[7:7] ;
assign n14158 =  ( n14157 ) == ( bv_1_0_n53 )  ;
assign n14159 =  ( wr_addr ) == ( bv_8_87_n243 )  ;
assign n14160 =  ( n14158 ) & (n14159 )  ;
assign n14161 =  ( n14160 ) & (wr )  ;
assign n14162 =  ( n14161 ) ? ( n4782 ) : ( iram_87 ) ;
assign n14163 = wr_addr[7:7] ;
assign n14164 =  ( n14163 ) == ( bv_1_0_n53 )  ;
assign n14165 =  ( wr_addr ) == ( bv_8_87_n243 )  ;
assign n14166 =  ( n14164 ) & (n14165 )  ;
assign n14167 =  ( n14166 ) & (wr )  ;
assign n14168 =  ( n14167 ) ? ( n4841 ) : ( iram_87 ) ;
assign n14169 = wr_addr[7:7] ;
assign n14170 =  ( n14169 ) == ( bv_1_0_n53 )  ;
assign n14171 =  ( wr_addr ) == ( bv_8_87_n243 )  ;
assign n14172 =  ( n14170 ) & (n14171 )  ;
assign n14173 =  ( n14172 ) & (wr )  ;
assign n14174 =  ( n14173 ) ? ( n5449 ) : ( iram_87 ) ;
assign n14175 = wr_addr[7:7] ;
assign n14176 =  ( n14175 ) == ( bv_1_0_n53 )  ;
assign n14177 =  ( wr_addr ) == ( bv_8_87_n243 )  ;
assign n14178 =  ( n14176 ) & (n14177 )  ;
assign n14179 =  ( n14178 ) & (wr )  ;
assign n14180 =  ( n14179 ) ? ( n4906 ) : ( iram_87 ) ;
assign n14181 = wr_addr[7:7] ;
assign n14182 =  ( n14181 ) == ( bv_1_0_n53 )  ;
assign n14183 =  ( wr_addr ) == ( bv_8_87_n243 )  ;
assign n14184 =  ( n14182 ) & (n14183 )  ;
assign n14185 =  ( n14184 ) & (wr )  ;
assign n14186 =  ( n14185 ) ? ( n5485 ) : ( iram_87 ) ;
assign n14187 = wr_addr[7:7] ;
assign n14188 =  ( n14187 ) == ( bv_1_0_n53 )  ;
assign n14189 =  ( wr_addr ) == ( bv_8_87_n243 )  ;
assign n14190 =  ( n14188 ) & (n14189 )  ;
assign n14191 =  ( n14190 ) & (wr )  ;
assign n14192 =  ( n14191 ) ? ( n5512 ) : ( iram_87 ) ;
assign n14193 = wr_addr[7:7] ;
assign n14194 =  ( n14193 ) == ( bv_1_0_n53 )  ;
assign n14195 =  ( wr_addr ) == ( bv_8_87_n243 )  ;
assign n14196 =  ( n14194 ) & (n14195 )  ;
assign n14197 =  ( n14196 ) & (wr )  ;
assign n14198 =  ( n14197 ) ? ( bv_8_0_n69 ) : ( iram_87 ) ;
assign n14199 = wr_addr[7:7] ;
assign n14200 =  ( n14199 ) == ( bv_1_0_n53 )  ;
assign n14201 =  ( wr_addr ) == ( bv_8_87_n243 )  ;
assign n14202 =  ( n14200 ) & (n14201 )  ;
assign n14203 =  ( n14202 ) & (wr )  ;
assign n14204 =  ( n14203 ) ? ( n5071 ) : ( iram_87 ) ;
assign n14205 = wr_addr[7:7] ;
assign n14206 =  ( n14205 ) == ( bv_1_0_n53 )  ;
assign n14207 =  ( wr_addr ) == ( bv_8_87_n243 )  ;
assign n14208 =  ( n14206 ) & (n14207 )  ;
assign n14209 =  ( n14208 ) & (wr )  ;
assign n14210 =  ( n14209 ) ? ( n5096 ) : ( iram_87 ) ;
assign n14211 = wr_addr[7:7] ;
assign n14212 =  ( n14211 ) == ( bv_1_0_n53 )  ;
assign n14213 =  ( wr_addr ) == ( bv_8_87_n243 )  ;
assign n14214 =  ( n14212 ) & (n14213 )  ;
assign n14215 =  ( n14214 ) & (wr )  ;
assign n14216 =  ( n14215 ) ? ( n5123 ) : ( iram_87 ) ;
assign n14217 = wr_addr[7:7] ;
assign n14218 =  ( n14217 ) == ( bv_1_0_n53 )  ;
assign n14219 =  ( wr_addr ) == ( bv_8_87_n243 )  ;
assign n14220 =  ( n14218 ) & (n14219 )  ;
assign n14221 =  ( n14220 ) & (wr )  ;
assign n14222 =  ( n14221 ) ? ( n5165 ) : ( iram_87 ) ;
assign n14223 = wr_addr[7:7] ;
assign n14224 =  ( n14223 ) == ( bv_1_0_n53 )  ;
assign n14225 =  ( wr_addr ) == ( bv_8_87_n243 )  ;
assign n14226 =  ( n14224 ) & (n14225 )  ;
assign n14227 =  ( n14226 ) & (wr )  ;
assign n14228 =  ( n14227 ) ? ( n5204 ) : ( iram_87 ) ;
assign n14229 = wr_addr[7:7] ;
assign n14230 =  ( n14229 ) == ( bv_1_0_n53 )  ;
assign n14231 =  ( wr_addr ) == ( bv_8_87_n243 )  ;
assign n14232 =  ( n14230 ) & (n14231 )  ;
assign n14233 =  ( n14232 ) & (wr )  ;
assign n14234 =  ( n14233 ) ? ( n5262 ) : ( iram_87 ) ;
assign n14235 = wr_addr[7:7] ;
assign n14236 =  ( n14235 ) == ( bv_1_0_n53 )  ;
assign n14237 =  ( wr_addr ) == ( bv_8_87_n243 )  ;
assign n14238 =  ( n14236 ) & (n14237 )  ;
assign n14239 =  ( n14238 ) & (wr )  ;
assign n14240 =  ( n14239 ) ? ( n5298 ) : ( iram_87 ) ;
assign n14241 = wr_addr[7:7] ;
assign n14242 =  ( n14241 ) == ( bv_1_0_n53 )  ;
assign n14243 =  ( wr_addr ) == ( bv_8_87_n243 )  ;
assign n14244 =  ( n14242 ) & (n14243 )  ;
assign n14245 =  ( n14244 ) & (wr )  ;
assign n14246 =  ( n14245 ) ? ( n5325 ) : ( iram_87 ) ;
assign n14247 = wr_addr[7:7] ;
assign n14248 =  ( n14247 ) == ( bv_1_0_n53 )  ;
assign n14249 =  ( wr_addr ) == ( bv_8_88_n245 )  ;
assign n14250 =  ( n14248 ) & (n14249 )  ;
assign n14251 =  ( n14250 ) & (wr )  ;
assign n14252 =  ( n14251 ) ? ( n4782 ) : ( iram_88 ) ;
assign n14253 = wr_addr[7:7] ;
assign n14254 =  ( n14253 ) == ( bv_1_0_n53 )  ;
assign n14255 =  ( wr_addr ) == ( bv_8_88_n245 )  ;
assign n14256 =  ( n14254 ) & (n14255 )  ;
assign n14257 =  ( n14256 ) & (wr )  ;
assign n14258 =  ( n14257 ) ? ( n4841 ) : ( iram_88 ) ;
assign n14259 = wr_addr[7:7] ;
assign n14260 =  ( n14259 ) == ( bv_1_0_n53 )  ;
assign n14261 =  ( wr_addr ) == ( bv_8_88_n245 )  ;
assign n14262 =  ( n14260 ) & (n14261 )  ;
assign n14263 =  ( n14262 ) & (wr )  ;
assign n14264 =  ( n14263 ) ? ( n5449 ) : ( iram_88 ) ;
assign n14265 = wr_addr[7:7] ;
assign n14266 =  ( n14265 ) == ( bv_1_0_n53 )  ;
assign n14267 =  ( wr_addr ) == ( bv_8_88_n245 )  ;
assign n14268 =  ( n14266 ) & (n14267 )  ;
assign n14269 =  ( n14268 ) & (wr )  ;
assign n14270 =  ( n14269 ) ? ( n4906 ) : ( iram_88 ) ;
assign n14271 = wr_addr[7:7] ;
assign n14272 =  ( n14271 ) == ( bv_1_0_n53 )  ;
assign n14273 =  ( wr_addr ) == ( bv_8_88_n245 )  ;
assign n14274 =  ( n14272 ) & (n14273 )  ;
assign n14275 =  ( n14274 ) & (wr )  ;
assign n14276 =  ( n14275 ) ? ( n5485 ) : ( iram_88 ) ;
assign n14277 = wr_addr[7:7] ;
assign n14278 =  ( n14277 ) == ( bv_1_0_n53 )  ;
assign n14279 =  ( wr_addr ) == ( bv_8_88_n245 )  ;
assign n14280 =  ( n14278 ) & (n14279 )  ;
assign n14281 =  ( n14280 ) & (wr )  ;
assign n14282 =  ( n14281 ) ? ( n5512 ) : ( iram_88 ) ;
assign n14283 = wr_addr[7:7] ;
assign n14284 =  ( n14283 ) == ( bv_1_0_n53 )  ;
assign n14285 =  ( wr_addr ) == ( bv_8_88_n245 )  ;
assign n14286 =  ( n14284 ) & (n14285 )  ;
assign n14287 =  ( n14286 ) & (wr )  ;
assign n14288 =  ( n14287 ) ? ( bv_8_0_n69 ) : ( iram_88 ) ;
assign n14289 = wr_addr[7:7] ;
assign n14290 =  ( n14289 ) == ( bv_1_0_n53 )  ;
assign n14291 =  ( wr_addr ) == ( bv_8_88_n245 )  ;
assign n14292 =  ( n14290 ) & (n14291 )  ;
assign n14293 =  ( n14292 ) & (wr )  ;
assign n14294 =  ( n14293 ) ? ( n5071 ) : ( iram_88 ) ;
assign n14295 = wr_addr[7:7] ;
assign n14296 =  ( n14295 ) == ( bv_1_0_n53 )  ;
assign n14297 =  ( wr_addr ) == ( bv_8_88_n245 )  ;
assign n14298 =  ( n14296 ) & (n14297 )  ;
assign n14299 =  ( n14298 ) & (wr )  ;
assign n14300 =  ( n14299 ) ? ( n5096 ) : ( iram_88 ) ;
assign n14301 = wr_addr[7:7] ;
assign n14302 =  ( n14301 ) == ( bv_1_0_n53 )  ;
assign n14303 =  ( wr_addr ) == ( bv_8_88_n245 )  ;
assign n14304 =  ( n14302 ) & (n14303 )  ;
assign n14305 =  ( n14304 ) & (wr )  ;
assign n14306 =  ( n14305 ) ? ( n5123 ) : ( iram_88 ) ;
assign n14307 = wr_addr[7:7] ;
assign n14308 =  ( n14307 ) == ( bv_1_0_n53 )  ;
assign n14309 =  ( wr_addr ) == ( bv_8_88_n245 )  ;
assign n14310 =  ( n14308 ) & (n14309 )  ;
assign n14311 =  ( n14310 ) & (wr )  ;
assign n14312 =  ( n14311 ) ? ( n5165 ) : ( iram_88 ) ;
assign n14313 = wr_addr[7:7] ;
assign n14314 =  ( n14313 ) == ( bv_1_0_n53 )  ;
assign n14315 =  ( wr_addr ) == ( bv_8_88_n245 )  ;
assign n14316 =  ( n14314 ) & (n14315 )  ;
assign n14317 =  ( n14316 ) & (wr )  ;
assign n14318 =  ( n14317 ) ? ( n5204 ) : ( iram_88 ) ;
assign n14319 = wr_addr[7:7] ;
assign n14320 =  ( n14319 ) == ( bv_1_0_n53 )  ;
assign n14321 =  ( wr_addr ) == ( bv_8_88_n245 )  ;
assign n14322 =  ( n14320 ) & (n14321 )  ;
assign n14323 =  ( n14322 ) & (wr )  ;
assign n14324 =  ( n14323 ) ? ( n5262 ) : ( iram_88 ) ;
assign n14325 = wr_addr[7:7] ;
assign n14326 =  ( n14325 ) == ( bv_1_0_n53 )  ;
assign n14327 =  ( wr_addr ) == ( bv_8_88_n245 )  ;
assign n14328 =  ( n14326 ) & (n14327 )  ;
assign n14329 =  ( n14328 ) & (wr )  ;
assign n14330 =  ( n14329 ) ? ( n5298 ) : ( iram_88 ) ;
assign n14331 = wr_addr[7:7] ;
assign n14332 =  ( n14331 ) == ( bv_1_0_n53 )  ;
assign n14333 =  ( wr_addr ) == ( bv_8_88_n245 )  ;
assign n14334 =  ( n14332 ) & (n14333 )  ;
assign n14335 =  ( n14334 ) & (wr )  ;
assign n14336 =  ( n14335 ) ? ( n5325 ) : ( iram_88 ) ;
assign n14337 = wr_addr[7:7] ;
assign n14338 =  ( n14337 ) == ( bv_1_0_n53 )  ;
assign n14339 =  ( wr_addr ) == ( bv_8_89_n247 )  ;
assign n14340 =  ( n14338 ) & (n14339 )  ;
assign n14341 =  ( n14340 ) & (wr )  ;
assign n14342 =  ( n14341 ) ? ( n4782 ) : ( iram_89 ) ;
assign n14343 = wr_addr[7:7] ;
assign n14344 =  ( n14343 ) == ( bv_1_0_n53 )  ;
assign n14345 =  ( wr_addr ) == ( bv_8_89_n247 )  ;
assign n14346 =  ( n14344 ) & (n14345 )  ;
assign n14347 =  ( n14346 ) & (wr )  ;
assign n14348 =  ( n14347 ) ? ( n4841 ) : ( iram_89 ) ;
assign n14349 = wr_addr[7:7] ;
assign n14350 =  ( n14349 ) == ( bv_1_0_n53 )  ;
assign n14351 =  ( wr_addr ) == ( bv_8_89_n247 )  ;
assign n14352 =  ( n14350 ) & (n14351 )  ;
assign n14353 =  ( n14352 ) & (wr )  ;
assign n14354 =  ( n14353 ) ? ( n5449 ) : ( iram_89 ) ;
assign n14355 = wr_addr[7:7] ;
assign n14356 =  ( n14355 ) == ( bv_1_0_n53 )  ;
assign n14357 =  ( wr_addr ) == ( bv_8_89_n247 )  ;
assign n14358 =  ( n14356 ) & (n14357 )  ;
assign n14359 =  ( n14358 ) & (wr )  ;
assign n14360 =  ( n14359 ) ? ( n4906 ) : ( iram_89 ) ;
assign n14361 = wr_addr[7:7] ;
assign n14362 =  ( n14361 ) == ( bv_1_0_n53 )  ;
assign n14363 =  ( wr_addr ) == ( bv_8_89_n247 )  ;
assign n14364 =  ( n14362 ) & (n14363 )  ;
assign n14365 =  ( n14364 ) & (wr )  ;
assign n14366 =  ( n14365 ) ? ( n5485 ) : ( iram_89 ) ;
assign n14367 = wr_addr[7:7] ;
assign n14368 =  ( n14367 ) == ( bv_1_0_n53 )  ;
assign n14369 =  ( wr_addr ) == ( bv_8_89_n247 )  ;
assign n14370 =  ( n14368 ) & (n14369 )  ;
assign n14371 =  ( n14370 ) & (wr )  ;
assign n14372 =  ( n14371 ) ? ( n5512 ) : ( iram_89 ) ;
assign n14373 = wr_addr[7:7] ;
assign n14374 =  ( n14373 ) == ( bv_1_0_n53 )  ;
assign n14375 =  ( wr_addr ) == ( bv_8_89_n247 )  ;
assign n14376 =  ( n14374 ) & (n14375 )  ;
assign n14377 =  ( n14376 ) & (wr )  ;
assign n14378 =  ( n14377 ) ? ( bv_8_0_n69 ) : ( iram_89 ) ;
assign n14379 = wr_addr[7:7] ;
assign n14380 =  ( n14379 ) == ( bv_1_0_n53 )  ;
assign n14381 =  ( wr_addr ) == ( bv_8_89_n247 )  ;
assign n14382 =  ( n14380 ) & (n14381 )  ;
assign n14383 =  ( n14382 ) & (wr )  ;
assign n14384 =  ( n14383 ) ? ( n5071 ) : ( iram_89 ) ;
assign n14385 = wr_addr[7:7] ;
assign n14386 =  ( n14385 ) == ( bv_1_0_n53 )  ;
assign n14387 =  ( wr_addr ) == ( bv_8_89_n247 )  ;
assign n14388 =  ( n14386 ) & (n14387 )  ;
assign n14389 =  ( n14388 ) & (wr )  ;
assign n14390 =  ( n14389 ) ? ( n5096 ) : ( iram_89 ) ;
assign n14391 = wr_addr[7:7] ;
assign n14392 =  ( n14391 ) == ( bv_1_0_n53 )  ;
assign n14393 =  ( wr_addr ) == ( bv_8_89_n247 )  ;
assign n14394 =  ( n14392 ) & (n14393 )  ;
assign n14395 =  ( n14394 ) & (wr )  ;
assign n14396 =  ( n14395 ) ? ( n5123 ) : ( iram_89 ) ;
assign n14397 = wr_addr[7:7] ;
assign n14398 =  ( n14397 ) == ( bv_1_0_n53 )  ;
assign n14399 =  ( wr_addr ) == ( bv_8_89_n247 )  ;
assign n14400 =  ( n14398 ) & (n14399 )  ;
assign n14401 =  ( n14400 ) & (wr )  ;
assign n14402 =  ( n14401 ) ? ( n5165 ) : ( iram_89 ) ;
assign n14403 = wr_addr[7:7] ;
assign n14404 =  ( n14403 ) == ( bv_1_0_n53 )  ;
assign n14405 =  ( wr_addr ) == ( bv_8_89_n247 )  ;
assign n14406 =  ( n14404 ) & (n14405 )  ;
assign n14407 =  ( n14406 ) & (wr )  ;
assign n14408 =  ( n14407 ) ? ( n5204 ) : ( iram_89 ) ;
assign n14409 = wr_addr[7:7] ;
assign n14410 =  ( n14409 ) == ( bv_1_0_n53 )  ;
assign n14411 =  ( wr_addr ) == ( bv_8_89_n247 )  ;
assign n14412 =  ( n14410 ) & (n14411 )  ;
assign n14413 =  ( n14412 ) & (wr )  ;
assign n14414 =  ( n14413 ) ? ( n5262 ) : ( iram_89 ) ;
assign n14415 = wr_addr[7:7] ;
assign n14416 =  ( n14415 ) == ( bv_1_0_n53 )  ;
assign n14417 =  ( wr_addr ) == ( bv_8_89_n247 )  ;
assign n14418 =  ( n14416 ) & (n14417 )  ;
assign n14419 =  ( n14418 ) & (wr )  ;
assign n14420 =  ( n14419 ) ? ( n5298 ) : ( iram_89 ) ;
assign n14421 = wr_addr[7:7] ;
assign n14422 =  ( n14421 ) == ( bv_1_0_n53 )  ;
assign n14423 =  ( wr_addr ) == ( bv_8_89_n247 )  ;
assign n14424 =  ( n14422 ) & (n14423 )  ;
assign n14425 =  ( n14424 ) & (wr )  ;
assign n14426 =  ( n14425 ) ? ( n5325 ) : ( iram_89 ) ;
assign n14427 = wr_addr[7:7] ;
assign n14428 =  ( n14427 ) == ( bv_1_0_n53 )  ;
assign n14429 =  ( wr_addr ) == ( bv_8_90_n249 )  ;
assign n14430 =  ( n14428 ) & (n14429 )  ;
assign n14431 =  ( n14430 ) & (wr )  ;
assign n14432 =  ( n14431 ) ? ( n4782 ) : ( iram_90 ) ;
assign n14433 = wr_addr[7:7] ;
assign n14434 =  ( n14433 ) == ( bv_1_0_n53 )  ;
assign n14435 =  ( wr_addr ) == ( bv_8_90_n249 )  ;
assign n14436 =  ( n14434 ) & (n14435 )  ;
assign n14437 =  ( n14436 ) & (wr )  ;
assign n14438 =  ( n14437 ) ? ( n4841 ) : ( iram_90 ) ;
assign n14439 = wr_addr[7:7] ;
assign n14440 =  ( n14439 ) == ( bv_1_0_n53 )  ;
assign n14441 =  ( wr_addr ) == ( bv_8_90_n249 )  ;
assign n14442 =  ( n14440 ) & (n14441 )  ;
assign n14443 =  ( n14442 ) & (wr )  ;
assign n14444 =  ( n14443 ) ? ( n5449 ) : ( iram_90 ) ;
assign n14445 = wr_addr[7:7] ;
assign n14446 =  ( n14445 ) == ( bv_1_0_n53 )  ;
assign n14447 =  ( wr_addr ) == ( bv_8_90_n249 )  ;
assign n14448 =  ( n14446 ) & (n14447 )  ;
assign n14449 =  ( n14448 ) & (wr )  ;
assign n14450 =  ( n14449 ) ? ( n4906 ) : ( iram_90 ) ;
assign n14451 = wr_addr[7:7] ;
assign n14452 =  ( n14451 ) == ( bv_1_0_n53 )  ;
assign n14453 =  ( wr_addr ) == ( bv_8_90_n249 )  ;
assign n14454 =  ( n14452 ) & (n14453 )  ;
assign n14455 =  ( n14454 ) & (wr )  ;
assign n14456 =  ( n14455 ) ? ( n5485 ) : ( iram_90 ) ;
assign n14457 = wr_addr[7:7] ;
assign n14458 =  ( n14457 ) == ( bv_1_0_n53 )  ;
assign n14459 =  ( wr_addr ) == ( bv_8_90_n249 )  ;
assign n14460 =  ( n14458 ) & (n14459 )  ;
assign n14461 =  ( n14460 ) & (wr )  ;
assign n14462 =  ( n14461 ) ? ( n5512 ) : ( iram_90 ) ;
assign n14463 = wr_addr[7:7] ;
assign n14464 =  ( n14463 ) == ( bv_1_0_n53 )  ;
assign n14465 =  ( wr_addr ) == ( bv_8_90_n249 )  ;
assign n14466 =  ( n14464 ) & (n14465 )  ;
assign n14467 =  ( n14466 ) & (wr )  ;
assign n14468 =  ( n14467 ) ? ( bv_8_0_n69 ) : ( iram_90 ) ;
assign n14469 = wr_addr[7:7] ;
assign n14470 =  ( n14469 ) == ( bv_1_0_n53 )  ;
assign n14471 =  ( wr_addr ) == ( bv_8_90_n249 )  ;
assign n14472 =  ( n14470 ) & (n14471 )  ;
assign n14473 =  ( n14472 ) & (wr )  ;
assign n14474 =  ( n14473 ) ? ( n5071 ) : ( iram_90 ) ;
assign n14475 = wr_addr[7:7] ;
assign n14476 =  ( n14475 ) == ( bv_1_0_n53 )  ;
assign n14477 =  ( wr_addr ) == ( bv_8_90_n249 )  ;
assign n14478 =  ( n14476 ) & (n14477 )  ;
assign n14479 =  ( n14478 ) & (wr )  ;
assign n14480 =  ( n14479 ) ? ( n5096 ) : ( iram_90 ) ;
assign n14481 = wr_addr[7:7] ;
assign n14482 =  ( n14481 ) == ( bv_1_0_n53 )  ;
assign n14483 =  ( wr_addr ) == ( bv_8_90_n249 )  ;
assign n14484 =  ( n14482 ) & (n14483 )  ;
assign n14485 =  ( n14484 ) & (wr )  ;
assign n14486 =  ( n14485 ) ? ( n5123 ) : ( iram_90 ) ;
assign n14487 = wr_addr[7:7] ;
assign n14488 =  ( n14487 ) == ( bv_1_0_n53 )  ;
assign n14489 =  ( wr_addr ) == ( bv_8_90_n249 )  ;
assign n14490 =  ( n14488 ) & (n14489 )  ;
assign n14491 =  ( n14490 ) & (wr )  ;
assign n14492 =  ( n14491 ) ? ( n5165 ) : ( iram_90 ) ;
assign n14493 = wr_addr[7:7] ;
assign n14494 =  ( n14493 ) == ( bv_1_0_n53 )  ;
assign n14495 =  ( wr_addr ) == ( bv_8_90_n249 )  ;
assign n14496 =  ( n14494 ) & (n14495 )  ;
assign n14497 =  ( n14496 ) & (wr )  ;
assign n14498 =  ( n14497 ) ? ( n5204 ) : ( iram_90 ) ;
assign n14499 = wr_addr[7:7] ;
assign n14500 =  ( n14499 ) == ( bv_1_0_n53 )  ;
assign n14501 =  ( wr_addr ) == ( bv_8_90_n249 )  ;
assign n14502 =  ( n14500 ) & (n14501 )  ;
assign n14503 =  ( n14502 ) & (wr )  ;
assign n14504 =  ( n14503 ) ? ( n5262 ) : ( iram_90 ) ;
assign n14505 = wr_addr[7:7] ;
assign n14506 =  ( n14505 ) == ( bv_1_0_n53 )  ;
assign n14507 =  ( wr_addr ) == ( bv_8_90_n249 )  ;
assign n14508 =  ( n14506 ) & (n14507 )  ;
assign n14509 =  ( n14508 ) & (wr )  ;
assign n14510 =  ( n14509 ) ? ( n5298 ) : ( iram_90 ) ;
assign n14511 = wr_addr[7:7] ;
assign n14512 =  ( n14511 ) == ( bv_1_0_n53 )  ;
assign n14513 =  ( wr_addr ) == ( bv_8_90_n249 )  ;
assign n14514 =  ( n14512 ) & (n14513 )  ;
assign n14515 =  ( n14514 ) & (wr )  ;
assign n14516 =  ( n14515 ) ? ( n5325 ) : ( iram_90 ) ;
assign n14517 = wr_addr[7:7] ;
assign n14518 =  ( n14517 ) == ( bv_1_0_n53 )  ;
assign n14519 =  ( wr_addr ) == ( bv_8_91_n251 )  ;
assign n14520 =  ( n14518 ) & (n14519 )  ;
assign n14521 =  ( n14520 ) & (wr )  ;
assign n14522 =  ( n14521 ) ? ( n4782 ) : ( iram_91 ) ;
assign n14523 = wr_addr[7:7] ;
assign n14524 =  ( n14523 ) == ( bv_1_0_n53 )  ;
assign n14525 =  ( wr_addr ) == ( bv_8_91_n251 )  ;
assign n14526 =  ( n14524 ) & (n14525 )  ;
assign n14527 =  ( n14526 ) & (wr )  ;
assign n14528 =  ( n14527 ) ? ( n4841 ) : ( iram_91 ) ;
assign n14529 = wr_addr[7:7] ;
assign n14530 =  ( n14529 ) == ( bv_1_0_n53 )  ;
assign n14531 =  ( wr_addr ) == ( bv_8_91_n251 )  ;
assign n14532 =  ( n14530 ) & (n14531 )  ;
assign n14533 =  ( n14532 ) & (wr )  ;
assign n14534 =  ( n14533 ) ? ( n5449 ) : ( iram_91 ) ;
assign n14535 = wr_addr[7:7] ;
assign n14536 =  ( n14535 ) == ( bv_1_0_n53 )  ;
assign n14537 =  ( wr_addr ) == ( bv_8_91_n251 )  ;
assign n14538 =  ( n14536 ) & (n14537 )  ;
assign n14539 =  ( n14538 ) & (wr )  ;
assign n14540 =  ( n14539 ) ? ( n4906 ) : ( iram_91 ) ;
assign n14541 = wr_addr[7:7] ;
assign n14542 =  ( n14541 ) == ( bv_1_0_n53 )  ;
assign n14543 =  ( wr_addr ) == ( bv_8_91_n251 )  ;
assign n14544 =  ( n14542 ) & (n14543 )  ;
assign n14545 =  ( n14544 ) & (wr )  ;
assign n14546 =  ( n14545 ) ? ( n5485 ) : ( iram_91 ) ;
assign n14547 = wr_addr[7:7] ;
assign n14548 =  ( n14547 ) == ( bv_1_0_n53 )  ;
assign n14549 =  ( wr_addr ) == ( bv_8_91_n251 )  ;
assign n14550 =  ( n14548 ) & (n14549 )  ;
assign n14551 =  ( n14550 ) & (wr )  ;
assign n14552 =  ( n14551 ) ? ( n5512 ) : ( iram_91 ) ;
assign n14553 = wr_addr[7:7] ;
assign n14554 =  ( n14553 ) == ( bv_1_0_n53 )  ;
assign n14555 =  ( wr_addr ) == ( bv_8_91_n251 )  ;
assign n14556 =  ( n14554 ) & (n14555 )  ;
assign n14557 =  ( n14556 ) & (wr )  ;
assign n14558 =  ( n14557 ) ? ( bv_8_0_n69 ) : ( iram_91 ) ;
assign n14559 = wr_addr[7:7] ;
assign n14560 =  ( n14559 ) == ( bv_1_0_n53 )  ;
assign n14561 =  ( wr_addr ) == ( bv_8_91_n251 )  ;
assign n14562 =  ( n14560 ) & (n14561 )  ;
assign n14563 =  ( n14562 ) & (wr )  ;
assign n14564 =  ( n14563 ) ? ( n5071 ) : ( iram_91 ) ;
assign n14565 = wr_addr[7:7] ;
assign n14566 =  ( n14565 ) == ( bv_1_0_n53 )  ;
assign n14567 =  ( wr_addr ) == ( bv_8_91_n251 )  ;
assign n14568 =  ( n14566 ) & (n14567 )  ;
assign n14569 =  ( n14568 ) & (wr )  ;
assign n14570 =  ( n14569 ) ? ( n5096 ) : ( iram_91 ) ;
assign n14571 = wr_addr[7:7] ;
assign n14572 =  ( n14571 ) == ( bv_1_0_n53 )  ;
assign n14573 =  ( wr_addr ) == ( bv_8_91_n251 )  ;
assign n14574 =  ( n14572 ) & (n14573 )  ;
assign n14575 =  ( n14574 ) & (wr )  ;
assign n14576 =  ( n14575 ) ? ( n5123 ) : ( iram_91 ) ;
assign n14577 = wr_addr[7:7] ;
assign n14578 =  ( n14577 ) == ( bv_1_0_n53 )  ;
assign n14579 =  ( wr_addr ) == ( bv_8_91_n251 )  ;
assign n14580 =  ( n14578 ) & (n14579 )  ;
assign n14581 =  ( n14580 ) & (wr )  ;
assign n14582 =  ( n14581 ) ? ( n5165 ) : ( iram_91 ) ;
assign n14583 = wr_addr[7:7] ;
assign n14584 =  ( n14583 ) == ( bv_1_0_n53 )  ;
assign n14585 =  ( wr_addr ) == ( bv_8_91_n251 )  ;
assign n14586 =  ( n14584 ) & (n14585 )  ;
assign n14587 =  ( n14586 ) & (wr )  ;
assign n14588 =  ( n14587 ) ? ( n5204 ) : ( iram_91 ) ;
assign n14589 = wr_addr[7:7] ;
assign n14590 =  ( n14589 ) == ( bv_1_0_n53 )  ;
assign n14591 =  ( wr_addr ) == ( bv_8_91_n251 )  ;
assign n14592 =  ( n14590 ) & (n14591 )  ;
assign n14593 =  ( n14592 ) & (wr )  ;
assign n14594 =  ( n14593 ) ? ( n5262 ) : ( iram_91 ) ;
assign n14595 = wr_addr[7:7] ;
assign n14596 =  ( n14595 ) == ( bv_1_0_n53 )  ;
assign n14597 =  ( wr_addr ) == ( bv_8_91_n251 )  ;
assign n14598 =  ( n14596 ) & (n14597 )  ;
assign n14599 =  ( n14598 ) & (wr )  ;
assign n14600 =  ( n14599 ) ? ( n5298 ) : ( iram_91 ) ;
assign n14601 = wr_addr[7:7] ;
assign n14602 =  ( n14601 ) == ( bv_1_0_n53 )  ;
assign n14603 =  ( wr_addr ) == ( bv_8_91_n251 )  ;
assign n14604 =  ( n14602 ) & (n14603 )  ;
assign n14605 =  ( n14604 ) & (wr )  ;
assign n14606 =  ( n14605 ) ? ( n5325 ) : ( iram_91 ) ;
assign n14607 = wr_addr[7:7] ;
assign n14608 =  ( n14607 ) == ( bv_1_0_n53 )  ;
assign n14609 =  ( wr_addr ) == ( bv_8_92_n253 )  ;
assign n14610 =  ( n14608 ) & (n14609 )  ;
assign n14611 =  ( n14610 ) & (wr )  ;
assign n14612 =  ( n14611 ) ? ( n4782 ) : ( iram_92 ) ;
assign n14613 = wr_addr[7:7] ;
assign n14614 =  ( n14613 ) == ( bv_1_0_n53 )  ;
assign n14615 =  ( wr_addr ) == ( bv_8_92_n253 )  ;
assign n14616 =  ( n14614 ) & (n14615 )  ;
assign n14617 =  ( n14616 ) & (wr )  ;
assign n14618 =  ( n14617 ) ? ( n4841 ) : ( iram_92 ) ;
assign n14619 = wr_addr[7:7] ;
assign n14620 =  ( n14619 ) == ( bv_1_0_n53 )  ;
assign n14621 =  ( wr_addr ) == ( bv_8_92_n253 )  ;
assign n14622 =  ( n14620 ) & (n14621 )  ;
assign n14623 =  ( n14622 ) & (wr )  ;
assign n14624 =  ( n14623 ) ? ( n5449 ) : ( iram_92 ) ;
assign n14625 = wr_addr[7:7] ;
assign n14626 =  ( n14625 ) == ( bv_1_0_n53 )  ;
assign n14627 =  ( wr_addr ) == ( bv_8_92_n253 )  ;
assign n14628 =  ( n14626 ) & (n14627 )  ;
assign n14629 =  ( n14628 ) & (wr )  ;
assign n14630 =  ( n14629 ) ? ( n4906 ) : ( iram_92 ) ;
assign n14631 = wr_addr[7:7] ;
assign n14632 =  ( n14631 ) == ( bv_1_0_n53 )  ;
assign n14633 =  ( wr_addr ) == ( bv_8_92_n253 )  ;
assign n14634 =  ( n14632 ) & (n14633 )  ;
assign n14635 =  ( n14634 ) & (wr )  ;
assign n14636 =  ( n14635 ) ? ( n5485 ) : ( iram_92 ) ;
assign n14637 = wr_addr[7:7] ;
assign n14638 =  ( n14637 ) == ( bv_1_0_n53 )  ;
assign n14639 =  ( wr_addr ) == ( bv_8_92_n253 )  ;
assign n14640 =  ( n14638 ) & (n14639 )  ;
assign n14641 =  ( n14640 ) & (wr )  ;
assign n14642 =  ( n14641 ) ? ( n5512 ) : ( iram_92 ) ;
assign n14643 = wr_addr[7:7] ;
assign n14644 =  ( n14643 ) == ( bv_1_0_n53 )  ;
assign n14645 =  ( wr_addr ) == ( bv_8_92_n253 )  ;
assign n14646 =  ( n14644 ) & (n14645 )  ;
assign n14647 =  ( n14646 ) & (wr )  ;
assign n14648 =  ( n14647 ) ? ( bv_8_0_n69 ) : ( iram_92 ) ;
assign n14649 = wr_addr[7:7] ;
assign n14650 =  ( n14649 ) == ( bv_1_0_n53 )  ;
assign n14651 =  ( wr_addr ) == ( bv_8_92_n253 )  ;
assign n14652 =  ( n14650 ) & (n14651 )  ;
assign n14653 =  ( n14652 ) & (wr )  ;
assign n14654 =  ( n14653 ) ? ( n5071 ) : ( iram_92 ) ;
assign n14655 = wr_addr[7:7] ;
assign n14656 =  ( n14655 ) == ( bv_1_0_n53 )  ;
assign n14657 =  ( wr_addr ) == ( bv_8_92_n253 )  ;
assign n14658 =  ( n14656 ) & (n14657 )  ;
assign n14659 =  ( n14658 ) & (wr )  ;
assign n14660 =  ( n14659 ) ? ( n5096 ) : ( iram_92 ) ;
assign n14661 = wr_addr[7:7] ;
assign n14662 =  ( n14661 ) == ( bv_1_0_n53 )  ;
assign n14663 =  ( wr_addr ) == ( bv_8_92_n253 )  ;
assign n14664 =  ( n14662 ) & (n14663 )  ;
assign n14665 =  ( n14664 ) & (wr )  ;
assign n14666 =  ( n14665 ) ? ( n5123 ) : ( iram_92 ) ;
assign n14667 = wr_addr[7:7] ;
assign n14668 =  ( n14667 ) == ( bv_1_0_n53 )  ;
assign n14669 =  ( wr_addr ) == ( bv_8_92_n253 )  ;
assign n14670 =  ( n14668 ) & (n14669 )  ;
assign n14671 =  ( n14670 ) & (wr )  ;
assign n14672 =  ( n14671 ) ? ( n5165 ) : ( iram_92 ) ;
assign n14673 = wr_addr[7:7] ;
assign n14674 =  ( n14673 ) == ( bv_1_0_n53 )  ;
assign n14675 =  ( wr_addr ) == ( bv_8_92_n253 )  ;
assign n14676 =  ( n14674 ) & (n14675 )  ;
assign n14677 =  ( n14676 ) & (wr )  ;
assign n14678 =  ( n14677 ) ? ( n5204 ) : ( iram_92 ) ;
assign n14679 = wr_addr[7:7] ;
assign n14680 =  ( n14679 ) == ( bv_1_0_n53 )  ;
assign n14681 =  ( wr_addr ) == ( bv_8_92_n253 )  ;
assign n14682 =  ( n14680 ) & (n14681 )  ;
assign n14683 =  ( n14682 ) & (wr )  ;
assign n14684 =  ( n14683 ) ? ( n5262 ) : ( iram_92 ) ;
assign n14685 = wr_addr[7:7] ;
assign n14686 =  ( n14685 ) == ( bv_1_0_n53 )  ;
assign n14687 =  ( wr_addr ) == ( bv_8_92_n253 )  ;
assign n14688 =  ( n14686 ) & (n14687 )  ;
assign n14689 =  ( n14688 ) & (wr )  ;
assign n14690 =  ( n14689 ) ? ( n5298 ) : ( iram_92 ) ;
assign n14691 = wr_addr[7:7] ;
assign n14692 =  ( n14691 ) == ( bv_1_0_n53 )  ;
assign n14693 =  ( wr_addr ) == ( bv_8_92_n253 )  ;
assign n14694 =  ( n14692 ) & (n14693 )  ;
assign n14695 =  ( n14694 ) & (wr )  ;
assign n14696 =  ( n14695 ) ? ( n5325 ) : ( iram_92 ) ;
assign n14697 = wr_addr[7:7] ;
assign n14698 =  ( n14697 ) == ( bv_1_0_n53 )  ;
assign n14699 =  ( wr_addr ) == ( bv_8_93_n255 )  ;
assign n14700 =  ( n14698 ) & (n14699 )  ;
assign n14701 =  ( n14700 ) & (wr )  ;
assign n14702 =  ( n14701 ) ? ( n4782 ) : ( iram_93 ) ;
assign n14703 = wr_addr[7:7] ;
assign n14704 =  ( n14703 ) == ( bv_1_0_n53 )  ;
assign n14705 =  ( wr_addr ) == ( bv_8_93_n255 )  ;
assign n14706 =  ( n14704 ) & (n14705 )  ;
assign n14707 =  ( n14706 ) & (wr )  ;
assign n14708 =  ( n14707 ) ? ( n4841 ) : ( iram_93 ) ;
assign n14709 = wr_addr[7:7] ;
assign n14710 =  ( n14709 ) == ( bv_1_0_n53 )  ;
assign n14711 =  ( wr_addr ) == ( bv_8_93_n255 )  ;
assign n14712 =  ( n14710 ) & (n14711 )  ;
assign n14713 =  ( n14712 ) & (wr )  ;
assign n14714 =  ( n14713 ) ? ( n5449 ) : ( iram_93 ) ;
assign n14715 = wr_addr[7:7] ;
assign n14716 =  ( n14715 ) == ( bv_1_0_n53 )  ;
assign n14717 =  ( wr_addr ) == ( bv_8_93_n255 )  ;
assign n14718 =  ( n14716 ) & (n14717 )  ;
assign n14719 =  ( n14718 ) & (wr )  ;
assign n14720 =  ( n14719 ) ? ( n4906 ) : ( iram_93 ) ;
assign n14721 = wr_addr[7:7] ;
assign n14722 =  ( n14721 ) == ( bv_1_0_n53 )  ;
assign n14723 =  ( wr_addr ) == ( bv_8_93_n255 )  ;
assign n14724 =  ( n14722 ) & (n14723 )  ;
assign n14725 =  ( n14724 ) & (wr )  ;
assign n14726 =  ( n14725 ) ? ( n5485 ) : ( iram_93 ) ;
assign n14727 = wr_addr[7:7] ;
assign n14728 =  ( n14727 ) == ( bv_1_0_n53 )  ;
assign n14729 =  ( wr_addr ) == ( bv_8_93_n255 )  ;
assign n14730 =  ( n14728 ) & (n14729 )  ;
assign n14731 =  ( n14730 ) & (wr )  ;
assign n14732 =  ( n14731 ) ? ( n5512 ) : ( iram_93 ) ;
assign n14733 = wr_addr[7:7] ;
assign n14734 =  ( n14733 ) == ( bv_1_0_n53 )  ;
assign n14735 =  ( wr_addr ) == ( bv_8_93_n255 )  ;
assign n14736 =  ( n14734 ) & (n14735 )  ;
assign n14737 =  ( n14736 ) & (wr )  ;
assign n14738 =  ( n14737 ) ? ( bv_8_0_n69 ) : ( iram_93 ) ;
assign n14739 = wr_addr[7:7] ;
assign n14740 =  ( n14739 ) == ( bv_1_0_n53 )  ;
assign n14741 =  ( wr_addr ) == ( bv_8_93_n255 )  ;
assign n14742 =  ( n14740 ) & (n14741 )  ;
assign n14743 =  ( n14742 ) & (wr )  ;
assign n14744 =  ( n14743 ) ? ( n5071 ) : ( iram_93 ) ;
assign n14745 = wr_addr[7:7] ;
assign n14746 =  ( n14745 ) == ( bv_1_0_n53 )  ;
assign n14747 =  ( wr_addr ) == ( bv_8_93_n255 )  ;
assign n14748 =  ( n14746 ) & (n14747 )  ;
assign n14749 =  ( n14748 ) & (wr )  ;
assign n14750 =  ( n14749 ) ? ( n5096 ) : ( iram_93 ) ;
assign n14751 = wr_addr[7:7] ;
assign n14752 =  ( n14751 ) == ( bv_1_0_n53 )  ;
assign n14753 =  ( wr_addr ) == ( bv_8_93_n255 )  ;
assign n14754 =  ( n14752 ) & (n14753 )  ;
assign n14755 =  ( n14754 ) & (wr )  ;
assign n14756 =  ( n14755 ) ? ( n5123 ) : ( iram_93 ) ;
assign n14757 = wr_addr[7:7] ;
assign n14758 =  ( n14757 ) == ( bv_1_0_n53 )  ;
assign n14759 =  ( wr_addr ) == ( bv_8_93_n255 )  ;
assign n14760 =  ( n14758 ) & (n14759 )  ;
assign n14761 =  ( n14760 ) & (wr )  ;
assign n14762 =  ( n14761 ) ? ( n5165 ) : ( iram_93 ) ;
assign n14763 = wr_addr[7:7] ;
assign n14764 =  ( n14763 ) == ( bv_1_0_n53 )  ;
assign n14765 =  ( wr_addr ) == ( bv_8_93_n255 )  ;
assign n14766 =  ( n14764 ) & (n14765 )  ;
assign n14767 =  ( n14766 ) & (wr )  ;
assign n14768 =  ( n14767 ) ? ( n5204 ) : ( iram_93 ) ;
assign n14769 = wr_addr[7:7] ;
assign n14770 =  ( n14769 ) == ( bv_1_0_n53 )  ;
assign n14771 =  ( wr_addr ) == ( bv_8_93_n255 )  ;
assign n14772 =  ( n14770 ) & (n14771 )  ;
assign n14773 =  ( n14772 ) & (wr )  ;
assign n14774 =  ( n14773 ) ? ( n5262 ) : ( iram_93 ) ;
assign n14775 = wr_addr[7:7] ;
assign n14776 =  ( n14775 ) == ( bv_1_0_n53 )  ;
assign n14777 =  ( wr_addr ) == ( bv_8_93_n255 )  ;
assign n14778 =  ( n14776 ) & (n14777 )  ;
assign n14779 =  ( n14778 ) & (wr )  ;
assign n14780 =  ( n14779 ) ? ( n5298 ) : ( iram_93 ) ;
assign n14781 = wr_addr[7:7] ;
assign n14782 =  ( n14781 ) == ( bv_1_0_n53 )  ;
assign n14783 =  ( wr_addr ) == ( bv_8_93_n255 )  ;
assign n14784 =  ( n14782 ) & (n14783 )  ;
assign n14785 =  ( n14784 ) & (wr )  ;
assign n14786 =  ( n14785 ) ? ( n5325 ) : ( iram_93 ) ;
assign n14787 = wr_addr[7:7] ;
assign n14788 =  ( n14787 ) == ( bv_1_0_n53 )  ;
assign n14789 =  ( wr_addr ) == ( bv_8_94_n257 )  ;
assign n14790 =  ( n14788 ) & (n14789 )  ;
assign n14791 =  ( n14790 ) & (wr )  ;
assign n14792 =  ( n14791 ) ? ( n4782 ) : ( iram_94 ) ;
assign n14793 = wr_addr[7:7] ;
assign n14794 =  ( n14793 ) == ( bv_1_0_n53 )  ;
assign n14795 =  ( wr_addr ) == ( bv_8_94_n257 )  ;
assign n14796 =  ( n14794 ) & (n14795 )  ;
assign n14797 =  ( n14796 ) & (wr )  ;
assign n14798 =  ( n14797 ) ? ( n4841 ) : ( iram_94 ) ;
assign n14799 = wr_addr[7:7] ;
assign n14800 =  ( n14799 ) == ( bv_1_0_n53 )  ;
assign n14801 =  ( wr_addr ) == ( bv_8_94_n257 )  ;
assign n14802 =  ( n14800 ) & (n14801 )  ;
assign n14803 =  ( n14802 ) & (wr )  ;
assign n14804 =  ( n14803 ) ? ( n5449 ) : ( iram_94 ) ;
assign n14805 = wr_addr[7:7] ;
assign n14806 =  ( n14805 ) == ( bv_1_0_n53 )  ;
assign n14807 =  ( wr_addr ) == ( bv_8_94_n257 )  ;
assign n14808 =  ( n14806 ) & (n14807 )  ;
assign n14809 =  ( n14808 ) & (wr )  ;
assign n14810 =  ( n14809 ) ? ( n4906 ) : ( iram_94 ) ;
assign n14811 = wr_addr[7:7] ;
assign n14812 =  ( n14811 ) == ( bv_1_0_n53 )  ;
assign n14813 =  ( wr_addr ) == ( bv_8_94_n257 )  ;
assign n14814 =  ( n14812 ) & (n14813 )  ;
assign n14815 =  ( n14814 ) & (wr )  ;
assign n14816 =  ( n14815 ) ? ( n5485 ) : ( iram_94 ) ;
assign n14817 = wr_addr[7:7] ;
assign n14818 =  ( n14817 ) == ( bv_1_0_n53 )  ;
assign n14819 =  ( wr_addr ) == ( bv_8_94_n257 )  ;
assign n14820 =  ( n14818 ) & (n14819 )  ;
assign n14821 =  ( n14820 ) & (wr )  ;
assign n14822 =  ( n14821 ) ? ( n5512 ) : ( iram_94 ) ;
assign n14823 = wr_addr[7:7] ;
assign n14824 =  ( n14823 ) == ( bv_1_0_n53 )  ;
assign n14825 =  ( wr_addr ) == ( bv_8_94_n257 )  ;
assign n14826 =  ( n14824 ) & (n14825 )  ;
assign n14827 =  ( n14826 ) & (wr )  ;
assign n14828 =  ( n14827 ) ? ( bv_8_0_n69 ) : ( iram_94 ) ;
assign n14829 = wr_addr[7:7] ;
assign n14830 =  ( n14829 ) == ( bv_1_0_n53 )  ;
assign n14831 =  ( wr_addr ) == ( bv_8_94_n257 )  ;
assign n14832 =  ( n14830 ) & (n14831 )  ;
assign n14833 =  ( n14832 ) & (wr )  ;
assign n14834 =  ( n14833 ) ? ( n5071 ) : ( iram_94 ) ;
assign n14835 = wr_addr[7:7] ;
assign n14836 =  ( n14835 ) == ( bv_1_0_n53 )  ;
assign n14837 =  ( wr_addr ) == ( bv_8_94_n257 )  ;
assign n14838 =  ( n14836 ) & (n14837 )  ;
assign n14839 =  ( n14838 ) & (wr )  ;
assign n14840 =  ( n14839 ) ? ( n5096 ) : ( iram_94 ) ;
assign n14841 = wr_addr[7:7] ;
assign n14842 =  ( n14841 ) == ( bv_1_0_n53 )  ;
assign n14843 =  ( wr_addr ) == ( bv_8_94_n257 )  ;
assign n14844 =  ( n14842 ) & (n14843 )  ;
assign n14845 =  ( n14844 ) & (wr )  ;
assign n14846 =  ( n14845 ) ? ( n5123 ) : ( iram_94 ) ;
assign n14847 = wr_addr[7:7] ;
assign n14848 =  ( n14847 ) == ( bv_1_0_n53 )  ;
assign n14849 =  ( wr_addr ) == ( bv_8_94_n257 )  ;
assign n14850 =  ( n14848 ) & (n14849 )  ;
assign n14851 =  ( n14850 ) & (wr )  ;
assign n14852 =  ( n14851 ) ? ( n5165 ) : ( iram_94 ) ;
assign n14853 = wr_addr[7:7] ;
assign n14854 =  ( n14853 ) == ( bv_1_0_n53 )  ;
assign n14855 =  ( wr_addr ) == ( bv_8_94_n257 )  ;
assign n14856 =  ( n14854 ) & (n14855 )  ;
assign n14857 =  ( n14856 ) & (wr )  ;
assign n14858 =  ( n14857 ) ? ( n5204 ) : ( iram_94 ) ;
assign n14859 = wr_addr[7:7] ;
assign n14860 =  ( n14859 ) == ( bv_1_0_n53 )  ;
assign n14861 =  ( wr_addr ) == ( bv_8_94_n257 )  ;
assign n14862 =  ( n14860 ) & (n14861 )  ;
assign n14863 =  ( n14862 ) & (wr )  ;
assign n14864 =  ( n14863 ) ? ( n5262 ) : ( iram_94 ) ;
assign n14865 = wr_addr[7:7] ;
assign n14866 =  ( n14865 ) == ( bv_1_0_n53 )  ;
assign n14867 =  ( wr_addr ) == ( bv_8_94_n257 )  ;
assign n14868 =  ( n14866 ) & (n14867 )  ;
assign n14869 =  ( n14868 ) & (wr )  ;
assign n14870 =  ( n14869 ) ? ( n5298 ) : ( iram_94 ) ;
assign n14871 = wr_addr[7:7] ;
assign n14872 =  ( n14871 ) == ( bv_1_0_n53 )  ;
assign n14873 =  ( wr_addr ) == ( bv_8_94_n257 )  ;
assign n14874 =  ( n14872 ) & (n14873 )  ;
assign n14875 =  ( n14874 ) & (wr )  ;
assign n14876 =  ( n14875 ) ? ( n5325 ) : ( iram_94 ) ;
assign n14877 = wr_addr[7:7] ;
assign n14878 =  ( n14877 ) == ( bv_1_0_n53 )  ;
assign n14879 =  ( wr_addr ) == ( bv_8_95_n259 )  ;
assign n14880 =  ( n14878 ) & (n14879 )  ;
assign n14881 =  ( n14880 ) & (wr )  ;
assign n14882 =  ( n14881 ) ? ( n4782 ) : ( iram_95 ) ;
assign n14883 = wr_addr[7:7] ;
assign n14884 =  ( n14883 ) == ( bv_1_0_n53 )  ;
assign n14885 =  ( wr_addr ) == ( bv_8_95_n259 )  ;
assign n14886 =  ( n14884 ) & (n14885 )  ;
assign n14887 =  ( n14886 ) & (wr )  ;
assign n14888 =  ( n14887 ) ? ( n4841 ) : ( iram_95 ) ;
assign n14889 = wr_addr[7:7] ;
assign n14890 =  ( n14889 ) == ( bv_1_0_n53 )  ;
assign n14891 =  ( wr_addr ) == ( bv_8_95_n259 )  ;
assign n14892 =  ( n14890 ) & (n14891 )  ;
assign n14893 =  ( n14892 ) & (wr )  ;
assign n14894 =  ( n14893 ) ? ( n5449 ) : ( iram_95 ) ;
assign n14895 = wr_addr[7:7] ;
assign n14896 =  ( n14895 ) == ( bv_1_0_n53 )  ;
assign n14897 =  ( wr_addr ) == ( bv_8_95_n259 )  ;
assign n14898 =  ( n14896 ) & (n14897 )  ;
assign n14899 =  ( n14898 ) & (wr )  ;
assign n14900 =  ( n14899 ) ? ( n4906 ) : ( iram_95 ) ;
assign n14901 = wr_addr[7:7] ;
assign n14902 =  ( n14901 ) == ( bv_1_0_n53 )  ;
assign n14903 =  ( wr_addr ) == ( bv_8_95_n259 )  ;
assign n14904 =  ( n14902 ) & (n14903 )  ;
assign n14905 =  ( n14904 ) & (wr )  ;
assign n14906 =  ( n14905 ) ? ( n5485 ) : ( iram_95 ) ;
assign n14907 = wr_addr[7:7] ;
assign n14908 =  ( n14907 ) == ( bv_1_0_n53 )  ;
assign n14909 =  ( wr_addr ) == ( bv_8_95_n259 )  ;
assign n14910 =  ( n14908 ) & (n14909 )  ;
assign n14911 =  ( n14910 ) & (wr )  ;
assign n14912 =  ( n14911 ) ? ( n5512 ) : ( iram_95 ) ;
assign n14913 = wr_addr[7:7] ;
assign n14914 =  ( n14913 ) == ( bv_1_0_n53 )  ;
assign n14915 =  ( wr_addr ) == ( bv_8_95_n259 )  ;
assign n14916 =  ( n14914 ) & (n14915 )  ;
assign n14917 =  ( n14916 ) & (wr )  ;
assign n14918 =  ( n14917 ) ? ( bv_8_0_n69 ) : ( iram_95 ) ;
assign n14919 = wr_addr[7:7] ;
assign n14920 =  ( n14919 ) == ( bv_1_0_n53 )  ;
assign n14921 =  ( wr_addr ) == ( bv_8_95_n259 )  ;
assign n14922 =  ( n14920 ) & (n14921 )  ;
assign n14923 =  ( n14922 ) & (wr )  ;
assign n14924 =  ( n14923 ) ? ( n5071 ) : ( iram_95 ) ;
assign n14925 = wr_addr[7:7] ;
assign n14926 =  ( n14925 ) == ( bv_1_0_n53 )  ;
assign n14927 =  ( wr_addr ) == ( bv_8_95_n259 )  ;
assign n14928 =  ( n14926 ) & (n14927 )  ;
assign n14929 =  ( n14928 ) & (wr )  ;
assign n14930 =  ( n14929 ) ? ( n5096 ) : ( iram_95 ) ;
assign n14931 = wr_addr[7:7] ;
assign n14932 =  ( n14931 ) == ( bv_1_0_n53 )  ;
assign n14933 =  ( wr_addr ) == ( bv_8_95_n259 )  ;
assign n14934 =  ( n14932 ) & (n14933 )  ;
assign n14935 =  ( n14934 ) & (wr )  ;
assign n14936 =  ( n14935 ) ? ( n5123 ) : ( iram_95 ) ;
assign n14937 = wr_addr[7:7] ;
assign n14938 =  ( n14937 ) == ( bv_1_0_n53 )  ;
assign n14939 =  ( wr_addr ) == ( bv_8_95_n259 )  ;
assign n14940 =  ( n14938 ) & (n14939 )  ;
assign n14941 =  ( n14940 ) & (wr )  ;
assign n14942 =  ( n14941 ) ? ( n5165 ) : ( iram_95 ) ;
assign n14943 = wr_addr[7:7] ;
assign n14944 =  ( n14943 ) == ( bv_1_0_n53 )  ;
assign n14945 =  ( wr_addr ) == ( bv_8_95_n259 )  ;
assign n14946 =  ( n14944 ) & (n14945 )  ;
assign n14947 =  ( n14946 ) & (wr )  ;
assign n14948 =  ( n14947 ) ? ( n5204 ) : ( iram_95 ) ;
assign n14949 = wr_addr[7:7] ;
assign n14950 =  ( n14949 ) == ( bv_1_0_n53 )  ;
assign n14951 =  ( wr_addr ) == ( bv_8_95_n259 )  ;
assign n14952 =  ( n14950 ) & (n14951 )  ;
assign n14953 =  ( n14952 ) & (wr )  ;
assign n14954 =  ( n14953 ) ? ( n5262 ) : ( iram_95 ) ;
assign n14955 = wr_addr[7:7] ;
assign n14956 =  ( n14955 ) == ( bv_1_0_n53 )  ;
assign n14957 =  ( wr_addr ) == ( bv_8_95_n259 )  ;
assign n14958 =  ( n14956 ) & (n14957 )  ;
assign n14959 =  ( n14958 ) & (wr )  ;
assign n14960 =  ( n14959 ) ? ( n5298 ) : ( iram_95 ) ;
assign n14961 = wr_addr[7:7] ;
assign n14962 =  ( n14961 ) == ( bv_1_0_n53 )  ;
assign n14963 =  ( wr_addr ) == ( bv_8_95_n259 )  ;
assign n14964 =  ( n14962 ) & (n14963 )  ;
assign n14965 =  ( n14964 ) & (wr )  ;
assign n14966 =  ( n14965 ) ? ( n5325 ) : ( iram_95 ) ;
assign n14967 = wr_addr[7:7] ;
assign n14968 =  ( n14967 ) == ( bv_1_0_n53 )  ;
assign n14969 =  ( wr_addr ) == ( bv_8_96_n261 )  ;
assign n14970 =  ( n14968 ) & (n14969 )  ;
assign n14971 =  ( n14970 ) & (wr )  ;
assign n14972 =  ( n14971 ) ? ( n4782 ) : ( iram_96 ) ;
assign n14973 = wr_addr[7:7] ;
assign n14974 =  ( n14973 ) == ( bv_1_0_n53 )  ;
assign n14975 =  ( wr_addr ) == ( bv_8_96_n261 )  ;
assign n14976 =  ( n14974 ) & (n14975 )  ;
assign n14977 =  ( n14976 ) & (wr )  ;
assign n14978 =  ( n14977 ) ? ( n4841 ) : ( iram_96 ) ;
assign n14979 = wr_addr[7:7] ;
assign n14980 =  ( n14979 ) == ( bv_1_0_n53 )  ;
assign n14981 =  ( wr_addr ) == ( bv_8_96_n261 )  ;
assign n14982 =  ( n14980 ) & (n14981 )  ;
assign n14983 =  ( n14982 ) & (wr )  ;
assign n14984 =  ( n14983 ) ? ( n5449 ) : ( iram_96 ) ;
assign n14985 = wr_addr[7:7] ;
assign n14986 =  ( n14985 ) == ( bv_1_0_n53 )  ;
assign n14987 =  ( wr_addr ) == ( bv_8_96_n261 )  ;
assign n14988 =  ( n14986 ) & (n14987 )  ;
assign n14989 =  ( n14988 ) & (wr )  ;
assign n14990 =  ( n14989 ) ? ( n4906 ) : ( iram_96 ) ;
assign n14991 = wr_addr[7:7] ;
assign n14992 =  ( n14991 ) == ( bv_1_0_n53 )  ;
assign n14993 =  ( wr_addr ) == ( bv_8_96_n261 )  ;
assign n14994 =  ( n14992 ) & (n14993 )  ;
assign n14995 =  ( n14994 ) & (wr )  ;
assign n14996 =  ( n14995 ) ? ( n5485 ) : ( iram_96 ) ;
assign n14997 = wr_addr[7:7] ;
assign n14998 =  ( n14997 ) == ( bv_1_0_n53 )  ;
assign n14999 =  ( wr_addr ) == ( bv_8_96_n261 )  ;
assign n15000 =  ( n14998 ) & (n14999 )  ;
assign n15001 =  ( n15000 ) & (wr )  ;
assign n15002 =  ( n15001 ) ? ( n5512 ) : ( iram_96 ) ;
assign n15003 = wr_addr[7:7] ;
assign n15004 =  ( n15003 ) == ( bv_1_0_n53 )  ;
assign n15005 =  ( wr_addr ) == ( bv_8_96_n261 )  ;
assign n15006 =  ( n15004 ) & (n15005 )  ;
assign n15007 =  ( n15006 ) & (wr )  ;
assign n15008 =  ( n15007 ) ? ( bv_8_0_n69 ) : ( iram_96 ) ;
assign n15009 = wr_addr[7:7] ;
assign n15010 =  ( n15009 ) == ( bv_1_0_n53 )  ;
assign n15011 =  ( wr_addr ) == ( bv_8_96_n261 )  ;
assign n15012 =  ( n15010 ) & (n15011 )  ;
assign n15013 =  ( n15012 ) & (wr )  ;
assign n15014 =  ( n15013 ) ? ( n5071 ) : ( iram_96 ) ;
assign n15015 = wr_addr[7:7] ;
assign n15016 =  ( n15015 ) == ( bv_1_0_n53 )  ;
assign n15017 =  ( wr_addr ) == ( bv_8_96_n261 )  ;
assign n15018 =  ( n15016 ) & (n15017 )  ;
assign n15019 =  ( n15018 ) & (wr )  ;
assign n15020 =  ( n15019 ) ? ( n5096 ) : ( iram_96 ) ;
assign n15021 = wr_addr[7:7] ;
assign n15022 =  ( n15021 ) == ( bv_1_0_n53 )  ;
assign n15023 =  ( wr_addr ) == ( bv_8_96_n261 )  ;
assign n15024 =  ( n15022 ) & (n15023 )  ;
assign n15025 =  ( n15024 ) & (wr )  ;
assign n15026 =  ( n15025 ) ? ( n5123 ) : ( iram_96 ) ;
assign n15027 = wr_addr[7:7] ;
assign n15028 =  ( n15027 ) == ( bv_1_0_n53 )  ;
assign n15029 =  ( wr_addr ) == ( bv_8_96_n261 )  ;
assign n15030 =  ( n15028 ) & (n15029 )  ;
assign n15031 =  ( n15030 ) & (wr )  ;
assign n15032 =  ( n15031 ) ? ( n5165 ) : ( iram_96 ) ;
assign n15033 = wr_addr[7:7] ;
assign n15034 =  ( n15033 ) == ( bv_1_0_n53 )  ;
assign n15035 =  ( wr_addr ) == ( bv_8_96_n261 )  ;
assign n15036 =  ( n15034 ) & (n15035 )  ;
assign n15037 =  ( n15036 ) & (wr )  ;
assign n15038 =  ( n15037 ) ? ( n5204 ) : ( iram_96 ) ;
assign n15039 = wr_addr[7:7] ;
assign n15040 =  ( n15039 ) == ( bv_1_0_n53 )  ;
assign n15041 =  ( wr_addr ) == ( bv_8_96_n261 )  ;
assign n15042 =  ( n15040 ) & (n15041 )  ;
assign n15043 =  ( n15042 ) & (wr )  ;
assign n15044 =  ( n15043 ) ? ( n5262 ) : ( iram_96 ) ;
assign n15045 = wr_addr[7:7] ;
assign n15046 =  ( n15045 ) == ( bv_1_0_n53 )  ;
assign n15047 =  ( wr_addr ) == ( bv_8_96_n261 )  ;
assign n15048 =  ( n15046 ) & (n15047 )  ;
assign n15049 =  ( n15048 ) & (wr )  ;
assign n15050 =  ( n15049 ) ? ( n5298 ) : ( iram_96 ) ;
assign n15051 = wr_addr[7:7] ;
assign n15052 =  ( n15051 ) == ( bv_1_0_n53 )  ;
assign n15053 =  ( wr_addr ) == ( bv_8_96_n261 )  ;
assign n15054 =  ( n15052 ) & (n15053 )  ;
assign n15055 =  ( n15054 ) & (wr )  ;
assign n15056 =  ( n15055 ) ? ( n5325 ) : ( iram_96 ) ;
assign n15057 = wr_addr[7:7] ;
assign n15058 =  ( n15057 ) == ( bv_1_0_n53 )  ;
assign n15059 =  ( wr_addr ) == ( bv_8_97_n263 )  ;
assign n15060 =  ( n15058 ) & (n15059 )  ;
assign n15061 =  ( n15060 ) & (wr )  ;
assign n15062 =  ( n15061 ) ? ( n4782 ) : ( iram_97 ) ;
assign n15063 = wr_addr[7:7] ;
assign n15064 =  ( n15063 ) == ( bv_1_0_n53 )  ;
assign n15065 =  ( wr_addr ) == ( bv_8_97_n263 )  ;
assign n15066 =  ( n15064 ) & (n15065 )  ;
assign n15067 =  ( n15066 ) & (wr )  ;
assign n15068 =  ( n15067 ) ? ( n4841 ) : ( iram_97 ) ;
assign n15069 = wr_addr[7:7] ;
assign n15070 =  ( n15069 ) == ( bv_1_0_n53 )  ;
assign n15071 =  ( wr_addr ) == ( bv_8_97_n263 )  ;
assign n15072 =  ( n15070 ) & (n15071 )  ;
assign n15073 =  ( n15072 ) & (wr )  ;
assign n15074 =  ( n15073 ) ? ( n5449 ) : ( iram_97 ) ;
assign n15075 = wr_addr[7:7] ;
assign n15076 =  ( n15075 ) == ( bv_1_0_n53 )  ;
assign n15077 =  ( wr_addr ) == ( bv_8_97_n263 )  ;
assign n15078 =  ( n15076 ) & (n15077 )  ;
assign n15079 =  ( n15078 ) & (wr )  ;
assign n15080 =  ( n15079 ) ? ( n4906 ) : ( iram_97 ) ;
assign n15081 = wr_addr[7:7] ;
assign n15082 =  ( n15081 ) == ( bv_1_0_n53 )  ;
assign n15083 =  ( wr_addr ) == ( bv_8_97_n263 )  ;
assign n15084 =  ( n15082 ) & (n15083 )  ;
assign n15085 =  ( n15084 ) & (wr )  ;
assign n15086 =  ( n15085 ) ? ( n5485 ) : ( iram_97 ) ;
assign n15087 = wr_addr[7:7] ;
assign n15088 =  ( n15087 ) == ( bv_1_0_n53 )  ;
assign n15089 =  ( wr_addr ) == ( bv_8_97_n263 )  ;
assign n15090 =  ( n15088 ) & (n15089 )  ;
assign n15091 =  ( n15090 ) & (wr )  ;
assign n15092 =  ( n15091 ) ? ( n5512 ) : ( iram_97 ) ;
assign n15093 = wr_addr[7:7] ;
assign n15094 =  ( n15093 ) == ( bv_1_0_n53 )  ;
assign n15095 =  ( wr_addr ) == ( bv_8_97_n263 )  ;
assign n15096 =  ( n15094 ) & (n15095 )  ;
assign n15097 =  ( n15096 ) & (wr )  ;
assign n15098 =  ( n15097 ) ? ( bv_8_0_n69 ) : ( iram_97 ) ;
assign n15099 = wr_addr[7:7] ;
assign n15100 =  ( n15099 ) == ( bv_1_0_n53 )  ;
assign n15101 =  ( wr_addr ) == ( bv_8_97_n263 )  ;
assign n15102 =  ( n15100 ) & (n15101 )  ;
assign n15103 =  ( n15102 ) & (wr )  ;
assign n15104 =  ( n15103 ) ? ( n5071 ) : ( iram_97 ) ;
assign n15105 = wr_addr[7:7] ;
assign n15106 =  ( n15105 ) == ( bv_1_0_n53 )  ;
assign n15107 =  ( wr_addr ) == ( bv_8_97_n263 )  ;
assign n15108 =  ( n15106 ) & (n15107 )  ;
assign n15109 =  ( n15108 ) & (wr )  ;
assign n15110 =  ( n15109 ) ? ( n5096 ) : ( iram_97 ) ;
assign n15111 = wr_addr[7:7] ;
assign n15112 =  ( n15111 ) == ( bv_1_0_n53 )  ;
assign n15113 =  ( wr_addr ) == ( bv_8_97_n263 )  ;
assign n15114 =  ( n15112 ) & (n15113 )  ;
assign n15115 =  ( n15114 ) & (wr )  ;
assign n15116 =  ( n15115 ) ? ( n5123 ) : ( iram_97 ) ;
assign n15117 = wr_addr[7:7] ;
assign n15118 =  ( n15117 ) == ( bv_1_0_n53 )  ;
assign n15119 =  ( wr_addr ) == ( bv_8_97_n263 )  ;
assign n15120 =  ( n15118 ) & (n15119 )  ;
assign n15121 =  ( n15120 ) & (wr )  ;
assign n15122 =  ( n15121 ) ? ( n5165 ) : ( iram_97 ) ;
assign n15123 = wr_addr[7:7] ;
assign n15124 =  ( n15123 ) == ( bv_1_0_n53 )  ;
assign n15125 =  ( wr_addr ) == ( bv_8_97_n263 )  ;
assign n15126 =  ( n15124 ) & (n15125 )  ;
assign n15127 =  ( n15126 ) & (wr )  ;
assign n15128 =  ( n15127 ) ? ( n5204 ) : ( iram_97 ) ;
assign n15129 = wr_addr[7:7] ;
assign n15130 =  ( n15129 ) == ( bv_1_0_n53 )  ;
assign n15131 =  ( wr_addr ) == ( bv_8_97_n263 )  ;
assign n15132 =  ( n15130 ) & (n15131 )  ;
assign n15133 =  ( n15132 ) & (wr )  ;
assign n15134 =  ( n15133 ) ? ( n5262 ) : ( iram_97 ) ;
assign n15135 = wr_addr[7:7] ;
assign n15136 =  ( n15135 ) == ( bv_1_0_n53 )  ;
assign n15137 =  ( wr_addr ) == ( bv_8_97_n263 )  ;
assign n15138 =  ( n15136 ) & (n15137 )  ;
assign n15139 =  ( n15138 ) & (wr )  ;
assign n15140 =  ( n15139 ) ? ( n5298 ) : ( iram_97 ) ;
assign n15141 = wr_addr[7:7] ;
assign n15142 =  ( n15141 ) == ( bv_1_0_n53 )  ;
assign n15143 =  ( wr_addr ) == ( bv_8_97_n263 )  ;
assign n15144 =  ( n15142 ) & (n15143 )  ;
assign n15145 =  ( n15144 ) & (wr )  ;
assign n15146 =  ( n15145 ) ? ( n5325 ) : ( iram_97 ) ;
assign n15147 = wr_addr[7:7] ;
assign n15148 =  ( n15147 ) == ( bv_1_0_n53 )  ;
assign n15149 =  ( wr_addr ) == ( bv_8_98_n265 )  ;
assign n15150 =  ( n15148 ) & (n15149 )  ;
assign n15151 =  ( n15150 ) & (wr )  ;
assign n15152 =  ( n15151 ) ? ( n4782 ) : ( iram_98 ) ;
assign n15153 = wr_addr[7:7] ;
assign n15154 =  ( n15153 ) == ( bv_1_0_n53 )  ;
assign n15155 =  ( wr_addr ) == ( bv_8_98_n265 )  ;
assign n15156 =  ( n15154 ) & (n15155 )  ;
assign n15157 =  ( n15156 ) & (wr )  ;
assign n15158 =  ( n15157 ) ? ( n4841 ) : ( iram_98 ) ;
assign n15159 = wr_addr[7:7] ;
assign n15160 =  ( n15159 ) == ( bv_1_0_n53 )  ;
assign n15161 =  ( wr_addr ) == ( bv_8_98_n265 )  ;
assign n15162 =  ( n15160 ) & (n15161 )  ;
assign n15163 =  ( n15162 ) & (wr )  ;
assign n15164 =  ( n15163 ) ? ( n5449 ) : ( iram_98 ) ;
assign n15165 = wr_addr[7:7] ;
assign n15166 =  ( n15165 ) == ( bv_1_0_n53 )  ;
assign n15167 =  ( wr_addr ) == ( bv_8_98_n265 )  ;
assign n15168 =  ( n15166 ) & (n15167 )  ;
assign n15169 =  ( n15168 ) & (wr )  ;
assign n15170 =  ( n15169 ) ? ( n4906 ) : ( iram_98 ) ;
assign n15171 = wr_addr[7:7] ;
assign n15172 =  ( n15171 ) == ( bv_1_0_n53 )  ;
assign n15173 =  ( wr_addr ) == ( bv_8_98_n265 )  ;
assign n15174 =  ( n15172 ) & (n15173 )  ;
assign n15175 =  ( n15174 ) & (wr )  ;
assign n15176 =  ( n15175 ) ? ( n5485 ) : ( iram_98 ) ;
assign n15177 = wr_addr[7:7] ;
assign n15178 =  ( n15177 ) == ( bv_1_0_n53 )  ;
assign n15179 =  ( wr_addr ) == ( bv_8_98_n265 )  ;
assign n15180 =  ( n15178 ) & (n15179 )  ;
assign n15181 =  ( n15180 ) & (wr )  ;
assign n15182 =  ( n15181 ) ? ( n5512 ) : ( iram_98 ) ;
assign n15183 = wr_addr[7:7] ;
assign n15184 =  ( n15183 ) == ( bv_1_0_n53 )  ;
assign n15185 =  ( wr_addr ) == ( bv_8_98_n265 )  ;
assign n15186 =  ( n15184 ) & (n15185 )  ;
assign n15187 =  ( n15186 ) & (wr )  ;
assign n15188 =  ( n15187 ) ? ( bv_8_0_n69 ) : ( iram_98 ) ;
assign n15189 = wr_addr[7:7] ;
assign n15190 =  ( n15189 ) == ( bv_1_0_n53 )  ;
assign n15191 =  ( wr_addr ) == ( bv_8_98_n265 )  ;
assign n15192 =  ( n15190 ) & (n15191 )  ;
assign n15193 =  ( n15192 ) & (wr )  ;
assign n15194 =  ( n15193 ) ? ( n5071 ) : ( iram_98 ) ;
assign n15195 = wr_addr[7:7] ;
assign n15196 =  ( n15195 ) == ( bv_1_0_n53 )  ;
assign n15197 =  ( wr_addr ) == ( bv_8_98_n265 )  ;
assign n15198 =  ( n15196 ) & (n15197 )  ;
assign n15199 =  ( n15198 ) & (wr )  ;
assign n15200 =  ( n15199 ) ? ( n5096 ) : ( iram_98 ) ;
assign n15201 = wr_addr[7:7] ;
assign n15202 =  ( n15201 ) == ( bv_1_0_n53 )  ;
assign n15203 =  ( wr_addr ) == ( bv_8_98_n265 )  ;
assign n15204 =  ( n15202 ) & (n15203 )  ;
assign n15205 =  ( n15204 ) & (wr )  ;
assign n15206 =  ( n15205 ) ? ( n5123 ) : ( iram_98 ) ;
assign n15207 = wr_addr[7:7] ;
assign n15208 =  ( n15207 ) == ( bv_1_0_n53 )  ;
assign n15209 =  ( wr_addr ) == ( bv_8_98_n265 )  ;
assign n15210 =  ( n15208 ) & (n15209 )  ;
assign n15211 =  ( n15210 ) & (wr )  ;
assign n15212 =  ( n15211 ) ? ( n5165 ) : ( iram_98 ) ;
assign n15213 = wr_addr[7:7] ;
assign n15214 =  ( n15213 ) == ( bv_1_0_n53 )  ;
assign n15215 =  ( wr_addr ) == ( bv_8_98_n265 )  ;
assign n15216 =  ( n15214 ) & (n15215 )  ;
assign n15217 =  ( n15216 ) & (wr )  ;
assign n15218 =  ( n15217 ) ? ( n5204 ) : ( iram_98 ) ;
assign n15219 = wr_addr[7:7] ;
assign n15220 =  ( n15219 ) == ( bv_1_0_n53 )  ;
assign n15221 =  ( wr_addr ) == ( bv_8_98_n265 )  ;
assign n15222 =  ( n15220 ) & (n15221 )  ;
assign n15223 =  ( n15222 ) & (wr )  ;
assign n15224 =  ( n15223 ) ? ( n5262 ) : ( iram_98 ) ;
assign n15225 = wr_addr[7:7] ;
assign n15226 =  ( n15225 ) == ( bv_1_0_n53 )  ;
assign n15227 =  ( wr_addr ) == ( bv_8_98_n265 )  ;
assign n15228 =  ( n15226 ) & (n15227 )  ;
assign n15229 =  ( n15228 ) & (wr )  ;
assign n15230 =  ( n15229 ) ? ( n5298 ) : ( iram_98 ) ;
assign n15231 = wr_addr[7:7] ;
assign n15232 =  ( n15231 ) == ( bv_1_0_n53 )  ;
assign n15233 =  ( wr_addr ) == ( bv_8_98_n265 )  ;
assign n15234 =  ( n15232 ) & (n15233 )  ;
assign n15235 =  ( n15234 ) & (wr )  ;
assign n15236 =  ( n15235 ) ? ( n5325 ) : ( iram_98 ) ;
assign n15237 = wr_addr[7:7] ;
assign n15238 =  ( n15237 ) == ( bv_1_0_n53 )  ;
assign n15239 =  ( wr_addr ) == ( bv_8_99_n267 )  ;
assign n15240 =  ( n15238 ) & (n15239 )  ;
assign n15241 =  ( n15240 ) & (wr )  ;
assign n15242 =  ( n15241 ) ? ( n4782 ) : ( iram_99 ) ;
assign n15243 = wr_addr[7:7] ;
assign n15244 =  ( n15243 ) == ( bv_1_0_n53 )  ;
assign n15245 =  ( wr_addr ) == ( bv_8_99_n267 )  ;
assign n15246 =  ( n15244 ) & (n15245 )  ;
assign n15247 =  ( n15246 ) & (wr )  ;
assign n15248 =  ( n15247 ) ? ( n4841 ) : ( iram_99 ) ;
assign n15249 = wr_addr[7:7] ;
assign n15250 =  ( n15249 ) == ( bv_1_0_n53 )  ;
assign n15251 =  ( wr_addr ) == ( bv_8_99_n267 )  ;
assign n15252 =  ( n15250 ) & (n15251 )  ;
assign n15253 =  ( n15252 ) & (wr )  ;
assign n15254 =  ( n15253 ) ? ( n5449 ) : ( iram_99 ) ;
assign n15255 = wr_addr[7:7] ;
assign n15256 =  ( n15255 ) == ( bv_1_0_n53 )  ;
assign n15257 =  ( wr_addr ) == ( bv_8_99_n267 )  ;
assign n15258 =  ( n15256 ) & (n15257 )  ;
assign n15259 =  ( n15258 ) & (wr )  ;
assign n15260 =  ( n15259 ) ? ( n4906 ) : ( iram_99 ) ;
assign n15261 = wr_addr[7:7] ;
assign n15262 =  ( n15261 ) == ( bv_1_0_n53 )  ;
assign n15263 =  ( wr_addr ) == ( bv_8_99_n267 )  ;
assign n15264 =  ( n15262 ) & (n15263 )  ;
assign n15265 =  ( n15264 ) & (wr )  ;
assign n15266 =  ( n15265 ) ? ( n5485 ) : ( iram_99 ) ;
assign n15267 = wr_addr[7:7] ;
assign n15268 =  ( n15267 ) == ( bv_1_0_n53 )  ;
assign n15269 =  ( wr_addr ) == ( bv_8_99_n267 )  ;
assign n15270 =  ( n15268 ) & (n15269 )  ;
assign n15271 =  ( n15270 ) & (wr )  ;
assign n15272 =  ( n15271 ) ? ( n5512 ) : ( iram_99 ) ;
assign n15273 = wr_addr[7:7] ;
assign n15274 =  ( n15273 ) == ( bv_1_0_n53 )  ;
assign n15275 =  ( wr_addr ) == ( bv_8_99_n267 )  ;
assign n15276 =  ( n15274 ) & (n15275 )  ;
assign n15277 =  ( n15276 ) & (wr )  ;
assign n15278 =  ( n15277 ) ? ( bv_8_0_n69 ) : ( iram_99 ) ;
assign n15279 = wr_addr[7:7] ;
assign n15280 =  ( n15279 ) == ( bv_1_0_n53 )  ;
assign n15281 =  ( wr_addr ) == ( bv_8_99_n267 )  ;
assign n15282 =  ( n15280 ) & (n15281 )  ;
assign n15283 =  ( n15282 ) & (wr )  ;
assign n15284 =  ( n15283 ) ? ( n5071 ) : ( iram_99 ) ;
assign n15285 = wr_addr[7:7] ;
assign n15286 =  ( n15285 ) == ( bv_1_0_n53 )  ;
assign n15287 =  ( wr_addr ) == ( bv_8_99_n267 )  ;
assign n15288 =  ( n15286 ) & (n15287 )  ;
assign n15289 =  ( n15288 ) & (wr )  ;
assign n15290 =  ( n15289 ) ? ( n5096 ) : ( iram_99 ) ;
assign n15291 = wr_addr[7:7] ;
assign n15292 =  ( n15291 ) == ( bv_1_0_n53 )  ;
assign n15293 =  ( wr_addr ) == ( bv_8_99_n267 )  ;
assign n15294 =  ( n15292 ) & (n15293 )  ;
assign n15295 =  ( n15294 ) & (wr )  ;
assign n15296 =  ( n15295 ) ? ( n5123 ) : ( iram_99 ) ;
assign n15297 = wr_addr[7:7] ;
assign n15298 =  ( n15297 ) == ( bv_1_0_n53 )  ;
assign n15299 =  ( wr_addr ) == ( bv_8_99_n267 )  ;
assign n15300 =  ( n15298 ) & (n15299 )  ;
assign n15301 =  ( n15300 ) & (wr )  ;
assign n15302 =  ( n15301 ) ? ( n5165 ) : ( iram_99 ) ;
assign n15303 = wr_addr[7:7] ;
assign n15304 =  ( n15303 ) == ( bv_1_0_n53 )  ;
assign n15305 =  ( wr_addr ) == ( bv_8_99_n267 )  ;
assign n15306 =  ( n15304 ) & (n15305 )  ;
assign n15307 =  ( n15306 ) & (wr )  ;
assign n15308 =  ( n15307 ) ? ( n5204 ) : ( iram_99 ) ;
assign n15309 = wr_addr[7:7] ;
assign n15310 =  ( n15309 ) == ( bv_1_0_n53 )  ;
assign n15311 =  ( wr_addr ) == ( bv_8_99_n267 )  ;
assign n15312 =  ( n15310 ) & (n15311 )  ;
assign n15313 =  ( n15312 ) & (wr )  ;
assign n15314 =  ( n15313 ) ? ( n5262 ) : ( iram_99 ) ;
assign n15315 = wr_addr[7:7] ;
assign n15316 =  ( n15315 ) == ( bv_1_0_n53 )  ;
assign n15317 =  ( wr_addr ) == ( bv_8_99_n267 )  ;
assign n15318 =  ( n15316 ) & (n15317 )  ;
assign n15319 =  ( n15318 ) & (wr )  ;
assign n15320 =  ( n15319 ) ? ( n5298 ) : ( iram_99 ) ;
assign n15321 = wr_addr[7:7] ;
assign n15322 =  ( n15321 ) == ( bv_1_0_n53 )  ;
assign n15323 =  ( wr_addr ) == ( bv_8_99_n267 )  ;
assign n15324 =  ( n15322 ) & (n15323 )  ;
assign n15325 =  ( n15324 ) & (wr )  ;
assign n15326 =  ( n15325 ) ? ( n5325 ) : ( iram_99 ) ;
assign n15327 = wr_addr[7:7] ;
assign n15328 =  ( n15327 ) == ( bv_1_0_n53 )  ;
assign n15329 =  ( wr_addr ) == ( bv_8_100_n269 )  ;
assign n15330 =  ( n15328 ) & (n15329 )  ;
assign n15331 =  ( n15330 ) & (wr )  ;
assign n15332 =  ( n15331 ) ? ( n4782 ) : ( iram_100 ) ;
assign n15333 = wr_addr[7:7] ;
assign n15334 =  ( n15333 ) == ( bv_1_0_n53 )  ;
assign n15335 =  ( wr_addr ) == ( bv_8_100_n269 )  ;
assign n15336 =  ( n15334 ) & (n15335 )  ;
assign n15337 =  ( n15336 ) & (wr )  ;
assign n15338 =  ( n15337 ) ? ( n4841 ) : ( iram_100 ) ;
assign n15339 = wr_addr[7:7] ;
assign n15340 =  ( n15339 ) == ( bv_1_0_n53 )  ;
assign n15341 =  ( wr_addr ) == ( bv_8_100_n269 )  ;
assign n15342 =  ( n15340 ) & (n15341 )  ;
assign n15343 =  ( n15342 ) & (wr )  ;
assign n15344 =  ( n15343 ) ? ( n5449 ) : ( iram_100 ) ;
assign n15345 = wr_addr[7:7] ;
assign n15346 =  ( n15345 ) == ( bv_1_0_n53 )  ;
assign n15347 =  ( wr_addr ) == ( bv_8_100_n269 )  ;
assign n15348 =  ( n15346 ) & (n15347 )  ;
assign n15349 =  ( n15348 ) & (wr )  ;
assign n15350 =  ( n15349 ) ? ( n4906 ) : ( iram_100 ) ;
assign n15351 = wr_addr[7:7] ;
assign n15352 =  ( n15351 ) == ( bv_1_0_n53 )  ;
assign n15353 =  ( wr_addr ) == ( bv_8_100_n269 )  ;
assign n15354 =  ( n15352 ) & (n15353 )  ;
assign n15355 =  ( n15354 ) & (wr )  ;
assign n15356 =  ( n15355 ) ? ( n5485 ) : ( iram_100 ) ;
assign n15357 = wr_addr[7:7] ;
assign n15358 =  ( n15357 ) == ( bv_1_0_n53 )  ;
assign n15359 =  ( wr_addr ) == ( bv_8_100_n269 )  ;
assign n15360 =  ( n15358 ) & (n15359 )  ;
assign n15361 =  ( n15360 ) & (wr )  ;
assign n15362 =  ( n15361 ) ? ( n5512 ) : ( iram_100 ) ;
assign n15363 = wr_addr[7:7] ;
assign n15364 =  ( n15363 ) == ( bv_1_0_n53 )  ;
assign n15365 =  ( wr_addr ) == ( bv_8_100_n269 )  ;
assign n15366 =  ( n15364 ) & (n15365 )  ;
assign n15367 =  ( n15366 ) & (wr )  ;
assign n15368 =  ( n15367 ) ? ( bv_8_0_n69 ) : ( iram_100 ) ;
assign n15369 = wr_addr[7:7] ;
assign n15370 =  ( n15369 ) == ( bv_1_0_n53 )  ;
assign n15371 =  ( wr_addr ) == ( bv_8_100_n269 )  ;
assign n15372 =  ( n15370 ) & (n15371 )  ;
assign n15373 =  ( n15372 ) & (wr )  ;
assign n15374 =  ( n15373 ) ? ( n5071 ) : ( iram_100 ) ;
assign n15375 = wr_addr[7:7] ;
assign n15376 =  ( n15375 ) == ( bv_1_0_n53 )  ;
assign n15377 =  ( wr_addr ) == ( bv_8_100_n269 )  ;
assign n15378 =  ( n15376 ) & (n15377 )  ;
assign n15379 =  ( n15378 ) & (wr )  ;
assign n15380 =  ( n15379 ) ? ( n5096 ) : ( iram_100 ) ;
assign n15381 = wr_addr[7:7] ;
assign n15382 =  ( n15381 ) == ( bv_1_0_n53 )  ;
assign n15383 =  ( wr_addr ) == ( bv_8_100_n269 )  ;
assign n15384 =  ( n15382 ) & (n15383 )  ;
assign n15385 =  ( n15384 ) & (wr )  ;
assign n15386 =  ( n15385 ) ? ( n5123 ) : ( iram_100 ) ;
assign n15387 = wr_addr[7:7] ;
assign n15388 =  ( n15387 ) == ( bv_1_0_n53 )  ;
assign n15389 =  ( wr_addr ) == ( bv_8_100_n269 )  ;
assign n15390 =  ( n15388 ) & (n15389 )  ;
assign n15391 =  ( n15390 ) & (wr )  ;
assign n15392 =  ( n15391 ) ? ( n5165 ) : ( iram_100 ) ;
assign n15393 = wr_addr[7:7] ;
assign n15394 =  ( n15393 ) == ( bv_1_0_n53 )  ;
assign n15395 =  ( wr_addr ) == ( bv_8_100_n269 )  ;
assign n15396 =  ( n15394 ) & (n15395 )  ;
assign n15397 =  ( n15396 ) & (wr )  ;
assign n15398 =  ( n15397 ) ? ( n5204 ) : ( iram_100 ) ;
assign n15399 = wr_addr[7:7] ;
assign n15400 =  ( n15399 ) == ( bv_1_0_n53 )  ;
assign n15401 =  ( wr_addr ) == ( bv_8_100_n269 )  ;
assign n15402 =  ( n15400 ) & (n15401 )  ;
assign n15403 =  ( n15402 ) & (wr )  ;
assign n15404 =  ( n15403 ) ? ( n5262 ) : ( iram_100 ) ;
assign n15405 = wr_addr[7:7] ;
assign n15406 =  ( n15405 ) == ( bv_1_0_n53 )  ;
assign n15407 =  ( wr_addr ) == ( bv_8_100_n269 )  ;
assign n15408 =  ( n15406 ) & (n15407 )  ;
assign n15409 =  ( n15408 ) & (wr )  ;
assign n15410 =  ( n15409 ) ? ( n5298 ) : ( iram_100 ) ;
assign n15411 = wr_addr[7:7] ;
assign n15412 =  ( n15411 ) == ( bv_1_0_n53 )  ;
assign n15413 =  ( wr_addr ) == ( bv_8_100_n269 )  ;
assign n15414 =  ( n15412 ) & (n15413 )  ;
assign n15415 =  ( n15414 ) & (wr )  ;
assign n15416 =  ( n15415 ) ? ( n5325 ) : ( iram_100 ) ;
assign n15417 = wr_addr[7:7] ;
assign n15418 =  ( n15417 ) == ( bv_1_0_n53 )  ;
assign n15419 =  ( wr_addr ) == ( bv_8_101_n271 )  ;
assign n15420 =  ( n15418 ) & (n15419 )  ;
assign n15421 =  ( n15420 ) & (wr )  ;
assign n15422 =  ( n15421 ) ? ( n4782 ) : ( iram_101 ) ;
assign n15423 = wr_addr[7:7] ;
assign n15424 =  ( n15423 ) == ( bv_1_0_n53 )  ;
assign n15425 =  ( wr_addr ) == ( bv_8_101_n271 )  ;
assign n15426 =  ( n15424 ) & (n15425 )  ;
assign n15427 =  ( n15426 ) & (wr )  ;
assign n15428 =  ( n15427 ) ? ( n4841 ) : ( iram_101 ) ;
assign n15429 = wr_addr[7:7] ;
assign n15430 =  ( n15429 ) == ( bv_1_0_n53 )  ;
assign n15431 =  ( wr_addr ) == ( bv_8_101_n271 )  ;
assign n15432 =  ( n15430 ) & (n15431 )  ;
assign n15433 =  ( n15432 ) & (wr )  ;
assign n15434 =  ( n15433 ) ? ( n5449 ) : ( iram_101 ) ;
assign n15435 = wr_addr[7:7] ;
assign n15436 =  ( n15435 ) == ( bv_1_0_n53 )  ;
assign n15437 =  ( wr_addr ) == ( bv_8_101_n271 )  ;
assign n15438 =  ( n15436 ) & (n15437 )  ;
assign n15439 =  ( n15438 ) & (wr )  ;
assign n15440 =  ( n15439 ) ? ( n4906 ) : ( iram_101 ) ;
assign n15441 = wr_addr[7:7] ;
assign n15442 =  ( n15441 ) == ( bv_1_0_n53 )  ;
assign n15443 =  ( wr_addr ) == ( bv_8_101_n271 )  ;
assign n15444 =  ( n15442 ) & (n15443 )  ;
assign n15445 =  ( n15444 ) & (wr )  ;
assign n15446 =  ( n15445 ) ? ( n5485 ) : ( iram_101 ) ;
assign n15447 = wr_addr[7:7] ;
assign n15448 =  ( n15447 ) == ( bv_1_0_n53 )  ;
assign n15449 =  ( wr_addr ) == ( bv_8_101_n271 )  ;
assign n15450 =  ( n15448 ) & (n15449 )  ;
assign n15451 =  ( n15450 ) & (wr )  ;
assign n15452 =  ( n15451 ) ? ( n5512 ) : ( iram_101 ) ;
assign n15453 = wr_addr[7:7] ;
assign n15454 =  ( n15453 ) == ( bv_1_0_n53 )  ;
assign n15455 =  ( wr_addr ) == ( bv_8_101_n271 )  ;
assign n15456 =  ( n15454 ) & (n15455 )  ;
assign n15457 =  ( n15456 ) & (wr )  ;
assign n15458 =  ( n15457 ) ? ( bv_8_0_n69 ) : ( iram_101 ) ;
assign n15459 = wr_addr[7:7] ;
assign n15460 =  ( n15459 ) == ( bv_1_0_n53 )  ;
assign n15461 =  ( wr_addr ) == ( bv_8_101_n271 )  ;
assign n15462 =  ( n15460 ) & (n15461 )  ;
assign n15463 =  ( n15462 ) & (wr )  ;
assign n15464 =  ( n15463 ) ? ( n5071 ) : ( iram_101 ) ;
assign n15465 = wr_addr[7:7] ;
assign n15466 =  ( n15465 ) == ( bv_1_0_n53 )  ;
assign n15467 =  ( wr_addr ) == ( bv_8_101_n271 )  ;
assign n15468 =  ( n15466 ) & (n15467 )  ;
assign n15469 =  ( n15468 ) & (wr )  ;
assign n15470 =  ( n15469 ) ? ( n5096 ) : ( iram_101 ) ;
assign n15471 = wr_addr[7:7] ;
assign n15472 =  ( n15471 ) == ( bv_1_0_n53 )  ;
assign n15473 =  ( wr_addr ) == ( bv_8_101_n271 )  ;
assign n15474 =  ( n15472 ) & (n15473 )  ;
assign n15475 =  ( n15474 ) & (wr )  ;
assign n15476 =  ( n15475 ) ? ( n5123 ) : ( iram_101 ) ;
assign n15477 = wr_addr[7:7] ;
assign n15478 =  ( n15477 ) == ( bv_1_0_n53 )  ;
assign n15479 =  ( wr_addr ) == ( bv_8_101_n271 )  ;
assign n15480 =  ( n15478 ) & (n15479 )  ;
assign n15481 =  ( n15480 ) & (wr )  ;
assign n15482 =  ( n15481 ) ? ( n5165 ) : ( iram_101 ) ;
assign n15483 = wr_addr[7:7] ;
assign n15484 =  ( n15483 ) == ( bv_1_0_n53 )  ;
assign n15485 =  ( wr_addr ) == ( bv_8_101_n271 )  ;
assign n15486 =  ( n15484 ) & (n15485 )  ;
assign n15487 =  ( n15486 ) & (wr )  ;
assign n15488 =  ( n15487 ) ? ( n5204 ) : ( iram_101 ) ;
assign n15489 = wr_addr[7:7] ;
assign n15490 =  ( n15489 ) == ( bv_1_0_n53 )  ;
assign n15491 =  ( wr_addr ) == ( bv_8_101_n271 )  ;
assign n15492 =  ( n15490 ) & (n15491 )  ;
assign n15493 =  ( n15492 ) & (wr )  ;
assign n15494 =  ( n15493 ) ? ( n5262 ) : ( iram_101 ) ;
assign n15495 = wr_addr[7:7] ;
assign n15496 =  ( n15495 ) == ( bv_1_0_n53 )  ;
assign n15497 =  ( wr_addr ) == ( bv_8_101_n271 )  ;
assign n15498 =  ( n15496 ) & (n15497 )  ;
assign n15499 =  ( n15498 ) & (wr )  ;
assign n15500 =  ( n15499 ) ? ( n5298 ) : ( iram_101 ) ;
assign n15501 = wr_addr[7:7] ;
assign n15502 =  ( n15501 ) == ( bv_1_0_n53 )  ;
assign n15503 =  ( wr_addr ) == ( bv_8_101_n271 )  ;
assign n15504 =  ( n15502 ) & (n15503 )  ;
assign n15505 =  ( n15504 ) & (wr )  ;
assign n15506 =  ( n15505 ) ? ( n5325 ) : ( iram_101 ) ;
assign n15507 = wr_addr[7:7] ;
assign n15508 =  ( n15507 ) == ( bv_1_0_n53 )  ;
assign n15509 =  ( wr_addr ) == ( bv_8_102_n273 )  ;
assign n15510 =  ( n15508 ) & (n15509 )  ;
assign n15511 =  ( n15510 ) & (wr )  ;
assign n15512 =  ( n15511 ) ? ( n4782 ) : ( iram_102 ) ;
assign n15513 = wr_addr[7:7] ;
assign n15514 =  ( n15513 ) == ( bv_1_0_n53 )  ;
assign n15515 =  ( wr_addr ) == ( bv_8_102_n273 )  ;
assign n15516 =  ( n15514 ) & (n15515 )  ;
assign n15517 =  ( n15516 ) & (wr )  ;
assign n15518 =  ( n15517 ) ? ( n4841 ) : ( iram_102 ) ;
assign n15519 = wr_addr[7:7] ;
assign n15520 =  ( n15519 ) == ( bv_1_0_n53 )  ;
assign n15521 =  ( wr_addr ) == ( bv_8_102_n273 )  ;
assign n15522 =  ( n15520 ) & (n15521 )  ;
assign n15523 =  ( n15522 ) & (wr )  ;
assign n15524 =  ( n15523 ) ? ( n5449 ) : ( iram_102 ) ;
assign n15525 = wr_addr[7:7] ;
assign n15526 =  ( n15525 ) == ( bv_1_0_n53 )  ;
assign n15527 =  ( wr_addr ) == ( bv_8_102_n273 )  ;
assign n15528 =  ( n15526 ) & (n15527 )  ;
assign n15529 =  ( n15528 ) & (wr )  ;
assign n15530 =  ( n15529 ) ? ( n4906 ) : ( iram_102 ) ;
assign n15531 = wr_addr[7:7] ;
assign n15532 =  ( n15531 ) == ( bv_1_0_n53 )  ;
assign n15533 =  ( wr_addr ) == ( bv_8_102_n273 )  ;
assign n15534 =  ( n15532 ) & (n15533 )  ;
assign n15535 =  ( n15534 ) & (wr )  ;
assign n15536 =  ( n15535 ) ? ( n5485 ) : ( iram_102 ) ;
assign n15537 = wr_addr[7:7] ;
assign n15538 =  ( n15537 ) == ( bv_1_0_n53 )  ;
assign n15539 =  ( wr_addr ) == ( bv_8_102_n273 )  ;
assign n15540 =  ( n15538 ) & (n15539 )  ;
assign n15541 =  ( n15540 ) & (wr )  ;
assign n15542 =  ( n15541 ) ? ( n5512 ) : ( iram_102 ) ;
assign n15543 = wr_addr[7:7] ;
assign n15544 =  ( n15543 ) == ( bv_1_0_n53 )  ;
assign n15545 =  ( wr_addr ) == ( bv_8_102_n273 )  ;
assign n15546 =  ( n15544 ) & (n15545 )  ;
assign n15547 =  ( n15546 ) & (wr )  ;
assign n15548 =  ( n15547 ) ? ( bv_8_0_n69 ) : ( iram_102 ) ;
assign n15549 = wr_addr[7:7] ;
assign n15550 =  ( n15549 ) == ( bv_1_0_n53 )  ;
assign n15551 =  ( wr_addr ) == ( bv_8_102_n273 )  ;
assign n15552 =  ( n15550 ) & (n15551 )  ;
assign n15553 =  ( n15552 ) & (wr )  ;
assign n15554 =  ( n15553 ) ? ( n5071 ) : ( iram_102 ) ;
assign n15555 = wr_addr[7:7] ;
assign n15556 =  ( n15555 ) == ( bv_1_0_n53 )  ;
assign n15557 =  ( wr_addr ) == ( bv_8_102_n273 )  ;
assign n15558 =  ( n15556 ) & (n15557 )  ;
assign n15559 =  ( n15558 ) & (wr )  ;
assign n15560 =  ( n15559 ) ? ( n5096 ) : ( iram_102 ) ;
assign n15561 = wr_addr[7:7] ;
assign n15562 =  ( n15561 ) == ( bv_1_0_n53 )  ;
assign n15563 =  ( wr_addr ) == ( bv_8_102_n273 )  ;
assign n15564 =  ( n15562 ) & (n15563 )  ;
assign n15565 =  ( n15564 ) & (wr )  ;
assign n15566 =  ( n15565 ) ? ( n5123 ) : ( iram_102 ) ;
assign n15567 = wr_addr[7:7] ;
assign n15568 =  ( n15567 ) == ( bv_1_0_n53 )  ;
assign n15569 =  ( wr_addr ) == ( bv_8_102_n273 )  ;
assign n15570 =  ( n15568 ) & (n15569 )  ;
assign n15571 =  ( n15570 ) & (wr )  ;
assign n15572 =  ( n15571 ) ? ( n5165 ) : ( iram_102 ) ;
assign n15573 = wr_addr[7:7] ;
assign n15574 =  ( n15573 ) == ( bv_1_0_n53 )  ;
assign n15575 =  ( wr_addr ) == ( bv_8_102_n273 )  ;
assign n15576 =  ( n15574 ) & (n15575 )  ;
assign n15577 =  ( n15576 ) & (wr )  ;
assign n15578 =  ( n15577 ) ? ( n5204 ) : ( iram_102 ) ;
assign n15579 = wr_addr[7:7] ;
assign n15580 =  ( n15579 ) == ( bv_1_0_n53 )  ;
assign n15581 =  ( wr_addr ) == ( bv_8_102_n273 )  ;
assign n15582 =  ( n15580 ) & (n15581 )  ;
assign n15583 =  ( n15582 ) & (wr )  ;
assign n15584 =  ( n15583 ) ? ( n5262 ) : ( iram_102 ) ;
assign n15585 = wr_addr[7:7] ;
assign n15586 =  ( n15585 ) == ( bv_1_0_n53 )  ;
assign n15587 =  ( wr_addr ) == ( bv_8_102_n273 )  ;
assign n15588 =  ( n15586 ) & (n15587 )  ;
assign n15589 =  ( n15588 ) & (wr )  ;
assign n15590 =  ( n15589 ) ? ( n5298 ) : ( iram_102 ) ;
assign n15591 = wr_addr[7:7] ;
assign n15592 =  ( n15591 ) == ( bv_1_0_n53 )  ;
assign n15593 =  ( wr_addr ) == ( bv_8_102_n273 )  ;
assign n15594 =  ( n15592 ) & (n15593 )  ;
assign n15595 =  ( n15594 ) & (wr )  ;
assign n15596 =  ( n15595 ) ? ( n5325 ) : ( iram_102 ) ;
assign n15597 = wr_addr[7:7] ;
assign n15598 =  ( n15597 ) == ( bv_1_0_n53 )  ;
assign n15599 =  ( wr_addr ) == ( bv_8_103_n275 )  ;
assign n15600 =  ( n15598 ) & (n15599 )  ;
assign n15601 =  ( n15600 ) & (wr )  ;
assign n15602 =  ( n15601 ) ? ( n4782 ) : ( iram_103 ) ;
assign n15603 = wr_addr[7:7] ;
assign n15604 =  ( n15603 ) == ( bv_1_0_n53 )  ;
assign n15605 =  ( wr_addr ) == ( bv_8_103_n275 )  ;
assign n15606 =  ( n15604 ) & (n15605 )  ;
assign n15607 =  ( n15606 ) & (wr )  ;
assign n15608 =  ( n15607 ) ? ( n4841 ) : ( iram_103 ) ;
assign n15609 = wr_addr[7:7] ;
assign n15610 =  ( n15609 ) == ( bv_1_0_n53 )  ;
assign n15611 =  ( wr_addr ) == ( bv_8_103_n275 )  ;
assign n15612 =  ( n15610 ) & (n15611 )  ;
assign n15613 =  ( n15612 ) & (wr )  ;
assign n15614 =  ( n15613 ) ? ( n5449 ) : ( iram_103 ) ;
assign n15615 = wr_addr[7:7] ;
assign n15616 =  ( n15615 ) == ( bv_1_0_n53 )  ;
assign n15617 =  ( wr_addr ) == ( bv_8_103_n275 )  ;
assign n15618 =  ( n15616 ) & (n15617 )  ;
assign n15619 =  ( n15618 ) & (wr )  ;
assign n15620 =  ( n15619 ) ? ( n4906 ) : ( iram_103 ) ;
assign n15621 = wr_addr[7:7] ;
assign n15622 =  ( n15621 ) == ( bv_1_0_n53 )  ;
assign n15623 =  ( wr_addr ) == ( bv_8_103_n275 )  ;
assign n15624 =  ( n15622 ) & (n15623 )  ;
assign n15625 =  ( n15624 ) & (wr )  ;
assign n15626 =  ( n15625 ) ? ( n5485 ) : ( iram_103 ) ;
assign n15627 = wr_addr[7:7] ;
assign n15628 =  ( n15627 ) == ( bv_1_0_n53 )  ;
assign n15629 =  ( wr_addr ) == ( bv_8_103_n275 )  ;
assign n15630 =  ( n15628 ) & (n15629 )  ;
assign n15631 =  ( n15630 ) & (wr )  ;
assign n15632 =  ( n15631 ) ? ( n5512 ) : ( iram_103 ) ;
assign n15633 = wr_addr[7:7] ;
assign n15634 =  ( n15633 ) == ( bv_1_0_n53 )  ;
assign n15635 =  ( wr_addr ) == ( bv_8_103_n275 )  ;
assign n15636 =  ( n15634 ) & (n15635 )  ;
assign n15637 =  ( n15636 ) & (wr )  ;
assign n15638 =  ( n15637 ) ? ( bv_8_0_n69 ) : ( iram_103 ) ;
assign n15639 = wr_addr[7:7] ;
assign n15640 =  ( n15639 ) == ( bv_1_0_n53 )  ;
assign n15641 =  ( wr_addr ) == ( bv_8_103_n275 )  ;
assign n15642 =  ( n15640 ) & (n15641 )  ;
assign n15643 =  ( n15642 ) & (wr )  ;
assign n15644 =  ( n15643 ) ? ( n5071 ) : ( iram_103 ) ;
assign n15645 = wr_addr[7:7] ;
assign n15646 =  ( n15645 ) == ( bv_1_0_n53 )  ;
assign n15647 =  ( wr_addr ) == ( bv_8_103_n275 )  ;
assign n15648 =  ( n15646 ) & (n15647 )  ;
assign n15649 =  ( n15648 ) & (wr )  ;
assign n15650 =  ( n15649 ) ? ( n5096 ) : ( iram_103 ) ;
assign n15651 = wr_addr[7:7] ;
assign n15652 =  ( n15651 ) == ( bv_1_0_n53 )  ;
assign n15653 =  ( wr_addr ) == ( bv_8_103_n275 )  ;
assign n15654 =  ( n15652 ) & (n15653 )  ;
assign n15655 =  ( n15654 ) & (wr )  ;
assign n15656 =  ( n15655 ) ? ( n5123 ) : ( iram_103 ) ;
assign n15657 = wr_addr[7:7] ;
assign n15658 =  ( n15657 ) == ( bv_1_0_n53 )  ;
assign n15659 =  ( wr_addr ) == ( bv_8_103_n275 )  ;
assign n15660 =  ( n15658 ) & (n15659 )  ;
assign n15661 =  ( n15660 ) & (wr )  ;
assign n15662 =  ( n15661 ) ? ( n5165 ) : ( iram_103 ) ;
assign n15663 = wr_addr[7:7] ;
assign n15664 =  ( n15663 ) == ( bv_1_0_n53 )  ;
assign n15665 =  ( wr_addr ) == ( bv_8_103_n275 )  ;
assign n15666 =  ( n15664 ) & (n15665 )  ;
assign n15667 =  ( n15666 ) & (wr )  ;
assign n15668 =  ( n15667 ) ? ( n5204 ) : ( iram_103 ) ;
assign n15669 = wr_addr[7:7] ;
assign n15670 =  ( n15669 ) == ( bv_1_0_n53 )  ;
assign n15671 =  ( wr_addr ) == ( bv_8_103_n275 )  ;
assign n15672 =  ( n15670 ) & (n15671 )  ;
assign n15673 =  ( n15672 ) & (wr )  ;
assign n15674 =  ( n15673 ) ? ( n5262 ) : ( iram_103 ) ;
assign n15675 = wr_addr[7:7] ;
assign n15676 =  ( n15675 ) == ( bv_1_0_n53 )  ;
assign n15677 =  ( wr_addr ) == ( bv_8_103_n275 )  ;
assign n15678 =  ( n15676 ) & (n15677 )  ;
assign n15679 =  ( n15678 ) & (wr )  ;
assign n15680 =  ( n15679 ) ? ( n5298 ) : ( iram_103 ) ;
assign n15681 = wr_addr[7:7] ;
assign n15682 =  ( n15681 ) == ( bv_1_0_n53 )  ;
assign n15683 =  ( wr_addr ) == ( bv_8_103_n275 )  ;
assign n15684 =  ( n15682 ) & (n15683 )  ;
assign n15685 =  ( n15684 ) & (wr )  ;
assign n15686 =  ( n15685 ) ? ( n5325 ) : ( iram_103 ) ;
assign n15687 = wr_addr[7:7] ;
assign n15688 =  ( n15687 ) == ( bv_1_0_n53 )  ;
assign n15689 =  ( wr_addr ) == ( bv_8_104_n277 )  ;
assign n15690 =  ( n15688 ) & (n15689 )  ;
assign n15691 =  ( n15690 ) & (wr )  ;
assign n15692 =  ( n15691 ) ? ( n4782 ) : ( iram_104 ) ;
assign n15693 = wr_addr[7:7] ;
assign n15694 =  ( n15693 ) == ( bv_1_0_n53 )  ;
assign n15695 =  ( wr_addr ) == ( bv_8_104_n277 )  ;
assign n15696 =  ( n15694 ) & (n15695 )  ;
assign n15697 =  ( n15696 ) & (wr )  ;
assign n15698 =  ( n15697 ) ? ( n4841 ) : ( iram_104 ) ;
assign n15699 = wr_addr[7:7] ;
assign n15700 =  ( n15699 ) == ( bv_1_0_n53 )  ;
assign n15701 =  ( wr_addr ) == ( bv_8_104_n277 )  ;
assign n15702 =  ( n15700 ) & (n15701 )  ;
assign n15703 =  ( n15702 ) & (wr )  ;
assign n15704 =  ( n15703 ) ? ( n5449 ) : ( iram_104 ) ;
assign n15705 = wr_addr[7:7] ;
assign n15706 =  ( n15705 ) == ( bv_1_0_n53 )  ;
assign n15707 =  ( wr_addr ) == ( bv_8_104_n277 )  ;
assign n15708 =  ( n15706 ) & (n15707 )  ;
assign n15709 =  ( n15708 ) & (wr )  ;
assign n15710 =  ( n15709 ) ? ( n4906 ) : ( iram_104 ) ;
assign n15711 = wr_addr[7:7] ;
assign n15712 =  ( n15711 ) == ( bv_1_0_n53 )  ;
assign n15713 =  ( wr_addr ) == ( bv_8_104_n277 )  ;
assign n15714 =  ( n15712 ) & (n15713 )  ;
assign n15715 =  ( n15714 ) & (wr )  ;
assign n15716 =  ( n15715 ) ? ( n5485 ) : ( iram_104 ) ;
assign n15717 = wr_addr[7:7] ;
assign n15718 =  ( n15717 ) == ( bv_1_0_n53 )  ;
assign n15719 =  ( wr_addr ) == ( bv_8_104_n277 )  ;
assign n15720 =  ( n15718 ) & (n15719 )  ;
assign n15721 =  ( n15720 ) & (wr )  ;
assign n15722 =  ( n15721 ) ? ( n5512 ) : ( iram_104 ) ;
assign n15723 = wr_addr[7:7] ;
assign n15724 =  ( n15723 ) == ( bv_1_0_n53 )  ;
assign n15725 =  ( wr_addr ) == ( bv_8_104_n277 )  ;
assign n15726 =  ( n15724 ) & (n15725 )  ;
assign n15727 =  ( n15726 ) & (wr )  ;
assign n15728 =  ( n15727 ) ? ( bv_8_0_n69 ) : ( iram_104 ) ;
assign n15729 = wr_addr[7:7] ;
assign n15730 =  ( n15729 ) == ( bv_1_0_n53 )  ;
assign n15731 =  ( wr_addr ) == ( bv_8_104_n277 )  ;
assign n15732 =  ( n15730 ) & (n15731 )  ;
assign n15733 =  ( n15732 ) & (wr )  ;
assign n15734 =  ( n15733 ) ? ( n5071 ) : ( iram_104 ) ;
assign n15735 = wr_addr[7:7] ;
assign n15736 =  ( n15735 ) == ( bv_1_0_n53 )  ;
assign n15737 =  ( wr_addr ) == ( bv_8_104_n277 )  ;
assign n15738 =  ( n15736 ) & (n15737 )  ;
assign n15739 =  ( n15738 ) & (wr )  ;
assign n15740 =  ( n15739 ) ? ( n5096 ) : ( iram_104 ) ;
assign n15741 = wr_addr[7:7] ;
assign n15742 =  ( n15741 ) == ( bv_1_0_n53 )  ;
assign n15743 =  ( wr_addr ) == ( bv_8_104_n277 )  ;
assign n15744 =  ( n15742 ) & (n15743 )  ;
assign n15745 =  ( n15744 ) & (wr )  ;
assign n15746 =  ( n15745 ) ? ( n5123 ) : ( iram_104 ) ;
assign n15747 = wr_addr[7:7] ;
assign n15748 =  ( n15747 ) == ( bv_1_0_n53 )  ;
assign n15749 =  ( wr_addr ) == ( bv_8_104_n277 )  ;
assign n15750 =  ( n15748 ) & (n15749 )  ;
assign n15751 =  ( n15750 ) & (wr )  ;
assign n15752 =  ( n15751 ) ? ( n5165 ) : ( iram_104 ) ;
assign n15753 = wr_addr[7:7] ;
assign n15754 =  ( n15753 ) == ( bv_1_0_n53 )  ;
assign n15755 =  ( wr_addr ) == ( bv_8_104_n277 )  ;
assign n15756 =  ( n15754 ) & (n15755 )  ;
assign n15757 =  ( n15756 ) & (wr )  ;
assign n15758 =  ( n15757 ) ? ( n5204 ) : ( iram_104 ) ;
assign n15759 = wr_addr[7:7] ;
assign n15760 =  ( n15759 ) == ( bv_1_0_n53 )  ;
assign n15761 =  ( wr_addr ) == ( bv_8_104_n277 )  ;
assign n15762 =  ( n15760 ) & (n15761 )  ;
assign n15763 =  ( n15762 ) & (wr )  ;
assign n15764 =  ( n15763 ) ? ( n5262 ) : ( iram_104 ) ;
assign n15765 = wr_addr[7:7] ;
assign n15766 =  ( n15765 ) == ( bv_1_0_n53 )  ;
assign n15767 =  ( wr_addr ) == ( bv_8_104_n277 )  ;
assign n15768 =  ( n15766 ) & (n15767 )  ;
assign n15769 =  ( n15768 ) & (wr )  ;
assign n15770 =  ( n15769 ) ? ( n5298 ) : ( iram_104 ) ;
assign n15771 = wr_addr[7:7] ;
assign n15772 =  ( n15771 ) == ( bv_1_0_n53 )  ;
assign n15773 =  ( wr_addr ) == ( bv_8_104_n277 )  ;
assign n15774 =  ( n15772 ) & (n15773 )  ;
assign n15775 =  ( n15774 ) & (wr )  ;
assign n15776 =  ( n15775 ) ? ( n5325 ) : ( iram_104 ) ;
assign n15777 = wr_addr[7:7] ;
assign n15778 =  ( n15777 ) == ( bv_1_0_n53 )  ;
assign n15779 =  ( wr_addr ) == ( bv_8_105_n279 )  ;
assign n15780 =  ( n15778 ) & (n15779 )  ;
assign n15781 =  ( n15780 ) & (wr )  ;
assign n15782 =  ( n15781 ) ? ( n4782 ) : ( iram_105 ) ;
assign n15783 = wr_addr[7:7] ;
assign n15784 =  ( n15783 ) == ( bv_1_0_n53 )  ;
assign n15785 =  ( wr_addr ) == ( bv_8_105_n279 )  ;
assign n15786 =  ( n15784 ) & (n15785 )  ;
assign n15787 =  ( n15786 ) & (wr )  ;
assign n15788 =  ( n15787 ) ? ( n4841 ) : ( iram_105 ) ;
assign n15789 = wr_addr[7:7] ;
assign n15790 =  ( n15789 ) == ( bv_1_0_n53 )  ;
assign n15791 =  ( wr_addr ) == ( bv_8_105_n279 )  ;
assign n15792 =  ( n15790 ) & (n15791 )  ;
assign n15793 =  ( n15792 ) & (wr )  ;
assign n15794 =  ( n15793 ) ? ( n5449 ) : ( iram_105 ) ;
assign n15795 = wr_addr[7:7] ;
assign n15796 =  ( n15795 ) == ( bv_1_0_n53 )  ;
assign n15797 =  ( wr_addr ) == ( bv_8_105_n279 )  ;
assign n15798 =  ( n15796 ) & (n15797 )  ;
assign n15799 =  ( n15798 ) & (wr )  ;
assign n15800 =  ( n15799 ) ? ( n4906 ) : ( iram_105 ) ;
assign n15801 = wr_addr[7:7] ;
assign n15802 =  ( n15801 ) == ( bv_1_0_n53 )  ;
assign n15803 =  ( wr_addr ) == ( bv_8_105_n279 )  ;
assign n15804 =  ( n15802 ) & (n15803 )  ;
assign n15805 =  ( n15804 ) & (wr )  ;
assign n15806 =  ( n15805 ) ? ( n5485 ) : ( iram_105 ) ;
assign n15807 = wr_addr[7:7] ;
assign n15808 =  ( n15807 ) == ( bv_1_0_n53 )  ;
assign n15809 =  ( wr_addr ) == ( bv_8_105_n279 )  ;
assign n15810 =  ( n15808 ) & (n15809 )  ;
assign n15811 =  ( n15810 ) & (wr )  ;
assign n15812 =  ( n15811 ) ? ( n5512 ) : ( iram_105 ) ;
assign n15813 = wr_addr[7:7] ;
assign n15814 =  ( n15813 ) == ( bv_1_0_n53 )  ;
assign n15815 =  ( wr_addr ) == ( bv_8_105_n279 )  ;
assign n15816 =  ( n15814 ) & (n15815 )  ;
assign n15817 =  ( n15816 ) & (wr )  ;
assign n15818 =  ( n15817 ) ? ( bv_8_0_n69 ) : ( iram_105 ) ;
assign n15819 = wr_addr[7:7] ;
assign n15820 =  ( n15819 ) == ( bv_1_0_n53 )  ;
assign n15821 =  ( wr_addr ) == ( bv_8_105_n279 )  ;
assign n15822 =  ( n15820 ) & (n15821 )  ;
assign n15823 =  ( n15822 ) & (wr )  ;
assign n15824 =  ( n15823 ) ? ( n5071 ) : ( iram_105 ) ;
assign n15825 = wr_addr[7:7] ;
assign n15826 =  ( n15825 ) == ( bv_1_0_n53 )  ;
assign n15827 =  ( wr_addr ) == ( bv_8_105_n279 )  ;
assign n15828 =  ( n15826 ) & (n15827 )  ;
assign n15829 =  ( n15828 ) & (wr )  ;
assign n15830 =  ( n15829 ) ? ( n5096 ) : ( iram_105 ) ;
assign n15831 = wr_addr[7:7] ;
assign n15832 =  ( n15831 ) == ( bv_1_0_n53 )  ;
assign n15833 =  ( wr_addr ) == ( bv_8_105_n279 )  ;
assign n15834 =  ( n15832 ) & (n15833 )  ;
assign n15835 =  ( n15834 ) & (wr )  ;
assign n15836 =  ( n15835 ) ? ( n5123 ) : ( iram_105 ) ;
assign n15837 = wr_addr[7:7] ;
assign n15838 =  ( n15837 ) == ( bv_1_0_n53 )  ;
assign n15839 =  ( wr_addr ) == ( bv_8_105_n279 )  ;
assign n15840 =  ( n15838 ) & (n15839 )  ;
assign n15841 =  ( n15840 ) & (wr )  ;
assign n15842 =  ( n15841 ) ? ( n5165 ) : ( iram_105 ) ;
assign n15843 = wr_addr[7:7] ;
assign n15844 =  ( n15843 ) == ( bv_1_0_n53 )  ;
assign n15845 =  ( wr_addr ) == ( bv_8_105_n279 )  ;
assign n15846 =  ( n15844 ) & (n15845 )  ;
assign n15847 =  ( n15846 ) & (wr )  ;
assign n15848 =  ( n15847 ) ? ( n5204 ) : ( iram_105 ) ;
assign n15849 = wr_addr[7:7] ;
assign n15850 =  ( n15849 ) == ( bv_1_0_n53 )  ;
assign n15851 =  ( wr_addr ) == ( bv_8_105_n279 )  ;
assign n15852 =  ( n15850 ) & (n15851 )  ;
assign n15853 =  ( n15852 ) & (wr )  ;
assign n15854 =  ( n15853 ) ? ( n5262 ) : ( iram_105 ) ;
assign n15855 = wr_addr[7:7] ;
assign n15856 =  ( n15855 ) == ( bv_1_0_n53 )  ;
assign n15857 =  ( wr_addr ) == ( bv_8_105_n279 )  ;
assign n15858 =  ( n15856 ) & (n15857 )  ;
assign n15859 =  ( n15858 ) & (wr )  ;
assign n15860 =  ( n15859 ) ? ( n5298 ) : ( iram_105 ) ;
assign n15861 = wr_addr[7:7] ;
assign n15862 =  ( n15861 ) == ( bv_1_0_n53 )  ;
assign n15863 =  ( wr_addr ) == ( bv_8_105_n279 )  ;
assign n15864 =  ( n15862 ) & (n15863 )  ;
assign n15865 =  ( n15864 ) & (wr )  ;
assign n15866 =  ( n15865 ) ? ( n5325 ) : ( iram_105 ) ;
assign n15867 = wr_addr[7:7] ;
assign n15868 =  ( n15867 ) == ( bv_1_0_n53 )  ;
assign n15869 =  ( wr_addr ) == ( bv_8_106_n281 )  ;
assign n15870 =  ( n15868 ) & (n15869 )  ;
assign n15871 =  ( n15870 ) & (wr )  ;
assign n15872 =  ( n15871 ) ? ( n4782 ) : ( iram_106 ) ;
assign n15873 = wr_addr[7:7] ;
assign n15874 =  ( n15873 ) == ( bv_1_0_n53 )  ;
assign n15875 =  ( wr_addr ) == ( bv_8_106_n281 )  ;
assign n15876 =  ( n15874 ) & (n15875 )  ;
assign n15877 =  ( n15876 ) & (wr )  ;
assign n15878 =  ( n15877 ) ? ( n4841 ) : ( iram_106 ) ;
assign n15879 = wr_addr[7:7] ;
assign n15880 =  ( n15879 ) == ( bv_1_0_n53 )  ;
assign n15881 =  ( wr_addr ) == ( bv_8_106_n281 )  ;
assign n15882 =  ( n15880 ) & (n15881 )  ;
assign n15883 =  ( n15882 ) & (wr )  ;
assign n15884 =  ( n15883 ) ? ( n5449 ) : ( iram_106 ) ;
assign n15885 = wr_addr[7:7] ;
assign n15886 =  ( n15885 ) == ( bv_1_0_n53 )  ;
assign n15887 =  ( wr_addr ) == ( bv_8_106_n281 )  ;
assign n15888 =  ( n15886 ) & (n15887 )  ;
assign n15889 =  ( n15888 ) & (wr )  ;
assign n15890 =  ( n15889 ) ? ( n4906 ) : ( iram_106 ) ;
assign n15891 = wr_addr[7:7] ;
assign n15892 =  ( n15891 ) == ( bv_1_0_n53 )  ;
assign n15893 =  ( wr_addr ) == ( bv_8_106_n281 )  ;
assign n15894 =  ( n15892 ) & (n15893 )  ;
assign n15895 =  ( n15894 ) & (wr )  ;
assign n15896 =  ( n15895 ) ? ( n5485 ) : ( iram_106 ) ;
assign n15897 = wr_addr[7:7] ;
assign n15898 =  ( n15897 ) == ( bv_1_0_n53 )  ;
assign n15899 =  ( wr_addr ) == ( bv_8_106_n281 )  ;
assign n15900 =  ( n15898 ) & (n15899 )  ;
assign n15901 =  ( n15900 ) & (wr )  ;
assign n15902 =  ( n15901 ) ? ( n5512 ) : ( iram_106 ) ;
assign n15903 = wr_addr[7:7] ;
assign n15904 =  ( n15903 ) == ( bv_1_0_n53 )  ;
assign n15905 =  ( wr_addr ) == ( bv_8_106_n281 )  ;
assign n15906 =  ( n15904 ) & (n15905 )  ;
assign n15907 =  ( n15906 ) & (wr )  ;
assign n15908 =  ( n15907 ) ? ( bv_8_0_n69 ) : ( iram_106 ) ;
assign n15909 = wr_addr[7:7] ;
assign n15910 =  ( n15909 ) == ( bv_1_0_n53 )  ;
assign n15911 =  ( wr_addr ) == ( bv_8_106_n281 )  ;
assign n15912 =  ( n15910 ) & (n15911 )  ;
assign n15913 =  ( n15912 ) & (wr )  ;
assign n15914 =  ( n15913 ) ? ( n5071 ) : ( iram_106 ) ;
assign n15915 = wr_addr[7:7] ;
assign n15916 =  ( n15915 ) == ( bv_1_0_n53 )  ;
assign n15917 =  ( wr_addr ) == ( bv_8_106_n281 )  ;
assign n15918 =  ( n15916 ) & (n15917 )  ;
assign n15919 =  ( n15918 ) & (wr )  ;
assign n15920 =  ( n15919 ) ? ( n5096 ) : ( iram_106 ) ;
assign n15921 = wr_addr[7:7] ;
assign n15922 =  ( n15921 ) == ( bv_1_0_n53 )  ;
assign n15923 =  ( wr_addr ) == ( bv_8_106_n281 )  ;
assign n15924 =  ( n15922 ) & (n15923 )  ;
assign n15925 =  ( n15924 ) & (wr )  ;
assign n15926 =  ( n15925 ) ? ( n5123 ) : ( iram_106 ) ;
assign n15927 = wr_addr[7:7] ;
assign n15928 =  ( n15927 ) == ( bv_1_0_n53 )  ;
assign n15929 =  ( wr_addr ) == ( bv_8_106_n281 )  ;
assign n15930 =  ( n15928 ) & (n15929 )  ;
assign n15931 =  ( n15930 ) & (wr )  ;
assign n15932 =  ( n15931 ) ? ( n5165 ) : ( iram_106 ) ;
assign n15933 = wr_addr[7:7] ;
assign n15934 =  ( n15933 ) == ( bv_1_0_n53 )  ;
assign n15935 =  ( wr_addr ) == ( bv_8_106_n281 )  ;
assign n15936 =  ( n15934 ) & (n15935 )  ;
assign n15937 =  ( n15936 ) & (wr )  ;
assign n15938 =  ( n15937 ) ? ( n5204 ) : ( iram_106 ) ;
assign n15939 = wr_addr[7:7] ;
assign n15940 =  ( n15939 ) == ( bv_1_0_n53 )  ;
assign n15941 =  ( wr_addr ) == ( bv_8_106_n281 )  ;
assign n15942 =  ( n15940 ) & (n15941 )  ;
assign n15943 =  ( n15942 ) & (wr )  ;
assign n15944 =  ( n15943 ) ? ( n5262 ) : ( iram_106 ) ;
assign n15945 = wr_addr[7:7] ;
assign n15946 =  ( n15945 ) == ( bv_1_0_n53 )  ;
assign n15947 =  ( wr_addr ) == ( bv_8_106_n281 )  ;
assign n15948 =  ( n15946 ) & (n15947 )  ;
assign n15949 =  ( n15948 ) & (wr )  ;
assign n15950 =  ( n15949 ) ? ( n5298 ) : ( iram_106 ) ;
assign n15951 = wr_addr[7:7] ;
assign n15952 =  ( n15951 ) == ( bv_1_0_n53 )  ;
assign n15953 =  ( wr_addr ) == ( bv_8_106_n281 )  ;
assign n15954 =  ( n15952 ) & (n15953 )  ;
assign n15955 =  ( n15954 ) & (wr )  ;
assign n15956 =  ( n15955 ) ? ( n5325 ) : ( iram_106 ) ;
assign n15957 = wr_addr[7:7] ;
assign n15958 =  ( n15957 ) == ( bv_1_0_n53 )  ;
assign n15959 =  ( wr_addr ) == ( bv_8_107_n283 )  ;
assign n15960 =  ( n15958 ) & (n15959 )  ;
assign n15961 =  ( n15960 ) & (wr )  ;
assign n15962 =  ( n15961 ) ? ( n4782 ) : ( iram_107 ) ;
assign n15963 = wr_addr[7:7] ;
assign n15964 =  ( n15963 ) == ( bv_1_0_n53 )  ;
assign n15965 =  ( wr_addr ) == ( bv_8_107_n283 )  ;
assign n15966 =  ( n15964 ) & (n15965 )  ;
assign n15967 =  ( n15966 ) & (wr )  ;
assign n15968 =  ( n15967 ) ? ( n4841 ) : ( iram_107 ) ;
assign n15969 = wr_addr[7:7] ;
assign n15970 =  ( n15969 ) == ( bv_1_0_n53 )  ;
assign n15971 =  ( wr_addr ) == ( bv_8_107_n283 )  ;
assign n15972 =  ( n15970 ) & (n15971 )  ;
assign n15973 =  ( n15972 ) & (wr )  ;
assign n15974 =  ( n15973 ) ? ( n5449 ) : ( iram_107 ) ;
assign n15975 = wr_addr[7:7] ;
assign n15976 =  ( n15975 ) == ( bv_1_0_n53 )  ;
assign n15977 =  ( wr_addr ) == ( bv_8_107_n283 )  ;
assign n15978 =  ( n15976 ) & (n15977 )  ;
assign n15979 =  ( n15978 ) & (wr )  ;
assign n15980 =  ( n15979 ) ? ( n4906 ) : ( iram_107 ) ;
assign n15981 = wr_addr[7:7] ;
assign n15982 =  ( n15981 ) == ( bv_1_0_n53 )  ;
assign n15983 =  ( wr_addr ) == ( bv_8_107_n283 )  ;
assign n15984 =  ( n15982 ) & (n15983 )  ;
assign n15985 =  ( n15984 ) & (wr )  ;
assign n15986 =  ( n15985 ) ? ( n5485 ) : ( iram_107 ) ;
assign n15987 = wr_addr[7:7] ;
assign n15988 =  ( n15987 ) == ( bv_1_0_n53 )  ;
assign n15989 =  ( wr_addr ) == ( bv_8_107_n283 )  ;
assign n15990 =  ( n15988 ) & (n15989 )  ;
assign n15991 =  ( n15990 ) & (wr )  ;
assign n15992 =  ( n15991 ) ? ( n5512 ) : ( iram_107 ) ;
assign n15993 = wr_addr[7:7] ;
assign n15994 =  ( n15993 ) == ( bv_1_0_n53 )  ;
assign n15995 =  ( wr_addr ) == ( bv_8_107_n283 )  ;
assign n15996 =  ( n15994 ) & (n15995 )  ;
assign n15997 =  ( n15996 ) & (wr )  ;
assign n15998 =  ( n15997 ) ? ( bv_8_0_n69 ) : ( iram_107 ) ;
assign n15999 = wr_addr[7:7] ;
assign n16000 =  ( n15999 ) == ( bv_1_0_n53 )  ;
assign n16001 =  ( wr_addr ) == ( bv_8_107_n283 )  ;
assign n16002 =  ( n16000 ) & (n16001 )  ;
assign n16003 =  ( n16002 ) & (wr )  ;
assign n16004 =  ( n16003 ) ? ( n5071 ) : ( iram_107 ) ;
assign n16005 = wr_addr[7:7] ;
assign n16006 =  ( n16005 ) == ( bv_1_0_n53 )  ;
assign n16007 =  ( wr_addr ) == ( bv_8_107_n283 )  ;
assign n16008 =  ( n16006 ) & (n16007 )  ;
assign n16009 =  ( n16008 ) & (wr )  ;
assign n16010 =  ( n16009 ) ? ( n5096 ) : ( iram_107 ) ;
assign n16011 = wr_addr[7:7] ;
assign n16012 =  ( n16011 ) == ( bv_1_0_n53 )  ;
assign n16013 =  ( wr_addr ) == ( bv_8_107_n283 )  ;
assign n16014 =  ( n16012 ) & (n16013 )  ;
assign n16015 =  ( n16014 ) & (wr )  ;
assign n16016 =  ( n16015 ) ? ( n5123 ) : ( iram_107 ) ;
assign n16017 = wr_addr[7:7] ;
assign n16018 =  ( n16017 ) == ( bv_1_0_n53 )  ;
assign n16019 =  ( wr_addr ) == ( bv_8_107_n283 )  ;
assign n16020 =  ( n16018 ) & (n16019 )  ;
assign n16021 =  ( n16020 ) & (wr )  ;
assign n16022 =  ( n16021 ) ? ( n5165 ) : ( iram_107 ) ;
assign n16023 = wr_addr[7:7] ;
assign n16024 =  ( n16023 ) == ( bv_1_0_n53 )  ;
assign n16025 =  ( wr_addr ) == ( bv_8_107_n283 )  ;
assign n16026 =  ( n16024 ) & (n16025 )  ;
assign n16027 =  ( n16026 ) & (wr )  ;
assign n16028 =  ( n16027 ) ? ( n5204 ) : ( iram_107 ) ;
assign n16029 = wr_addr[7:7] ;
assign n16030 =  ( n16029 ) == ( bv_1_0_n53 )  ;
assign n16031 =  ( wr_addr ) == ( bv_8_107_n283 )  ;
assign n16032 =  ( n16030 ) & (n16031 )  ;
assign n16033 =  ( n16032 ) & (wr )  ;
assign n16034 =  ( n16033 ) ? ( n5262 ) : ( iram_107 ) ;
assign n16035 = wr_addr[7:7] ;
assign n16036 =  ( n16035 ) == ( bv_1_0_n53 )  ;
assign n16037 =  ( wr_addr ) == ( bv_8_107_n283 )  ;
assign n16038 =  ( n16036 ) & (n16037 )  ;
assign n16039 =  ( n16038 ) & (wr )  ;
assign n16040 =  ( n16039 ) ? ( n5298 ) : ( iram_107 ) ;
assign n16041 = wr_addr[7:7] ;
assign n16042 =  ( n16041 ) == ( bv_1_0_n53 )  ;
assign n16043 =  ( wr_addr ) == ( bv_8_107_n283 )  ;
assign n16044 =  ( n16042 ) & (n16043 )  ;
assign n16045 =  ( n16044 ) & (wr )  ;
assign n16046 =  ( n16045 ) ? ( n5325 ) : ( iram_107 ) ;
assign n16047 = wr_addr[7:7] ;
assign n16048 =  ( n16047 ) == ( bv_1_0_n53 )  ;
assign n16049 =  ( wr_addr ) == ( bv_8_108_n285 )  ;
assign n16050 =  ( n16048 ) & (n16049 )  ;
assign n16051 =  ( n16050 ) & (wr )  ;
assign n16052 =  ( n16051 ) ? ( n4782 ) : ( iram_108 ) ;
assign n16053 = wr_addr[7:7] ;
assign n16054 =  ( n16053 ) == ( bv_1_0_n53 )  ;
assign n16055 =  ( wr_addr ) == ( bv_8_108_n285 )  ;
assign n16056 =  ( n16054 ) & (n16055 )  ;
assign n16057 =  ( n16056 ) & (wr )  ;
assign n16058 =  ( n16057 ) ? ( n4841 ) : ( iram_108 ) ;
assign n16059 = wr_addr[7:7] ;
assign n16060 =  ( n16059 ) == ( bv_1_0_n53 )  ;
assign n16061 =  ( wr_addr ) == ( bv_8_108_n285 )  ;
assign n16062 =  ( n16060 ) & (n16061 )  ;
assign n16063 =  ( n16062 ) & (wr )  ;
assign n16064 =  ( n16063 ) ? ( n5449 ) : ( iram_108 ) ;
assign n16065 = wr_addr[7:7] ;
assign n16066 =  ( n16065 ) == ( bv_1_0_n53 )  ;
assign n16067 =  ( wr_addr ) == ( bv_8_108_n285 )  ;
assign n16068 =  ( n16066 ) & (n16067 )  ;
assign n16069 =  ( n16068 ) & (wr )  ;
assign n16070 =  ( n16069 ) ? ( n4906 ) : ( iram_108 ) ;
assign n16071 = wr_addr[7:7] ;
assign n16072 =  ( n16071 ) == ( bv_1_0_n53 )  ;
assign n16073 =  ( wr_addr ) == ( bv_8_108_n285 )  ;
assign n16074 =  ( n16072 ) & (n16073 )  ;
assign n16075 =  ( n16074 ) & (wr )  ;
assign n16076 =  ( n16075 ) ? ( n5485 ) : ( iram_108 ) ;
assign n16077 = wr_addr[7:7] ;
assign n16078 =  ( n16077 ) == ( bv_1_0_n53 )  ;
assign n16079 =  ( wr_addr ) == ( bv_8_108_n285 )  ;
assign n16080 =  ( n16078 ) & (n16079 )  ;
assign n16081 =  ( n16080 ) & (wr )  ;
assign n16082 =  ( n16081 ) ? ( n5512 ) : ( iram_108 ) ;
assign n16083 = wr_addr[7:7] ;
assign n16084 =  ( n16083 ) == ( bv_1_0_n53 )  ;
assign n16085 =  ( wr_addr ) == ( bv_8_108_n285 )  ;
assign n16086 =  ( n16084 ) & (n16085 )  ;
assign n16087 =  ( n16086 ) & (wr )  ;
assign n16088 =  ( n16087 ) ? ( bv_8_0_n69 ) : ( iram_108 ) ;
assign n16089 = wr_addr[7:7] ;
assign n16090 =  ( n16089 ) == ( bv_1_0_n53 )  ;
assign n16091 =  ( wr_addr ) == ( bv_8_108_n285 )  ;
assign n16092 =  ( n16090 ) & (n16091 )  ;
assign n16093 =  ( n16092 ) & (wr )  ;
assign n16094 =  ( n16093 ) ? ( n5071 ) : ( iram_108 ) ;
assign n16095 = wr_addr[7:7] ;
assign n16096 =  ( n16095 ) == ( bv_1_0_n53 )  ;
assign n16097 =  ( wr_addr ) == ( bv_8_108_n285 )  ;
assign n16098 =  ( n16096 ) & (n16097 )  ;
assign n16099 =  ( n16098 ) & (wr )  ;
assign n16100 =  ( n16099 ) ? ( n5096 ) : ( iram_108 ) ;
assign n16101 = wr_addr[7:7] ;
assign n16102 =  ( n16101 ) == ( bv_1_0_n53 )  ;
assign n16103 =  ( wr_addr ) == ( bv_8_108_n285 )  ;
assign n16104 =  ( n16102 ) & (n16103 )  ;
assign n16105 =  ( n16104 ) & (wr )  ;
assign n16106 =  ( n16105 ) ? ( n5123 ) : ( iram_108 ) ;
assign n16107 = wr_addr[7:7] ;
assign n16108 =  ( n16107 ) == ( bv_1_0_n53 )  ;
assign n16109 =  ( wr_addr ) == ( bv_8_108_n285 )  ;
assign n16110 =  ( n16108 ) & (n16109 )  ;
assign n16111 =  ( n16110 ) & (wr )  ;
assign n16112 =  ( n16111 ) ? ( n5165 ) : ( iram_108 ) ;
assign n16113 = wr_addr[7:7] ;
assign n16114 =  ( n16113 ) == ( bv_1_0_n53 )  ;
assign n16115 =  ( wr_addr ) == ( bv_8_108_n285 )  ;
assign n16116 =  ( n16114 ) & (n16115 )  ;
assign n16117 =  ( n16116 ) & (wr )  ;
assign n16118 =  ( n16117 ) ? ( n5204 ) : ( iram_108 ) ;
assign n16119 = wr_addr[7:7] ;
assign n16120 =  ( n16119 ) == ( bv_1_0_n53 )  ;
assign n16121 =  ( wr_addr ) == ( bv_8_108_n285 )  ;
assign n16122 =  ( n16120 ) & (n16121 )  ;
assign n16123 =  ( n16122 ) & (wr )  ;
assign n16124 =  ( n16123 ) ? ( n5262 ) : ( iram_108 ) ;
assign n16125 = wr_addr[7:7] ;
assign n16126 =  ( n16125 ) == ( bv_1_0_n53 )  ;
assign n16127 =  ( wr_addr ) == ( bv_8_108_n285 )  ;
assign n16128 =  ( n16126 ) & (n16127 )  ;
assign n16129 =  ( n16128 ) & (wr )  ;
assign n16130 =  ( n16129 ) ? ( n5298 ) : ( iram_108 ) ;
assign n16131 = wr_addr[7:7] ;
assign n16132 =  ( n16131 ) == ( bv_1_0_n53 )  ;
assign n16133 =  ( wr_addr ) == ( bv_8_108_n285 )  ;
assign n16134 =  ( n16132 ) & (n16133 )  ;
assign n16135 =  ( n16134 ) & (wr )  ;
assign n16136 =  ( n16135 ) ? ( n5325 ) : ( iram_108 ) ;
assign n16137 = wr_addr[7:7] ;
assign n16138 =  ( n16137 ) == ( bv_1_0_n53 )  ;
assign n16139 =  ( wr_addr ) == ( bv_8_109_n287 )  ;
assign n16140 =  ( n16138 ) & (n16139 )  ;
assign n16141 =  ( n16140 ) & (wr )  ;
assign n16142 =  ( n16141 ) ? ( n4782 ) : ( iram_109 ) ;
assign n16143 = wr_addr[7:7] ;
assign n16144 =  ( n16143 ) == ( bv_1_0_n53 )  ;
assign n16145 =  ( wr_addr ) == ( bv_8_109_n287 )  ;
assign n16146 =  ( n16144 ) & (n16145 )  ;
assign n16147 =  ( n16146 ) & (wr )  ;
assign n16148 =  ( n16147 ) ? ( n4841 ) : ( iram_109 ) ;
assign n16149 = wr_addr[7:7] ;
assign n16150 =  ( n16149 ) == ( bv_1_0_n53 )  ;
assign n16151 =  ( wr_addr ) == ( bv_8_109_n287 )  ;
assign n16152 =  ( n16150 ) & (n16151 )  ;
assign n16153 =  ( n16152 ) & (wr )  ;
assign n16154 =  ( n16153 ) ? ( n5449 ) : ( iram_109 ) ;
assign n16155 = wr_addr[7:7] ;
assign n16156 =  ( n16155 ) == ( bv_1_0_n53 )  ;
assign n16157 =  ( wr_addr ) == ( bv_8_109_n287 )  ;
assign n16158 =  ( n16156 ) & (n16157 )  ;
assign n16159 =  ( n16158 ) & (wr )  ;
assign n16160 =  ( n16159 ) ? ( n4906 ) : ( iram_109 ) ;
assign n16161 = wr_addr[7:7] ;
assign n16162 =  ( n16161 ) == ( bv_1_0_n53 )  ;
assign n16163 =  ( wr_addr ) == ( bv_8_109_n287 )  ;
assign n16164 =  ( n16162 ) & (n16163 )  ;
assign n16165 =  ( n16164 ) & (wr )  ;
assign n16166 =  ( n16165 ) ? ( n5485 ) : ( iram_109 ) ;
assign n16167 = wr_addr[7:7] ;
assign n16168 =  ( n16167 ) == ( bv_1_0_n53 )  ;
assign n16169 =  ( wr_addr ) == ( bv_8_109_n287 )  ;
assign n16170 =  ( n16168 ) & (n16169 )  ;
assign n16171 =  ( n16170 ) & (wr )  ;
assign n16172 =  ( n16171 ) ? ( n5512 ) : ( iram_109 ) ;
assign n16173 = wr_addr[7:7] ;
assign n16174 =  ( n16173 ) == ( bv_1_0_n53 )  ;
assign n16175 =  ( wr_addr ) == ( bv_8_109_n287 )  ;
assign n16176 =  ( n16174 ) & (n16175 )  ;
assign n16177 =  ( n16176 ) & (wr )  ;
assign n16178 =  ( n16177 ) ? ( bv_8_0_n69 ) : ( iram_109 ) ;
assign n16179 = wr_addr[7:7] ;
assign n16180 =  ( n16179 ) == ( bv_1_0_n53 )  ;
assign n16181 =  ( wr_addr ) == ( bv_8_109_n287 )  ;
assign n16182 =  ( n16180 ) & (n16181 )  ;
assign n16183 =  ( n16182 ) & (wr )  ;
assign n16184 =  ( n16183 ) ? ( n5071 ) : ( iram_109 ) ;
assign n16185 = wr_addr[7:7] ;
assign n16186 =  ( n16185 ) == ( bv_1_0_n53 )  ;
assign n16187 =  ( wr_addr ) == ( bv_8_109_n287 )  ;
assign n16188 =  ( n16186 ) & (n16187 )  ;
assign n16189 =  ( n16188 ) & (wr )  ;
assign n16190 =  ( n16189 ) ? ( n5096 ) : ( iram_109 ) ;
assign n16191 = wr_addr[7:7] ;
assign n16192 =  ( n16191 ) == ( bv_1_0_n53 )  ;
assign n16193 =  ( wr_addr ) == ( bv_8_109_n287 )  ;
assign n16194 =  ( n16192 ) & (n16193 )  ;
assign n16195 =  ( n16194 ) & (wr )  ;
assign n16196 =  ( n16195 ) ? ( n5123 ) : ( iram_109 ) ;
assign n16197 = wr_addr[7:7] ;
assign n16198 =  ( n16197 ) == ( bv_1_0_n53 )  ;
assign n16199 =  ( wr_addr ) == ( bv_8_109_n287 )  ;
assign n16200 =  ( n16198 ) & (n16199 )  ;
assign n16201 =  ( n16200 ) & (wr )  ;
assign n16202 =  ( n16201 ) ? ( n5165 ) : ( iram_109 ) ;
assign n16203 = wr_addr[7:7] ;
assign n16204 =  ( n16203 ) == ( bv_1_0_n53 )  ;
assign n16205 =  ( wr_addr ) == ( bv_8_109_n287 )  ;
assign n16206 =  ( n16204 ) & (n16205 )  ;
assign n16207 =  ( n16206 ) & (wr )  ;
assign n16208 =  ( n16207 ) ? ( n5204 ) : ( iram_109 ) ;
assign n16209 = wr_addr[7:7] ;
assign n16210 =  ( n16209 ) == ( bv_1_0_n53 )  ;
assign n16211 =  ( wr_addr ) == ( bv_8_109_n287 )  ;
assign n16212 =  ( n16210 ) & (n16211 )  ;
assign n16213 =  ( n16212 ) & (wr )  ;
assign n16214 =  ( n16213 ) ? ( n5262 ) : ( iram_109 ) ;
assign n16215 = wr_addr[7:7] ;
assign n16216 =  ( n16215 ) == ( bv_1_0_n53 )  ;
assign n16217 =  ( wr_addr ) == ( bv_8_109_n287 )  ;
assign n16218 =  ( n16216 ) & (n16217 )  ;
assign n16219 =  ( n16218 ) & (wr )  ;
assign n16220 =  ( n16219 ) ? ( n5298 ) : ( iram_109 ) ;
assign n16221 = wr_addr[7:7] ;
assign n16222 =  ( n16221 ) == ( bv_1_0_n53 )  ;
assign n16223 =  ( wr_addr ) == ( bv_8_109_n287 )  ;
assign n16224 =  ( n16222 ) & (n16223 )  ;
assign n16225 =  ( n16224 ) & (wr )  ;
assign n16226 =  ( n16225 ) ? ( n5325 ) : ( iram_109 ) ;
assign n16227 = wr_addr[7:7] ;
assign n16228 =  ( n16227 ) == ( bv_1_0_n53 )  ;
assign n16229 =  ( wr_addr ) == ( bv_8_110_n289 )  ;
assign n16230 =  ( n16228 ) & (n16229 )  ;
assign n16231 =  ( n16230 ) & (wr )  ;
assign n16232 =  ( n16231 ) ? ( n4782 ) : ( iram_110 ) ;
assign n16233 = wr_addr[7:7] ;
assign n16234 =  ( n16233 ) == ( bv_1_0_n53 )  ;
assign n16235 =  ( wr_addr ) == ( bv_8_110_n289 )  ;
assign n16236 =  ( n16234 ) & (n16235 )  ;
assign n16237 =  ( n16236 ) & (wr )  ;
assign n16238 =  ( n16237 ) ? ( n4841 ) : ( iram_110 ) ;
assign n16239 = wr_addr[7:7] ;
assign n16240 =  ( n16239 ) == ( bv_1_0_n53 )  ;
assign n16241 =  ( wr_addr ) == ( bv_8_110_n289 )  ;
assign n16242 =  ( n16240 ) & (n16241 )  ;
assign n16243 =  ( n16242 ) & (wr )  ;
assign n16244 =  ( n16243 ) ? ( n5449 ) : ( iram_110 ) ;
assign n16245 = wr_addr[7:7] ;
assign n16246 =  ( n16245 ) == ( bv_1_0_n53 )  ;
assign n16247 =  ( wr_addr ) == ( bv_8_110_n289 )  ;
assign n16248 =  ( n16246 ) & (n16247 )  ;
assign n16249 =  ( n16248 ) & (wr )  ;
assign n16250 =  ( n16249 ) ? ( n4906 ) : ( iram_110 ) ;
assign n16251 = wr_addr[7:7] ;
assign n16252 =  ( n16251 ) == ( bv_1_0_n53 )  ;
assign n16253 =  ( wr_addr ) == ( bv_8_110_n289 )  ;
assign n16254 =  ( n16252 ) & (n16253 )  ;
assign n16255 =  ( n16254 ) & (wr )  ;
assign n16256 =  ( n16255 ) ? ( n5485 ) : ( iram_110 ) ;
assign n16257 = wr_addr[7:7] ;
assign n16258 =  ( n16257 ) == ( bv_1_0_n53 )  ;
assign n16259 =  ( wr_addr ) == ( bv_8_110_n289 )  ;
assign n16260 =  ( n16258 ) & (n16259 )  ;
assign n16261 =  ( n16260 ) & (wr )  ;
assign n16262 =  ( n16261 ) ? ( n5512 ) : ( iram_110 ) ;
assign n16263 = wr_addr[7:7] ;
assign n16264 =  ( n16263 ) == ( bv_1_0_n53 )  ;
assign n16265 =  ( wr_addr ) == ( bv_8_110_n289 )  ;
assign n16266 =  ( n16264 ) & (n16265 )  ;
assign n16267 =  ( n16266 ) & (wr )  ;
assign n16268 =  ( n16267 ) ? ( bv_8_0_n69 ) : ( iram_110 ) ;
assign n16269 = wr_addr[7:7] ;
assign n16270 =  ( n16269 ) == ( bv_1_0_n53 )  ;
assign n16271 =  ( wr_addr ) == ( bv_8_110_n289 )  ;
assign n16272 =  ( n16270 ) & (n16271 )  ;
assign n16273 =  ( n16272 ) & (wr )  ;
assign n16274 =  ( n16273 ) ? ( n5071 ) : ( iram_110 ) ;
assign n16275 = wr_addr[7:7] ;
assign n16276 =  ( n16275 ) == ( bv_1_0_n53 )  ;
assign n16277 =  ( wr_addr ) == ( bv_8_110_n289 )  ;
assign n16278 =  ( n16276 ) & (n16277 )  ;
assign n16279 =  ( n16278 ) & (wr )  ;
assign n16280 =  ( n16279 ) ? ( n5096 ) : ( iram_110 ) ;
assign n16281 = wr_addr[7:7] ;
assign n16282 =  ( n16281 ) == ( bv_1_0_n53 )  ;
assign n16283 =  ( wr_addr ) == ( bv_8_110_n289 )  ;
assign n16284 =  ( n16282 ) & (n16283 )  ;
assign n16285 =  ( n16284 ) & (wr )  ;
assign n16286 =  ( n16285 ) ? ( n5123 ) : ( iram_110 ) ;
assign n16287 = wr_addr[7:7] ;
assign n16288 =  ( n16287 ) == ( bv_1_0_n53 )  ;
assign n16289 =  ( wr_addr ) == ( bv_8_110_n289 )  ;
assign n16290 =  ( n16288 ) & (n16289 )  ;
assign n16291 =  ( n16290 ) & (wr )  ;
assign n16292 =  ( n16291 ) ? ( n5165 ) : ( iram_110 ) ;
assign n16293 = wr_addr[7:7] ;
assign n16294 =  ( n16293 ) == ( bv_1_0_n53 )  ;
assign n16295 =  ( wr_addr ) == ( bv_8_110_n289 )  ;
assign n16296 =  ( n16294 ) & (n16295 )  ;
assign n16297 =  ( n16296 ) & (wr )  ;
assign n16298 =  ( n16297 ) ? ( n5204 ) : ( iram_110 ) ;
assign n16299 = wr_addr[7:7] ;
assign n16300 =  ( n16299 ) == ( bv_1_0_n53 )  ;
assign n16301 =  ( wr_addr ) == ( bv_8_110_n289 )  ;
assign n16302 =  ( n16300 ) & (n16301 )  ;
assign n16303 =  ( n16302 ) & (wr )  ;
assign n16304 =  ( n16303 ) ? ( n5262 ) : ( iram_110 ) ;
assign n16305 = wr_addr[7:7] ;
assign n16306 =  ( n16305 ) == ( bv_1_0_n53 )  ;
assign n16307 =  ( wr_addr ) == ( bv_8_110_n289 )  ;
assign n16308 =  ( n16306 ) & (n16307 )  ;
assign n16309 =  ( n16308 ) & (wr )  ;
assign n16310 =  ( n16309 ) ? ( n5298 ) : ( iram_110 ) ;
assign n16311 = wr_addr[7:7] ;
assign n16312 =  ( n16311 ) == ( bv_1_0_n53 )  ;
assign n16313 =  ( wr_addr ) == ( bv_8_110_n289 )  ;
assign n16314 =  ( n16312 ) & (n16313 )  ;
assign n16315 =  ( n16314 ) & (wr )  ;
assign n16316 =  ( n16315 ) ? ( n5325 ) : ( iram_110 ) ;
assign n16317 = wr_addr[7:7] ;
assign n16318 =  ( n16317 ) == ( bv_1_0_n53 )  ;
assign n16319 =  ( wr_addr ) == ( bv_8_111_n291 )  ;
assign n16320 =  ( n16318 ) & (n16319 )  ;
assign n16321 =  ( n16320 ) & (wr )  ;
assign n16322 =  ( n16321 ) ? ( n4782 ) : ( iram_111 ) ;
assign n16323 = wr_addr[7:7] ;
assign n16324 =  ( n16323 ) == ( bv_1_0_n53 )  ;
assign n16325 =  ( wr_addr ) == ( bv_8_111_n291 )  ;
assign n16326 =  ( n16324 ) & (n16325 )  ;
assign n16327 =  ( n16326 ) & (wr )  ;
assign n16328 =  ( n16327 ) ? ( n4841 ) : ( iram_111 ) ;
assign n16329 = wr_addr[7:7] ;
assign n16330 =  ( n16329 ) == ( bv_1_0_n53 )  ;
assign n16331 =  ( wr_addr ) == ( bv_8_111_n291 )  ;
assign n16332 =  ( n16330 ) & (n16331 )  ;
assign n16333 =  ( n16332 ) & (wr )  ;
assign n16334 =  ( n16333 ) ? ( n5449 ) : ( iram_111 ) ;
assign n16335 = wr_addr[7:7] ;
assign n16336 =  ( n16335 ) == ( bv_1_0_n53 )  ;
assign n16337 =  ( wr_addr ) == ( bv_8_111_n291 )  ;
assign n16338 =  ( n16336 ) & (n16337 )  ;
assign n16339 =  ( n16338 ) & (wr )  ;
assign n16340 =  ( n16339 ) ? ( n4906 ) : ( iram_111 ) ;
assign n16341 = wr_addr[7:7] ;
assign n16342 =  ( n16341 ) == ( bv_1_0_n53 )  ;
assign n16343 =  ( wr_addr ) == ( bv_8_111_n291 )  ;
assign n16344 =  ( n16342 ) & (n16343 )  ;
assign n16345 =  ( n16344 ) & (wr )  ;
assign n16346 =  ( n16345 ) ? ( n5485 ) : ( iram_111 ) ;
assign n16347 = wr_addr[7:7] ;
assign n16348 =  ( n16347 ) == ( bv_1_0_n53 )  ;
assign n16349 =  ( wr_addr ) == ( bv_8_111_n291 )  ;
assign n16350 =  ( n16348 ) & (n16349 )  ;
assign n16351 =  ( n16350 ) & (wr )  ;
assign n16352 =  ( n16351 ) ? ( n5512 ) : ( iram_111 ) ;
assign n16353 = wr_addr[7:7] ;
assign n16354 =  ( n16353 ) == ( bv_1_0_n53 )  ;
assign n16355 =  ( wr_addr ) == ( bv_8_111_n291 )  ;
assign n16356 =  ( n16354 ) & (n16355 )  ;
assign n16357 =  ( n16356 ) & (wr )  ;
assign n16358 =  ( n16357 ) ? ( bv_8_0_n69 ) : ( iram_111 ) ;
assign n16359 = wr_addr[7:7] ;
assign n16360 =  ( n16359 ) == ( bv_1_0_n53 )  ;
assign n16361 =  ( wr_addr ) == ( bv_8_111_n291 )  ;
assign n16362 =  ( n16360 ) & (n16361 )  ;
assign n16363 =  ( n16362 ) & (wr )  ;
assign n16364 =  ( n16363 ) ? ( n5071 ) : ( iram_111 ) ;
assign n16365 = wr_addr[7:7] ;
assign n16366 =  ( n16365 ) == ( bv_1_0_n53 )  ;
assign n16367 =  ( wr_addr ) == ( bv_8_111_n291 )  ;
assign n16368 =  ( n16366 ) & (n16367 )  ;
assign n16369 =  ( n16368 ) & (wr )  ;
assign n16370 =  ( n16369 ) ? ( n5096 ) : ( iram_111 ) ;
assign n16371 = wr_addr[7:7] ;
assign n16372 =  ( n16371 ) == ( bv_1_0_n53 )  ;
assign n16373 =  ( wr_addr ) == ( bv_8_111_n291 )  ;
assign n16374 =  ( n16372 ) & (n16373 )  ;
assign n16375 =  ( n16374 ) & (wr )  ;
assign n16376 =  ( n16375 ) ? ( n5123 ) : ( iram_111 ) ;
assign n16377 = wr_addr[7:7] ;
assign n16378 =  ( n16377 ) == ( bv_1_0_n53 )  ;
assign n16379 =  ( wr_addr ) == ( bv_8_111_n291 )  ;
assign n16380 =  ( n16378 ) & (n16379 )  ;
assign n16381 =  ( n16380 ) & (wr )  ;
assign n16382 =  ( n16381 ) ? ( n5165 ) : ( iram_111 ) ;
assign n16383 = wr_addr[7:7] ;
assign n16384 =  ( n16383 ) == ( bv_1_0_n53 )  ;
assign n16385 =  ( wr_addr ) == ( bv_8_111_n291 )  ;
assign n16386 =  ( n16384 ) & (n16385 )  ;
assign n16387 =  ( n16386 ) & (wr )  ;
assign n16388 =  ( n16387 ) ? ( n5204 ) : ( iram_111 ) ;
assign n16389 = wr_addr[7:7] ;
assign n16390 =  ( n16389 ) == ( bv_1_0_n53 )  ;
assign n16391 =  ( wr_addr ) == ( bv_8_111_n291 )  ;
assign n16392 =  ( n16390 ) & (n16391 )  ;
assign n16393 =  ( n16392 ) & (wr )  ;
assign n16394 =  ( n16393 ) ? ( n5262 ) : ( iram_111 ) ;
assign n16395 = wr_addr[7:7] ;
assign n16396 =  ( n16395 ) == ( bv_1_0_n53 )  ;
assign n16397 =  ( wr_addr ) == ( bv_8_111_n291 )  ;
assign n16398 =  ( n16396 ) & (n16397 )  ;
assign n16399 =  ( n16398 ) & (wr )  ;
assign n16400 =  ( n16399 ) ? ( n5298 ) : ( iram_111 ) ;
assign n16401 = wr_addr[7:7] ;
assign n16402 =  ( n16401 ) == ( bv_1_0_n53 )  ;
assign n16403 =  ( wr_addr ) == ( bv_8_111_n291 )  ;
assign n16404 =  ( n16402 ) & (n16403 )  ;
assign n16405 =  ( n16404 ) & (wr )  ;
assign n16406 =  ( n16405 ) ? ( n5325 ) : ( iram_111 ) ;
assign n16407 = wr_addr[7:7] ;
assign n16408 =  ( n16407 ) == ( bv_1_0_n53 )  ;
assign n16409 =  ( wr_addr ) == ( bv_8_112_n293 )  ;
assign n16410 =  ( n16408 ) & (n16409 )  ;
assign n16411 =  ( n16410 ) & (wr )  ;
assign n16412 =  ( n16411 ) ? ( n4782 ) : ( iram_112 ) ;
assign n16413 = wr_addr[7:7] ;
assign n16414 =  ( n16413 ) == ( bv_1_0_n53 )  ;
assign n16415 =  ( wr_addr ) == ( bv_8_112_n293 )  ;
assign n16416 =  ( n16414 ) & (n16415 )  ;
assign n16417 =  ( n16416 ) & (wr )  ;
assign n16418 =  ( n16417 ) ? ( n4841 ) : ( iram_112 ) ;
assign n16419 = wr_addr[7:7] ;
assign n16420 =  ( n16419 ) == ( bv_1_0_n53 )  ;
assign n16421 =  ( wr_addr ) == ( bv_8_112_n293 )  ;
assign n16422 =  ( n16420 ) & (n16421 )  ;
assign n16423 =  ( n16422 ) & (wr )  ;
assign n16424 =  ( n16423 ) ? ( n5449 ) : ( iram_112 ) ;
assign n16425 = wr_addr[7:7] ;
assign n16426 =  ( n16425 ) == ( bv_1_0_n53 )  ;
assign n16427 =  ( wr_addr ) == ( bv_8_112_n293 )  ;
assign n16428 =  ( n16426 ) & (n16427 )  ;
assign n16429 =  ( n16428 ) & (wr )  ;
assign n16430 =  ( n16429 ) ? ( n4906 ) : ( iram_112 ) ;
assign n16431 = wr_addr[7:7] ;
assign n16432 =  ( n16431 ) == ( bv_1_0_n53 )  ;
assign n16433 =  ( wr_addr ) == ( bv_8_112_n293 )  ;
assign n16434 =  ( n16432 ) & (n16433 )  ;
assign n16435 =  ( n16434 ) & (wr )  ;
assign n16436 =  ( n16435 ) ? ( n5485 ) : ( iram_112 ) ;
assign n16437 = wr_addr[7:7] ;
assign n16438 =  ( n16437 ) == ( bv_1_0_n53 )  ;
assign n16439 =  ( wr_addr ) == ( bv_8_112_n293 )  ;
assign n16440 =  ( n16438 ) & (n16439 )  ;
assign n16441 =  ( n16440 ) & (wr )  ;
assign n16442 =  ( n16441 ) ? ( n5512 ) : ( iram_112 ) ;
assign n16443 = wr_addr[7:7] ;
assign n16444 =  ( n16443 ) == ( bv_1_0_n53 )  ;
assign n16445 =  ( wr_addr ) == ( bv_8_112_n293 )  ;
assign n16446 =  ( n16444 ) & (n16445 )  ;
assign n16447 =  ( n16446 ) & (wr )  ;
assign n16448 =  ( n16447 ) ? ( bv_8_0_n69 ) : ( iram_112 ) ;
assign n16449 = wr_addr[7:7] ;
assign n16450 =  ( n16449 ) == ( bv_1_0_n53 )  ;
assign n16451 =  ( wr_addr ) == ( bv_8_112_n293 )  ;
assign n16452 =  ( n16450 ) & (n16451 )  ;
assign n16453 =  ( n16452 ) & (wr )  ;
assign n16454 =  ( n16453 ) ? ( n5071 ) : ( iram_112 ) ;
assign n16455 = wr_addr[7:7] ;
assign n16456 =  ( n16455 ) == ( bv_1_0_n53 )  ;
assign n16457 =  ( wr_addr ) == ( bv_8_112_n293 )  ;
assign n16458 =  ( n16456 ) & (n16457 )  ;
assign n16459 =  ( n16458 ) & (wr )  ;
assign n16460 =  ( n16459 ) ? ( n5096 ) : ( iram_112 ) ;
assign n16461 = wr_addr[7:7] ;
assign n16462 =  ( n16461 ) == ( bv_1_0_n53 )  ;
assign n16463 =  ( wr_addr ) == ( bv_8_112_n293 )  ;
assign n16464 =  ( n16462 ) & (n16463 )  ;
assign n16465 =  ( n16464 ) & (wr )  ;
assign n16466 =  ( n16465 ) ? ( n5123 ) : ( iram_112 ) ;
assign n16467 = wr_addr[7:7] ;
assign n16468 =  ( n16467 ) == ( bv_1_0_n53 )  ;
assign n16469 =  ( wr_addr ) == ( bv_8_112_n293 )  ;
assign n16470 =  ( n16468 ) & (n16469 )  ;
assign n16471 =  ( n16470 ) & (wr )  ;
assign n16472 =  ( n16471 ) ? ( n5165 ) : ( iram_112 ) ;
assign n16473 = wr_addr[7:7] ;
assign n16474 =  ( n16473 ) == ( bv_1_0_n53 )  ;
assign n16475 =  ( wr_addr ) == ( bv_8_112_n293 )  ;
assign n16476 =  ( n16474 ) & (n16475 )  ;
assign n16477 =  ( n16476 ) & (wr )  ;
assign n16478 =  ( n16477 ) ? ( n5204 ) : ( iram_112 ) ;
assign n16479 = wr_addr[7:7] ;
assign n16480 =  ( n16479 ) == ( bv_1_0_n53 )  ;
assign n16481 =  ( wr_addr ) == ( bv_8_112_n293 )  ;
assign n16482 =  ( n16480 ) & (n16481 )  ;
assign n16483 =  ( n16482 ) & (wr )  ;
assign n16484 =  ( n16483 ) ? ( n5262 ) : ( iram_112 ) ;
assign n16485 = wr_addr[7:7] ;
assign n16486 =  ( n16485 ) == ( bv_1_0_n53 )  ;
assign n16487 =  ( wr_addr ) == ( bv_8_112_n293 )  ;
assign n16488 =  ( n16486 ) & (n16487 )  ;
assign n16489 =  ( n16488 ) & (wr )  ;
assign n16490 =  ( n16489 ) ? ( n5298 ) : ( iram_112 ) ;
assign n16491 = wr_addr[7:7] ;
assign n16492 =  ( n16491 ) == ( bv_1_0_n53 )  ;
assign n16493 =  ( wr_addr ) == ( bv_8_112_n293 )  ;
assign n16494 =  ( n16492 ) & (n16493 )  ;
assign n16495 =  ( n16494 ) & (wr )  ;
assign n16496 =  ( n16495 ) ? ( n5325 ) : ( iram_112 ) ;
assign n16497 = wr_addr[7:7] ;
assign n16498 =  ( n16497 ) == ( bv_1_0_n53 )  ;
assign n16499 =  ( wr_addr ) == ( bv_8_113_n295 )  ;
assign n16500 =  ( n16498 ) & (n16499 )  ;
assign n16501 =  ( n16500 ) & (wr )  ;
assign n16502 =  ( n16501 ) ? ( n4782 ) : ( iram_113 ) ;
assign n16503 = wr_addr[7:7] ;
assign n16504 =  ( n16503 ) == ( bv_1_0_n53 )  ;
assign n16505 =  ( wr_addr ) == ( bv_8_113_n295 )  ;
assign n16506 =  ( n16504 ) & (n16505 )  ;
assign n16507 =  ( n16506 ) & (wr )  ;
assign n16508 =  ( n16507 ) ? ( n4841 ) : ( iram_113 ) ;
assign n16509 = wr_addr[7:7] ;
assign n16510 =  ( n16509 ) == ( bv_1_0_n53 )  ;
assign n16511 =  ( wr_addr ) == ( bv_8_113_n295 )  ;
assign n16512 =  ( n16510 ) & (n16511 )  ;
assign n16513 =  ( n16512 ) & (wr )  ;
assign n16514 =  ( n16513 ) ? ( n5449 ) : ( iram_113 ) ;
assign n16515 = wr_addr[7:7] ;
assign n16516 =  ( n16515 ) == ( bv_1_0_n53 )  ;
assign n16517 =  ( wr_addr ) == ( bv_8_113_n295 )  ;
assign n16518 =  ( n16516 ) & (n16517 )  ;
assign n16519 =  ( n16518 ) & (wr )  ;
assign n16520 =  ( n16519 ) ? ( n4906 ) : ( iram_113 ) ;
assign n16521 = wr_addr[7:7] ;
assign n16522 =  ( n16521 ) == ( bv_1_0_n53 )  ;
assign n16523 =  ( wr_addr ) == ( bv_8_113_n295 )  ;
assign n16524 =  ( n16522 ) & (n16523 )  ;
assign n16525 =  ( n16524 ) & (wr )  ;
assign n16526 =  ( n16525 ) ? ( n5485 ) : ( iram_113 ) ;
assign n16527 = wr_addr[7:7] ;
assign n16528 =  ( n16527 ) == ( bv_1_0_n53 )  ;
assign n16529 =  ( wr_addr ) == ( bv_8_113_n295 )  ;
assign n16530 =  ( n16528 ) & (n16529 )  ;
assign n16531 =  ( n16530 ) & (wr )  ;
assign n16532 =  ( n16531 ) ? ( n5512 ) : ( iram_113 ) ;
assign n16533 = wr_addr[7:7] ;
assign n16534 =  ( n16533 ) == ( bv_1_0_n53 )  ;
assign n16535 =  ( wr_addr ) == ( bv_8_113_n295 )  ;
assign n16536 =  ( n16534 ) & (n16535 )  ;
assign n16537 =  ( n16536 ) & (wr )  ;
assign n16538 =  ( n16537 ) ? ( bv_8_0_n69 ) : ( iram_113 ) ;
assign n16539 = wr_addr[7:7] ;
assign n16540 =  ( n16539 ) == ( bv_1_0_n53 )  ;
assign n16541 =  ( wr_addr ) == ( bv_8_113_n295 )  ;
assign n16542 =  ( n16540 ) & (n16541 )  ;
assign n16543 =  ( n16542 ) & (wr )  ;
assign n16544 =  ( n16543 ) ? ( n5071 ) : ( iram_113 ) ;
assign n16545 = wr_addr[7:7] ;
assign n16546 =  ( n16545 ) == ( bv_1_0_n53 )  ;
assign n16547 =  ( wr_addr ) == ( bv_8_113_n295 )  ;
assign n16548 =  ( n16546 ) & (n16547 )  ;
assign n16549 =  ( n16548 ) & (wr )  ;
assign n16550 =  ( n16549 ) ? ( n5096 ) : ( iram_113 ) ;
assign n16551 = wr_addr[7:7] ;
assign n16552 =  ( n16551 ) == ( bv_1_0_n53 )  ;
assign n16553 =  ( wr_addr ) == ( bv_8_113_n295 )  ;
assign n16554 =  ( n16552 ) & (n16553 )  ;
assign n16555 =  ( n16554 ) & (wr )  ;
assign n16556 =  ( n16555 ) ? ( n5123 ) : ( iram_113 ) ;
assign n16557 = wr_addr[7:7] ;
assign n16558 =  ( n16557 ) == ( bv_1_0_n53 )  ;
assign n16559 =  ( wr_addr ) == ( bv_8_113_n295 )  ;
assign n16560 =  ( n16558 ) & (n16559 )  ;
assign n16561 =  ( n16560 ) & (wr )  ;
assign n16562 =  ( n16561 ) ? ( n5165 ) : ( iram_113 ) ;
assign n16563 = wr_addr[7:7] ;
assign n16564 =  ( n16563 ) == ( bv_1_0_n53 )  ;
assign n16565 =  ( wr_addr ) == ( bv_8_113_n295 )  ;
assign n16566 =  ( n16564 ) & (n16565 )  ;
assign n16567 =  ( n16566 ) & (wr )  ;
assign n16568 =  ( n16567 ) ? ( n5204 ) : ( iram_113 ) ;
assign n16569 = wr_addr[7:7] ;
assign n16570 =  ( n16569 ) == ( bv_1_0_n53 )  ;
assign n16571 =  ( wr_addr ) == ( bv_8_113_n295 )  ;
assign n16572 =  ( n16570 ) & (n16571 )  ;
assign n16573 =  ( n16572 ) & (wr )  ;
assign n16574 =  ( n16573 ) ? ( n5262 ) : ( iram_113 ) ;
assign n16575 = wr_addr[7:7] ;
assign n16576 =  ( n16575 ) == ( bv_1_0_n53 )  ;
assign n16577 =  ( wr_addr ) == ( bv_8_113_n295 )  ;
assign n16578 =  ( n16576 ) & (n16577 )  ;
assign n16579 =  ( n16578 ) & (wr )  ;
assign n16580 =  ( n16579 ) ? ( n5298 ) : ( iram_113 ) ;
assign n16581 = wr_addr[7:7] ;
assign n16582 =  ( n16581 ) == ( bv_1_0_n53 )  ;
assign n16583 =  ( wr_addr ) == ( bv_8_113_n295 )  ;
assign n16584 =  ( n16582 ) & (n16583 )  ;
assign n16585 =  ( n16584 ) & (wr )  ;
assign n16586 =  ( n16585 ) ? ( n5325 ) : ( iram_113 ) ;
assign n16587 = wr_addr[7:7] ;
assign n16588 =  ( n16587 ) == ( bv_1_0_n53 )  ;
assign n16589 =  ( wr_addr ) == ( bv_8_114_n297 )  ;
assign n16590 =  ( n16588 ) & (n16589 )  ;
assign n16591 =  ( n16590 ) & (wr )  ;
assign n16592 =  ( n16591 ) ? ( n4782 ) : ( iram_114 ) ;
assign n16593 = wr_addr[7:7] ;
assign n16594 =  ( n16593 ) == ( bv_1_0_n53 )  ;
assign n16595 =  ( wr_addr ) == ( bv_8_114_n297 )  ;
assign n16596 =  ( n16594 ) & (n16595 )  ;
assign n16597 =  ( n16596 ) & (wr )  ;
assign n16598 =  ( n16597 ) ? ( n4841 ) : ( iram_114 ) ;
assign n16599 = wr_addr[7:7] ;
assign n16600 =  ( n16599 ) == ( bv_1_0_n53 )  ;
assign n16601 =  ( wr_addr ) == ( bv_8_114_n297 )  ;
assign n16602 =  ( n16600 ) & (n16601 )  ;
assign n16603 =  ( n16602 ) & (wr )  ;
assign n16604 =  ( n16603 ) ? ( n5449 ) : ( iram_114 ) ;
assign n16605 = wr_addr[7:7] ;
assign n16606 =  ( n16605 ) == ( bv_1_0_n53 )  ;
assign n16607 =  ( wr_addr ) == ( bv_8_114_n297 )  ;
assign n16608 =  ( n16606 ) & (n16607 )  ;
assign n16609 =  ( n16608 ) & (wr )  ;
assign n16610 =  ( n16609 ) ? ( n4906 ) : ( iram_114 ) ;
assign n16611 = wr_addr[7:7] ;
assign n16612 =  ( n16611 ) == ( bv_1_0_n53 )  ;
assign n16613 =  ( wr_addr ) == ( bv_8_114_n297 )  ;
assign n16614 =  ( n16612 ) & (n16613 )  ;
assign n16615 =  ( n16614 ) & (wr )  ;
assign n16616 =  ( n16615 ) ? ( n5485 ) : ( iram_114 ) ;
assign n16617 = wr_addr[7:7] ;
assign n16618 =  ( n16617 ) == ( bv_1_0_n53 )  ;
assign n16619 =  ( wr_addr ) == ( bv_8_114_n297 )  ;
assign n16620 =  ( n16618 ) & (n16619 )  ;
assign n16621 =  ( n16620 ) & (wr )  ;
assign n16622 =  ( n16621 ) ? ( n5512 ) : ( iram_114 ) ;
assign n16623 = wr_addr[7:7] ;
assign n16624 =  ( n16623 ) == ( bv_1_0_n53 )  ;
assign n16625 =  ( wr_addr ) == ( bv_8_114_n297 )  ;
assign n16626 =  ( n16624 ) & (n16625 )  ;
assign n16627 =  ( n16626 ) & (wr )  ;
assign n16628 =  ( n16627 ) ? ( bv_8_0_n69 ) : ( iram_114 ) ;
assign n16629 = wr_addr[7:7] ;
assign n16630 =  ( n16629 ) == ( bv_1_0_n53 )  ;
assign n16631 =  ( wr_addr ) == ( bv_8_114_n297 )  ;
assign n16632 =  ( n16630 ) & (n16631 )  ;
assign n16633 =  ( n16632 ) & (wr )  ;
assign n16634 =  ( n16633 ) ? ( n5071 ) : ( iram_114 ) ;
assign n16635 = wr_addr[7:7] ;
assign n16636 =  ( n16635 ) == ( bv_1_0_n53 )  ;
assign n16637 =  ( wr_addr ) == ( bv_8_114_n297 )  ;
assign n16638 =  ( n16636 ) & (n16637 )  ;
assign n16639 =  ( n16638 ) & (wr )  ;
assign n16640 =  ( n16639 ) ? ( n5096 ) : ( iram_114 ) ;
assign n16641 = wr_addr[7:7] ;
assign n16642 =  ( n16641 ) == ( bv_1_0_n53 )  ;
assign n16643 =  ( wr_addr ) == ( bv_8_114_n297 )  ;
assign n16644 =  ( n16642 ) & (n16643 )  ;
assign n16645 =  ( n16644 ) & (wr )  ;
assign n16646 =  ( n16645 ) ? ( n5123 ) : ( iram_114 ) ;
assign n16647 = wr_addr[7:7] ;
assign n16648 =  ( n16647 ) == ( bv_1_0_n53 )  ;
assign n16649 =  ( wr_addr ) == ( bv_8_114_n297 )  ;
assign n16650 =  ( n16648 ) & (n16649 )  ;
assign n16651 =  ( n16650 ) & (wr )  ;
assign n16652 =  ( n16651 ) ? ( n5165 ) : ( iram_114 ) ;
assign n16653 = wr_addr[7:7] ;
assign n16654 =  ( n16653 ) == ( bv_1_0_n53 )  ;
assign n16655 =  ( wr_addr ) == ( bv_8_114_n297 )  ;
assign n16656 =  ( n16654 ) & (n16655 )  ;
assign n16657 =  ( n16656 ) & (wr )  ;
assign n16658 =  ( n16657 ) ? ( n5204 ) : ( iram_114 ) ;
assign n16659 = wr_addr[7:7] ;
assign n16660 =  ( n16659 ) == ( bv_1_0_n53 )  ;
assign n16661 =  ( wr_addr ) == ( bv_8_114_n297 )  ;
assign n16662 =  ( n16660 ) & (n16661 )  ;
assign n16663 =  ( n16662 ) & (wr )  ;
assign n16664 =  ( n16663 ) ? ( n5262 ) : ( iram_114 ) ;
assign n16665 = wr_addr[7:7] ;
assign n16666 =  ( n16665 ) == ( bv_1_0_n53 )  ;
assign n16667 =  ( wr_addr ) == ( bv_8_114_n297 )  ;
assign n16668 =  ( n16666 ) & (n16667 )  ;
assign n16669 =  ( n16668 ) & (wr )  ;
assign n16670 =  ( n16669 ) ? ( n5298 ) : ( iram_114 ) ;
assign n16671 = wr_addr[7:7] ;
assign n16672 =  ( n16671 ) == ( bv_1_0_n53 )  ;
assign n16673 =  ( wr_addr ) == ( bv_8_114_n297 )  ;
assign n16674 =  ( n16672 ) & (n16673 )  ;
assign n16675 =  ( n16674 ) & (wr )  ;
assign n16676 =  ( n16675 ) ? ( n5325 ) : ( iram_114 ) ;
assign n16677 = wr_addr[7:7] ;
assign n16678 =  ( n16677 ) == ( bv_1_0_n53 )  ;
assign n16679 =  ( wr_addr ) == ( bv_8_115_n299 )  ;
assign n16680 =  ( n16678 ) & (n16679 )  ;
assign n16681 =  ( n16680 ) & (wr )  ;
assign n16682 =  ( n16681 ) ? ( n4782 ) : ( iram_115 ) ;
assign n16683 = wr_addr[7:7] ;
assign n16684 =  ( n16683 ) == ( bv_1_0_n53 )  ;
assign n16685 =  ( wr_addr ) == ( bv_8_115_n299 )  ;
assign n16686 =  ( n16684 ) & (n16685 )  ;
assign n16687 =  ( n16686 ) & (wr )  ;
assign n16688 =  ( n16687 ) ? ( n4841 ) : ( iram_115 ) ;
assign n16689 = wr_addr[7:7] ;
assign n16690 =  ( n16689 ) == ( bv_1_0_n53 )  ;
assign n16691 =  ( wr_addr ) == ( bv_8_115_n299 )  ;
assign n16692 =  ( n16690 ) & (n16691 )  ;
assign n16693 =  ( n16692 ) & (wr )  ;
assign n16694 =  ( n16693 ) ? ( n5449 ) : ( iram_115 ) ;
assign n16695 = wr_addr[7:7] ;
assign n16696 =  ( n16695 ) == ( bv_1_0_n53 )  ;
assign n16697 =  ( wr_addr ) == ( bv_8_115_n299 )  ;
assign n16698 =  ( n16696 ) & (n16697 )  ;
assign n16699 =  ( n16698 ) & (wr )  ;
assign n16700 =  ( n16699 ) ? ( n4906 ) : ( iram_115 ) ;
assign n16701 = wr_addr[7:7] ;
assign n16702 =  ( n16701 ) == ( bv_1_0_n53 )  ;
assign n16703 =  ( wr_addr ) == ( bv_8_115_n299 )  ;
assign n16704 =  ( n16702 ) & (n16703 )  ;
assign n16705 =  ( n16704 ) & (wr )  ;
assign n16706 =  ( n16705 ) ? ( n5485 ) : ( iram_115 ) ;
assign n16707 = wr_addr[7:7] ;
assign n16708 =  ( n16707 ) == ( bv_1_0_n53 )  ;
assign n16709 =  ( wr_addr ) == ( bv_8_115_n299 )  ;
assign n16710 =  ( n16708 ) & (n16709 )  ;
assign n16711 =  ( n16710 ) & (wr )  ;
assign n16712 =  ( n16711 ) ? ( n5512 ) : ( iram_115 ) ;
assign n16713 = wr_addr[7:7] ;
assign n16714 =  ( n16713 ) == ( bv_1_0_n53 )  ;
assign n16715 =  ( wr_addr ) == ( bv_8_115_n299 )  ;
assign n16716 =  ( n16714 ) & (n16715 )  ;
assign n16717 =  ( n16716 ) & (wr )  ;
assign n16718 =  ( n16717 ) ? ( bv_8_0_n69 ) : ( iram_115 ) ;
assign n16719 = wr_addr[7:7] ;
assign n16720 =  ( n16719 ) == ( bv_1_0_n53 )  ;
assign n16721 =  ( wr_addr ) == ( bv_8_115_n299 )  ;
assign n16722 =  ( n16720 ) & (n16721 )  ;
assign n16723 =  ( n16722 ) & (wr )  ;
assign n16724 =  ( n16723 ) ? ( n5071 ) : ( iram_115 ) ;
assign n16725 = wr_addr[7:7] ;
assign n16726 =  ( n16725 ) == ( bv_1_0_n53 )  ;
assign n16727 =  ( wr_addr ) == ( bv_8_115_n299 )  ;
assign n16728 =  ( n16726 ) & (n16727 )  ;
assign n16729 =  ( n16728 ) & (wr )  ;
assign n16730 =  ( n16729 ) ? ( n5096 ) : ( iram_115 ) ;
assign n16731 = wr_addr[7:7] ;
assign n16732 =  ( n16731 ) == ( bv_1_0_n53 )  ;
assign n16733 =  ( wr_addr ) == ( bv_8_115_n299 )  ;
assign n16734 =  ( n16732 ) & (n16733 )  ;
assign n16735 =  ( n16734 ) & (wr )  ;
assign n16736 =  ( n16735 ) ? ( n5123 ) : ( iram_115 ) ;
assign n16737 = wr_addr[7:7] ;
assign n16738 =  ( n16737 ) == ( bv_1_0_n53 )  ;
assign n16739 =  ( wr_addr ) == ( bv_8_115_n299 )  ;
assign n16740 =  ( n16738 ) & (n16739 )  ;
assign n16741 =  ( n16740 ) & (wr )  ;
assign n16742 =  ( n16741 ) ? ( n5165 ) : ( iram_115 ) ;
assign n16743 = wr_addr[7:7] ;
assign n16744 =  ( n16743 ) == ( bv_1_0_n53 )  ;
assign n16745 =  ( wr_addr ) == ( bv_8_115_n299 )  ;
assign n16746 =  ( n16744 ) & (n16745 )  ;
assign n16747 =  ( n16746 ) & (wr )  ;
assign n16748 =  ( n16747 ) ? ( n5204 ) : ( iram_115 ) ;
assign n16749 = wr_addr[7:7] ;
assign n16750 =  ( n16749 ) == ( bv_1_0_n53 )  ;
assign n16751 =  ( wr_addr ) == ( bv_8_115_n299 )  ;
assign n16752 =  ( n16750 ) & (n16751 )  ;
assign n16753 =  ( n16752 ) & (wr )  ;
assign n16754 =  ( n16753 ) ? ( n5262 ) : ( iram_115 ) ;
assign n16755 = wr_addr[7:7] ;
assign n16756 =  ( n16755 ) == ( bv_1_0_n53 )  ;
assign n16757 =  ( wr_addr ) == ( bv_8_115_n299 )  ;
assign n16758 =  ( n16756 ) & (n16757 )  ;
assign n16759 =  ( n16758 ) & (wr )  ;
assign n16760 =  ( n16759 ) ? ( n5298 ) : ( iram_115 ) ;
assign n16761 = wr_addr[7:7] ;
assign n16762 =  ( n16761 ) == ( bv_1_0_n53 )  ;
assign n16763 =  ( wr_addr ) == ( bv_8_115_n299 )  ;
assign n16764 =  ( n16762 ) & (n16763 )  ;
assign n16765 =  ( n16764 ) & (wr )  ;
assign n16766 =  ( n16765 ) ? ( n5325 ) : ( iram_115 ) ;
assign n16767 = wr_addr[7:7] ;
assign n16768 =  ( n16767 ) == ( bv_1_0_n53 )  ;
assign n16769 =  ( wr_addr ) == ( bv_8_116_n301 )  ;
assign n16770 =  ( n16768 ) & (n16769 )  ;
assign n16771 =  ( n16770 ) & (wr )  ;
assign n16772 =  ( n16771 ) ? ( n4782 ) : ( iram_116 ) ;
assign n16773 = wr_addr[7:7] ;
assign n16774 =  ( n16773 ) == ( bv_1_0_n53 )  ;
assign n16775 =  ( wr_addr ) == ( bv_8_116_n301 )  ;
assign n16776 =  ( n16774 ) & (n16775 )  ;
assign n16777 =  ( n16776 ) & (wr )  ;
assign n16778 =  ( n16777 ) ? ( n4841 ) : ( iram_116 ) ;
assign n16779 = wr_addr[7:7] ;
assign n16780 =  ( n16779 ) == ( bv_1_0_n53 )  ;
assign n16781 =  ( wr_addr ) == ( bv_8_116_n301 )  ;
assign n16782 =  ( n16780 ) & (n16781 )  ;
assign n16783 =  ( n16782 ) & (wr )  ;
assign n16784 =  ( n16783 ) ? ( n5449 ) : ( iram_116 ) ;
assign n16785 = wr_addr[7:7] ;
assign n16786 =  ( n16785 ) == ( bv_1_0_n53 )  ;
assign n16787 =  ( wr_addr ) == ( bv_8_116_n301 )  ;
assign n16788 =  ( n16786 ) & (n16787 )  ;
assign n16789 =  ( n16788 ) & (wr )  ;
assign n16790 =  ( n16789 ) ? ( n4906 ) : ( iram_116 ) ;
assign n16791 = wr_addr[7:7] ;
assign n16792 =  ( n16791 ) == ( bv_1_0_n53 )  ;
assign n16793 =  ( wr_addr ) == ( bv_8_116_n301 )  ;
assign n16794 =  ( n16792 ) & (n16793 )  ;
assign n16795 =  ( n16794 ) & (wr )  ;
assign n16796 =  ( n16795 ) ? ( n5485 ) : ( iram_116 ) ;
assign n16797 = wr_addr[7:7] ;
assign n16798 =  ( n16797 ) == ( bv_1_0_n53 )  ;
assign n16799 =  ( wr_addr ) == ( bv_8_116_n301 )  ;
assign n16800 =  ( n16798 ) & (n16799 )  ;
assign n16801 =  ( n16800 ) & (wr )  ;
assign n16802 =  ( n16801 ) ? ( n5512 ) : ( iram_116 ) ;
assign n16803 = wr_addr[7:7] ;
assign n16804 =  ( n16803 ) == ( bv_1_0_n53 )  ;
assign n16805 =  ( wr_addr ) == ( bv_8_116_n301 )  ;
assign n16806 =  ( n16804 ) & (n16805 )  ;
assign n16807 =  ( n16806 ) & (wr )  ;
assign n16808 =  ( n16807 ) ? ( bv_8_0_n69 ) : ( iram_116 ) ;
assign n16809 = wr_addr[7:7] ;
assign n16810 =  ( n16809 ) == ( bv_1_0_n53 )  ;
assign n16811 =  ( wr_addr ) == ( bv_8_116_n301 )  ;
assign n16812 =  ( n16810 ) & (n16811 )  ;
assign n16813 =  ( n16812 ) & (wr )  ;
assign n16814 =  ( n16813 ) ? ( n5071 ) : ( iram_116 ) ;
assign n16815 = wr_addr[7:7] ;
assign n16816 =  ( n16815 ) == ( bv_1_0_n53 )  ;
assign n16817 =  ( wr_addr ) == ( bv_8_116_n301 )  ;
assign n16818 =  ( n16816 ) & (n16817 )  ;
assign n16819 =  ( n16818 ) & (wr )  ;
assign n16820 =  ( n16819 ) ? ( n5096 ) : ( iram_116 ) ;
assign n16821 = wr_addr[7:7] ;
assign n16822 =  ( n16821 ) == ( bv_1_0_n53 )  ;
assign n16823 =  ( wr_addr ) == ( bv_8_116_n301 )  ;
assign n16824 =  ( n16822 ) & (n16823 )  ;
assign n16825 =  ( n16824 ) & (wr )  ;
assign n16826 =  ( n16825 ) ? ( n5123 ) : ( iram_116 ) ;
assign n16827 = wr_addr[7:7] ;
assign n16828 =  ( n16827 ) == ( bv_1_0_n53 )  ;
assign n16829 =  ( wr_addr ) == ( bv_8_116_n301 )  ;
assign n16830 =  ( n16828 ) & (n16829 )  ;
assign n16831 =  ( n16830 ) & (wr )  ;
assign n16832 =  ( n16831 ) ? ( n5165 ) : ( iram_116 ) ;
assign n16833 = wr_addr[7:7] ;
assign n16834 =  ( n16833 ) == ( bv_1_0_n53 )  ;
assign n16835 =  ( wr_addr ) == ( bv_8_116_n301 )  ;
assign n16836 =  ( n16834 ) & (n16835 )  ;
assign n16837 =  ( n16836 ) & (wr )  ;
assign n16838 =  ( n16837 ) ? ( n5204 ) : ( iram_116 ) ;
assign n16839 = wr_addr[7:7] ;
assign n16840 =  ( n16839 ) == ( bv_1_0_n53 )  ;
assign n16841 =  ( wr_addr ) == ( bv_8_116_n301 )  ;
assign n16842 =  ( n16840 ) & (n16841 )  ;
assign n16843 =  ( n16842 ) & (wr )  ;
assign n16844 =  ( n16843 ) ? ( n5262 ) : ( iram_116 ) ;
assign n16845 = wr_addr[7:7] ;
assign n16846 =  ( n16845 ) == ( bv_1_0_n53 )  ;
assign n16847 =  ( wr_addr ) == ( bv_8_116_n301 )  ;
assign n16848 =  ( n16846 ) & (n16847 )  ;
assign n16849 =  ( n16848 ) & (wr )  ;
assign n16850 =  ( n16849 ) ? ( n5298 ) : ( iram_116 ) ;
assign n16851 = wr_addr[7:7] ;
assign n16852 =  ( n16851 ) == ( bv_1_0_n53 )  ;
assign n16853 =  ( wr_addr ) == ( bv_8_116_n301 )  ;
assign n16854 =  ( n16852 ) & (n16853 )  ;
assign n16855 =  ( n16854 ) & (wr )  ;
assign n16856 =  ( n16855 ) ? ( n5325 ) : ( iram_116 ) ;
assign n16857 = wr_addr[7:7] ;
assign n16858 =  ( n16857 ) == ( bv_1_0_n53 )  ;
assign n16859 =  ( wr_addr ) == ( bv_8_117_n303 )  ;
assign n16860 =  ( n16858 ) & (n16859 )  ;
assign n16861 =  ( n16860 ) & (wr )  ;
assign n16862 =  ( n16861 ) ? ( n4782 ) : ( iram_117 ) ;
assign n16863 = wr_addr[7:7] ;
assign n16864 =  ( n16863 ) == ( bv_1_0_n53 )  ;
assign n16865 =  ( wr_addr ) == ( bv_8_117_n303 )  ;
assign n16866 =  ( n16864 ) & (n16865 )  ;
assign n16867 =  ( n16866 ) & (wr )  ;
assign n16868 =  ( n16867 ) ? ( n4841 ) : ( iram_117 ) ;
assign n16869 = wr_addr[7:7] ;
assign n16870 =  ( n16869 ) == ( bv_1_0_n53 )  ;
assign n16871 =  ( wr_addr ) == ( bv_8_117_n303 )  ;
assign n16872 =  ( n16870 ) & (n16871 )  ;
assign n16873 =  ( n16872 ) & (wr )  ;
assign n16874 =  ( n16873 ) ? ( n5449 ) : ( iram_117 ) ;
assign n16875 = wr_addr[7:7] ;
assign n16876 =  ( n16875 ) == ( bv_1_0_n53 )  ;
assign n16877 =  ( wr_addr ) == ( bv_8_117_n303 )  ;
assign n16878 =  ( n16876 ) & (n16877 )  ;
assign n16879 =  ( n16878 ) & (wr )  ;
assign n16880 =  ( n16879 ) ? ( n4906 ) : ( iram_117 ) ;
assign n16881 = wr_addr[7:7] ;
assign n16882 =  ( n16881 ) == ( bv_1_0_n53 )  ;
assign n16883 =  ( wr_addr ) == ( bv_8_117_n303 )  ;
assign n16884 =  ( n16882 ) & (n16883 )  ;
assign n16885 =  ( n16884 ) & (wr )  ;
assign n16886 =  ( n16885 ) ? ( n5485 ) : ( iram_117 ) ;
assign n16887 = wr_addr[7:7] ;
assign n16888 =  ( n16887 ) == ( bv_1_0_n53 )  ;
assign n16889 =  ( wr_addr ) == ( bv_8_117_n303 )  ;
assign n16890 =  ( n16888 ) & (n16889 )  ;
assign n16891 =  ( n16890 ) & (wr )  ;
assign n16892 =  ( n16891 ) ? ( n5512 ) : ( iram_117 ) ;
assign n16893 = wr_addr[7:7] ;
assign n16894 =  ( n16893 ) == ( bv_1_0_n53 )  ;
assign n16895 =  ( wr_addr ) == ( bv_8_117_n303 )  ;
assign n16896 =  ( n16894 ) & (n16895 )  ;
assign n16897 =  ( n16896 ) & (wr )  ;
assign n16898 =  ( n16897 ) ? ( bv_8_0_n69 ) : ( iram_117 ) ;
assign n16899 = wr_addr[7:7] ;
assign n16900 =  ( n16899 ) == ( bv_1_0_n53 )  ;
assign n16901 =  ( wr_addr ) == ( bv_8_117_n303 )  ;
assign n16902 =  ( n16900 ) & (n16901 )  ;
assign n16903 =  ( n16902 ) & (wr )  ;
assign n16904 =  ( n16903 ) ? ( n5071 ) : ( iram_117 ) ;
assign n16905 = wr_addr[7:7] ;
assign n16906 =  ( n16905 ) == ( bv_1_0_n53 )  ;
assign n16907 =  ( wr_addr ) == ( bv_8_117_n303 )  ;
assign n16908 =  ( n16906 ) & (n16907 )  ;
assign n16909 =  ( n16908 ) & (wr )  ;
assign n16910 =  ( n16909 ) ? ( n5096 ) : ( iram_117 ) ;
assign n16911 = wr_addr[7:7] ;
assign n16912 =  ( n16911 ) == ( bv_1_0_n53 )  ;
assign n16913 =  ( wr_addr ) == ( bv_8_117_n303 )  ;
assign n16914 =  ( n16912 ) & (n16913 )  ;
assign n16915 =  ( n16914 ) & (wr )  ;
assign n16916 =  ( n16915 ) ? ( n5123 ) : ( iram_117 ) ;
assign n16917 = wr_addr[7:7] ;
assign n16918 =  ( n16917 ) == ( bv_1_0_n53 )  ;
assign n16919 =  ( wr_addr ) == ( bv_8_117_n303 )  ;
assign n16920 =  ( n16918 ) & (n16919 )  ;
assign n16921 =  ( n16920 ) & (wr )  ;
assign n16922 =  ( n16921 ) ? ( n5165 ) : ( iram_117 ) ;
assign n16923 = wr_addr[7:7] ;
assign n16924 =  ( n16923 ) == ( bv_1_0_n53 )  ;
assign n16925 =  ( wr_addr ) == ( bv_8_117_n303 )  ;
assign n16926 =  ( n16924 ) & (n16925 )  ;
assign n16927 =  ( n16926 ) & (wr )  ;
assign n16928 =  ( n16927 ) ? ( n5204 ) : ( iram_117 ) ;
assign n16929 = wr_addr[7:7] ;
assign n16930 =  ( n16929 ) == ( bv_1_0_n53 )  ;
assign n16931 =  ( wr_addr ) == ( bv_8_117_n303 )  ;
assign n16932 =  ( n16930 ) & (n16931 )  ;
assign n16933 =  ( n16932 ) & (wr )  ;
assign n16934 =  ( n16933 ) ? ( n5262 ) : ( iram_117 ) ;
assign n16935 = wr_addr[7:7] ;
assign n16936 =  ( n16935 ) == ( bv_1_0_n53 )  ;
assign n16937 =  ( wr_addr ) == ( bv_8_117_n303 )  ;
assign n16938 =  ( n16936 ) & (n16937 )  ;
assign n16939 =  ( n16938 ) & (wr )  ;
assign n16940 =  ( n16939 ) ? ( n5298 ) : ( iram_117 ) ;
assign n16941 = wr_addr[7:7] ;
assign n16942 =  ( n16941 ) == ( bv_1_0_n53 )  ;
assign n16943 =  ( wr_addr ) == ( bv_8_117_n303 )  ;
assign n16944 =  ( n16942 ) & (n16943 )  ;
assign n16945 =  ( n16944 ) & (wr )  ;
assign n16946 =  ( n16945 ) ? ( n5325 ) : ( iram_117 ) ;
assign n16947 = wr_addr[7:7] ;
assign n16948 =  ( n16947 ) == ( bv_1_0_n53 )  ;
assign n16949 =  ( wr_addr ) == ( bv_8_118_n305 )  ;
assign n16950 =  ( n16948 ) & (n16949 )  ;
assign n16951 =  ( n16950 ) & (wr )  ;
assign n16952 =  ( n16951 ) ? ( n4782 ) : ( iram_118 ) ;
assign n16953 = wr_addr[7:7] ;
assign n16954 =  ( n16953 ) == ( bv_1_0_n53 )  ;
assign n16955 =  ( wr_addr ) == ( bv_8_118_n305 )  ;
assign n16956 =  ( n16954 ) & (n16955 )  ;
assign n16957 =  ( n16956 ) & (wr )  ;
assign n16958 =  ( n16957 ) ? ( n4841 ) : ( iram_118 ) ;
assign n16959 = wr_addr[7:7] ;
assign n16960 =  ( n16959 ) == ( bv_1_0_n53 )  ;
assign n16961 =  ( wr_addr ) == ( bv_8_118_n305 )  ;
assign n16962 =  ( n16960 ) & (n16961 )  ;
assign n16963 =  ( n16962 ) & (wr )  ;
assign n16964 =  ( n16963 ) ? ( n5449 ) : ( iram_118 ) ;
assign n16965 = wr_addr[7:7] ;
assign n16966 =  ( n16965 ) == ( bv_1_0_n53 )  ;
assign n16967 =  ( wr_addr ) == ( bv_8_118_n305 )  ;
assign n16968 =  ( n16966 ) & (n16967 )  ;
assign n16969 =  ( n16968 ) & (wr )  ;
assign n16970 =  ( n16969 ) ? ( n4906 ) : ( iram_118 ) ;
assign n16971 = wr_addr[7:7] ;
assign n16972 =  ( n16971 ) == ( bv_1_0_n53 )  ;
assign n16973 =  ( wr_addr ) == ( bv_8_118_n305 )  ;
assign n16974 =  ( n16972 ) & (n16973 )  ;
assign n16975 =  ( n16974 ) & (wr )  ;
assign n16976 =  ( n16975 ) ? ( n5485 ) : ( iram_118 ) ;
assign n16977 = wr_addr[7:7] ;
assign n16978 =  ( n16977 ) == ( bv_1_0_n53 )  ;
assign n16979 =  ( wr_addr ) == ( bv_8_118_n305 )  ;
assign n16980 =  ( n16978 ) & (n16979 )  ;
assign n16981 =  ( n16980 ) & (wr )  ;
assign n16982 =  ( n16981 ) ? ( n5512 ) : ( iram_118 ) ;
assign n16983 = wr_addr[7:7] ;
assign n16984 =  ( n16983 ) == ( bv_1_0_n53 )  ;
assign n16985 =  ( wr_addr ) == ( bv_8_118_n305 )  ;
assign n16986 =  ( n16984 ) & (n16985 )  ;
assign n16987 =  ( n16986 ) & (wr )  ;
assign n16988 =  ( n16987 ) ? ( bv_8_0_n69 ) : ( iram_118 ) ;
assign n16989 = wr_addr[7:7] ;
assign n16990 =  ( n16989 ) == ( bv_1_0_n53 )  ;
assign n16991 =  ( wr_addr ) == ( bv_8_118_n305 )  ;
assign n16992 =  ( n16990 ) & (n16991 )  ;
assign n16993 =  ( n16992 ) & (wr )  ;
assign n16994 =  ( n16993 ) ? ( n5071 ) : ( iram_118 ) ;
assign n16995 = wr_addr[7:7] ;
assign n16996 =  ( n16995 ) == ( bv_1_0_n53 )  ;
assign n16997 =  ( wr_addr ) == ( bv_8_118_n305 )  ;
assign n16998 =  ( n16996 ) & (n16997 )  ;
assign n16999 =  ( n16998 ) & (wr )  ;
assign n17000 =  ( n16999 ) ? ( n5096 ) : ( iram_118 ) ;
assign n17001 = wr_addr[7:7] ;
assign n17002 =  ( n17001 ) == ( bv_1_0_n53 )  ;
assign n17003 =  ( wr_addr ) == ( bv_8_118_n305 )  ;
assign n17004 =  ( n17002 ) & (n17003 )  ;
assign n17005 =  ( n17004 ) & (wr )  ;
assign n17006 =  ( n17005 ) ? ( n5123 ) : ( iram_118 ) ;
assign n17007 = wr_addr[7:7] ;
assign n17008 =  ( n17007 ) == ( bv_1_0_n53 )  ;
assign n17009 =  ( wr_addr ) == ( bv_8_118_n305 )  ;
assign n17010 =  ( n17008 ) & (n17009 )  ;
assign n17011 =  ( n17010 ) & (wr )  ;
assign n17012 =  ( n17011 ) ? ( n5165 ) : ( iram_118 ) ;
assign n17013 = wr_addr[7:7] ;
assign n17014 =  ( n17013 ) == ( bv_1_0_n53 )  ;
assign n17015 =  ( wr_addr ) == ( bv_8_118_n305 )  ;
assign n17016 =  ( n17014 ) & (n17015 )  ;
assign n17017 =  ( n17016 ) & (wr )  ;
assign n17018 =  ( n17017 ) ? ( n5204 ) : ( iram_118 ) ;
assign n17019 = wr_addr[7:7] ;
assign n17020 =  ( n17019 ) == ( bv_1_0_n53 )  ;
assign n17021 =  ( wr_addr ) == ( bv_8_118_n305 )  ;
assign n17022 =  ( n17020 ) & (n17021 )  ;
assign n17023 =  ( n17022 ) & (wr )  ;
assign n17024 =  ( n17023 ) ? ( n5262 ) : ( iram_118 ) ;
assign n17025 = wr_addr[7:7] ;
assign n17026 =  ( n17025 ) == ( bv_1_0_n53 )  ;
assign n17027 =  ( wr_addr ) == ( bv_8_118_n305 )  ;
assign n17028 =  ( n17026 ) & (n17027 )  ;
assign n17029 =  ( n17028 ) & (wr )  ;
assign n17030 =  ( n17029 ) ? ( n5298 ) : ( iram_118 ) ;
assign n17031 = wr_addr[7:7] ;
assign n17032 =  ( n17031 ) == ( bv_1_0_n53 )  ;
assign n17033 =  ( wr_addr ) == ( bv_8_118_n305 )  ;
assign n17034 =  ( n17032 ) & (n17033 )  ;
assign n17035 =  ( n17034 ) & (wr )  ;
assign n17036 =  ( n17035 ) ? ( n5325 ) : ( iram_118 ) ;
assign n17037 = wr_addr[7:7] ;
assign n17038 =  ( n17037 ) == ( bv_1_0_n53 )  ;
assign n17039 =  ( wr_addr ) == ( bv_8_119_n307 )  ;
assign n17040 =  ( n17038 ) & (n17039 )  ;
assign n17041 =  ( n17040 ) & (wr )  ;
assign n17042 =  ( n17041 ) ? ( n4782 ) : ( iram_119 ) ;
assign n17043 = wr_addr[7:7] ;
assign n17044 =  ( n17043 ) == ( bv_1_0_n53 )  ;
assign n17045 =  ( wr_addr ) == ( bv_8_119_n307 )  ;
assign n17046 =  ( n17044 ) & (n17045 )  ;
assign n17047 =  ( n17046 ) & (wr )  ;
assign n17048 =  ( n17047 ) ? ( n4841 ) : ( iram_119 ) ;
assign n17049 = wr_addr[7:7] ;
assign n17050 =  ( n17049 ) == ( bv_1_0_n53 )  ;
assign n17051 =  ( wr_addr ) == ( bv_8_119_n307 )  ;
assign n17052 =  ( n17050 ) & (n17051 )  ;
assign n17053 =  ( n17052 ) & (wr )  ;
assign n17054 =  ( n17053 ) ? ( n5449 ) : ( iram_119 ) ;
assign n17055 = wr_addr[7:7] ;
assign n17056 =  ( n17055 ) == ( bv_1_0_n53 )  ;
assign n17057 =  ( wr_addr ) == ( bv_8_119_n307 )  ;
assign n17058 =  ( n17056 ) & (n17057 )  ;
assign n17059 =  ( n17058 ) & (wr )  ;
assign n17060 =  ( n17059 ) ? ( n4906 ) : ( iram_119 ) ;
assign n17061 = wr_addr[7:7] ;
assign n17062 =  ( n17061 ) == ( bv_1_0_n53 )  ;
assign n17063 =  ( wr_addr ) == ( bv_8_119_n307 )  ;
assign n17064 =  ( n17062 ) & (n17063 )  ;
assign n17065 =  ( n17064 ) & (wr )  ;
assign n17066 =  ( n17065 ) ? ( n5485 ) : ( iram_119 ) ;
assign n17067 = wr_addr[7:7] ;
assign n17068 =  ( n17067 ) == ( bv_1_0_n53 )  ;
assign n17069 =  ( wr_addr ) == ( bv_8_119_n307 )  ;
assign n17070 =  ( n17068 ) & (n17069 )  ;
assign n17071 =  ( n17070 ) & (wr )  ;
assign n17072 =  ( n17071 ) ? ( n5512 ) : ( iram_119 ) ;
assign n17073 = wr_addr[7:7] ;
assign n17074 =  ( n17073 ) == ( bv_1_0_n53 )  ;
assign n17075 =  ( wr_addr ) == ( bv_8_119_n307 )  ;
assign n17076 =  ( n17074 ) & (n17075 )  ;
assign n17077 =  ( n17076 ) & (wr )  ;
assign n17078 =  ( n17077 ) ? ( bv_8_0_n69 ) : ( iram_119 ) ;
assign n17079 = wr_addr[7:7] ;
assign n17080 =  ( n17079 ) == ( bv_1_0_n53 )  ;
assign n17081 =  ( wr_addr ) == ( bv_8_119_n307 )  ;
assign n17082 =  ( n17080 ) & (n17081 )  ;
assign n17083 =  ( n17082 ) & (wr )  ;
assign n17084 =  ( n17083 ) ? ( n5071 ) : ( iram_119 ) ;
assign n17085 = wr_addr[7:7] ;
assign n17086 =  ( n17085 ) == ( bv_1_0_n53 )  ;
assign n17087 =  ( wr_addr ) == ( bv_8_119_n307 )  ;
assign n17088 =  ( n17086 ) & (n17087 )  ;
assign n17089 =  ( n17088 ) & (wr )  ;
assign n17090 =  ( n17089 ) ? ( n5096 ) : ( iram_119 ) ;
assign n17091 = wr_addr[7:7] ;
assign n17092 =  ( n17091 ) == ( bv_1_0_n53 )  ;
assign n17093 =  ( wr_addr ) == ( bv_8_119_n307 )  ;
assign n17094 =  ( n17092 ) & (n17093 )  ;
assign n17095 =  ( n17094 ) & (wr )  ;
assign n17096 =  ( n17095 ) ? ( n5123 ) : ( iram_119 ) ;
assign n17097 = wr_addr[7:7] ;
assign n17098 =  ( n17097 ) == ( bv_1_0_n53 )  ;
assign n17099 =  ( wr_addr ) == ( bv_8_119_n307 )  ;
assign n17100 =  ( n17098 ) & (n17099 )  ;
assign n17101 =  ( n17100 ) & (wr )  ;
assign n17102 =  ( n17101 ) ? ( n5165 ) : ( iram_119 ) ;
assign n17103 = wr_addr[7:7] ;
assign n17104 =  ( n17103 ) == ( bv_1_0_n53 )  ;
assign n17105 =  ( wr_addr ) == ( bv_8_119_n307 )  ;
assign n17106 =  ( n17104 ) & (n17105 )  ;
assign n17107 =  ( n17106 ) & (wr )  ;
assign n17108 =  ( n17107 ) ? ( n5204 ) : ( iram_119 ) ;
assign n17109 = wr_addr[7:7] ;
assign n17110 =  ( n17109 ) == ( bv_1_0_n53 )  ;
assign n17111 =  ( wr_addr ) == ( bv_8_119_n307 )  ;
assign n17112 =  ( n17110 ) & (n17111 )  ;
assign n17113 =  ( n17112 ) & (wr )  ;
assign n17114 =  ( n17113 ) ? ( n5262 ) : ( iram_119 ) ;
assign n17115 = wr_addr[7:7] ;
assign n17116 =  ( n17115 ) == ( bv_1_0_n53 )  ;
assign n17117 =  ( wr_addr ) == ( bv_8_119_n307 )  ;
assign n17118 =  ( n17116 ) & (n17117 )  ;
assign n17119 =  ( n17118 ) & (wr )  ;
assign n17120 =  ( n17119 ) ? ( n5298 ) : ( iram_119 ) ;
assign n17121 = wr_addr[7:7] ;
assign n17122 =  ( n17121 ) == ( bv_1_0_n53 )  ;
assign n17123 =  ( wr_addr ) == ( bv_8_119_n307 )  ;
assign n17124 =  ( n17122 ) & (n17123 )  ;
assign n17125 =  ( n17124 ) & (wr )  ;
assign n17126 =  ( n17125 ) ? ( n5325 ) : ( iram_119 ) ;
assign n17127 = wr_addr[7:7] ;
assign n17128 =  ( n17127 ) == ( bv_1_0_n53 )  ;
assign n17129 =  ( wr_addr ) == ( bv_8_120_n309 )  ;
assign n17130 =  ( n17128 ) & (n17129 )  ;
assign n17131 =  ( n17130 ) & (wr )  ;
assign n17132 =  ( n17131 ) ? ( n4782 ) : ( iram_120 ) ;
assign n17133 = wr_addr[7:7] ;
assign n17134 =  ( n17133 ) == ( bv_1_0_n53 )  ;
assign n17135 =  ( wr_addr ) == ( bv_8_120_n309 )  ;
assign n17136 =  ( n17134 ) & (n17135 )  ;
assign n17137 =  ( n17136 ) & (wr )  ;
assign n17138 =  ( n17137 ) ? ( n4841 ) : ( iram_120 ) ;
assign n17139 = wr_addr[7:7] ;
assign n17140 =  ( n17139 ) == ( bv_1_0_n53 )  ;
assign n17141 =  ( wr_addr ) == ( bv_8_120_n309 )  ;
assign n17142 =  ( n17140 ) & (n17141 )  ;
assign n17143 =  ( n17142 ) & (wr )  ;
assign n17144 =  ( n17143 ) ? ( n5449 ) : ( iram_120 ) ;
assign n17145 = wr_addr[7:7] ;
assign n17146 =  ( n17145 ) == ( bv_1_0_n53 )  ;
assign n17147 =  ( wr_addr ) == ( bv_8_120_n309 )  ;
assign n17148 =  ( n17146 ) & (n17147 )  ;
assign n17149 =  ( n17148 ) & (wr )  ;
assign n17150 =  ( n17149 ) ? ( n4906 ) : ( iram_120 ) ;
assign n17151 = wr_addr[7:7] ;
assign n17152 =  ( n17151 ) == ( bv_1_0_n53 )  ;
assign n17153 =  ( wr_addr ) == ( bv_8_120_n309 )  ;
assign n17154 =  ( n17152 ) & (n17153 )  ;
assign n17155 =  ( n17154 ) & (wr )  ;
assign n17156 =  ( n17155 ) ? ( n5485 ) : ( iram_120 ) ;
assign n17157 = wr_addr[7:7] ;
assign n17158 =  ( n17157 ) == ( bv_1_0_n53 )  ;
assign n17159 =  ( wr_addr ) == ( bv_8_120_n309 )  ;
assign n17160 =  ( n17158 ) & (n17159 )  ;
assign n17161 =  ( n17160 ) & (wr )  ;
assign n17162 =  ( n17161 ) ? ( n5512 ) : ( iram_120 ) ;
assign n17163 = wr_addr[7:7] ;
assign n17164 =  ( n17163 ) == ( bv_1_0_n53 )  ;
assign n17165 =  ( wr_addr ) == ( bv_8_120_n309 )  ;
assign n17166 =  ( n17164 ) & (n17165 )  ;
assign n17167 =  ( n17166 ) & (wr )  ;
assign n17168 =  ( n17167 ) ? ( bv_8_0_n69 ) : ( iram_120 ) ;
assign n17169 = wr_addr[7:7] ;
assign n17170 =  ( n17169 ) == ( bv_1_0_n53 )  ;
assign n17171 =  ( wr_addr ) == ( bv_8_120_n309 )  ;
assign n17172 =  ( n17170 ) & (n17171 )  ;
assign n17173 =  ( n17172 ) & (wr )  ;
assign n17174 =  ( n17173 ) ? ( n5071 ) : ( iram_120 ) ;
assign n17175 = wr_addr[7:7] ;
assign n17176 =  ( n17175 ) == ( bv_1_0_n53 )  ;
assign n17177 =  ( wr_addr ) == ( bv_8_120_n309 )  ;
assign n17178 =  ( n17176 ) & (n17177 )  ;
assign n17179 =  ( n17178 ) & (wr )  ;
assign n17180 =  ( n17179 ) ? ( n5096 ) : ( iram_120 ) ;
assign n17181 = wr_addr[7:7] ;
assign n17182 =  ( n17181 ) == ( bv_1_0_n53 )  ;
assign n17183 =  ( wr_addr ) == ( bv_8_120_n309 )  ;
assign n17184 =  ( n17182 ) & (n17183 )  ;
assign n17185 =  ( n17184 ) & (wr )  ;
assign n17186 =  ( n17185 ) ? ( n5123 ) : ( iram_120 ) ;
assign n17187 = wr_addr[7:7] ;
assign n17188 =  ( n17187 ) == ( bv_1_0_n53 )  ;
assign n17189 =  ( wr_addr ) == ( bv_8_120_n309 )  ;
assign n17190 =  ( n17188 ) & (n17189 )  ;
assign n17191 =  ( n17190 ) & (wr )  ;
assign n17192 =  ( n17191 ) ? ( n5165 ) : ( iram_120 ) ;
assign n17193 = wr_addr[7:7] ;
assign n17194 =  ( n17193 ) == ( bv_1_0_n53 )  ;
assign n17195 =  ( wr_addr ) == ( bv_8_120_n309 )  ;
assign n17196 =  ( n17194 ) & (n17195 )  ;
assign n17197 =  ( n17196 ) & (wr )  ;
assign n17198 =  ( n17197 ) ? ( n5204 ) : ( iram_120 ) ;
assign n17199 = wr_addr[7:7] ;
assign n17200 =  ( n17199 ) == ( bv_1_0_n53 )  ;
assign n17201 =  ( wr_addr ) == ( bv_8_120_n309 )  ;
assign n17202 =  ( n17200 ) & (n17201 )  ;
assign n17203 =  ( n17202 ) & (wr )  ;
assign n17204 =  ( n17203 ) ? ( n5262 ) : ( iram_120 ) ;
assign n17205 = wr_addr[7:7] ;
assign n17206 =  ( n17205 ) == ( bv_1_0_n53 )  ;
assign n17207 =  ( wr_addr ) == ( bv_8_120_n309 )  ;
assign n17208 =  ( n17206 ) & (n17207 )  ;
assign n17209 =  ( n17208 ) & (wr )  ;
assign n17210 =  ( n17209 ) ? ( n5298 ) : ( iram_120 ) ;
assign n17211 = wr_addr[7:7] ;
assign n17212 =  ( n17211 ) == ( bv_1_0_n53 )  ;
assign n17213 =  ( wr_addr ) == ( bv_8_120_n309 )  ;
assign n17214 =  ( n17212 ) & (n17213 )  ;
assign n17215 =  ( n17214 ) & (wr )  ;
assign n17216 =  ( n17215 ) ? ( n5325 ) : ( iram_120 ) ;
assign n17217 = wr_addr[7:7] ;
assign n17218 =  ( n17217 ) == ( bv_1_0_n53 )  ;
assign n17219 =  ( wr_addr ) == ( bv_8_121_n311 )  ;
assign n17220 =  ( n17218 ) & (n17219 )  ;
assign n17221 =  ( n17220 ) & (wr )  ;
assign n17222 =  ( n17221 ) ? ( n4782 ) : ( iram_121 ) ;
assign n17223 = wr_addr[7:7] ;
assign n17224 =  ( n17223 ) == ( bv_1_0_n53 )  ;
assign n17225 =  ( wr_addr ) == ( bv_8_121_n311 )  ;
assign n17226 =  ( n17224 ) & (n17225 )  ;
assign n17227 =  ( n17226 ) & (wr )  ;
assign n17228 =  ( n17227 ) ? ( n4841 ) : ( iram_121 ) ;
assign n17229 = wr_addr[7:7] ;
assign n17230 =  ( n17229 ) == ( bv_1_0_n53 )  ;
assign n17231 =  ( wr_addr ) == ( bv_8_121_n311 )  ;
assign n17232 =  ( n17230 ) & (n17231 )  ;
assign n17233 =  ( n17232 ) & (wr )  ;
assign n17234 =  ( n17233 ) ? ( n5449 ) : ( iram_121 ) ;
assign n17235 = wr_addr[7:7] ;
assign n17236 =  ( n17235 ) == ( bv_1_0_n53 )  ;
assign n17237 =  ( wr_addr ) == ( bv_8_121_n311 )  ;
assign n17238 =  ( n17236 ) & (n17237 )  ;
assign n17239 =  ( n17238 ) & (wr )  ;
assign n17240 =  ( n17239 ) ? ( n4906 ) : ( iram_121 ) ;
assign n17241 = wr_addr[7:7] ;
assign n17242 =  ( n17241 ) == ( bv_1_0_n53 )  ;
assign n17243 =  ( wr_addr ) == ( bv_8_121_n311 )  ;
assign n17244 =  ( n17242 ) & (n17243 )  ;
assign n17245 =  ( n17244 ) & (wr )  ;
assign n17246 =  ( n17245 ) ? ( n5485 ) : ( iram_121 ) ;
assign n17247 = wr_addr[7:7] ;
assign n17248 =  ( n17247 ) == ( bv_1_0_n53 )  ;
assign n17249 =  ( wr_addr ) == ( bv_8_121_n311 )  ;
assign n17250 =  ( n17248 ) & (n17249 )  ;
assign n17251 =  ( n17250 ) & (wr )  ;
assign n17252 =  ( n17251 ) ? ( n5512 ) : ( iram_121 ) ;
assign n17253 = wr_addr[7:7] ;
assign n17254 =  ( n17253 ) == ( bv_1_0_n53 )  ;
assign n17255 =  ( wr_addr ) == ( bv_8_121_n311 )  ;
assign n17256 =  ( n17254 ) & (n17255 )  ;
assign n17257 =  ( n17256 ) & (wr )  ;
assign n17258 =  ( n17257 ) ? ( bv_8_0_n69 ) : ( iram_121 ) ;
assign n17259 = wr_addr[7:7] ;
assign n17260 =  ( n17259 ) == ( bv_1_0_n53 )  ;
assign n17261 =  ( wr_addr ) == ( bv_8_121_n311 )  ;
assign n17262 =  ( n17260 ) & (n17261 )  ;
assign n17263 =  ( n17262 ) & (wr )  ;
assign n17264 =  ( n17263 ) ? ( n5071 ) : ( iram_121 ) ;
assign n17265 = wr_addr[7:7] ;
assign n17266 =  ( n17265 ) == ( bv_1_0_n53 )  ;
assign n17267 =  ( wr_addr ) == ( bv_8_121_n311 )  ;
assign n17268 =  ( n17266 ) & (n17267 )  ;
assign n17269 =  ( n17268 ) & (wr )  ;
assign n17270 =  ( n17269 ) ? ( n5096 ) : ( iram_121 ) ;
assign n17271 = wr_addr[7:7] ;
assign n17272 =  ( n17271 ) == ( bv_1_0_n53 )  ;
assign n17273 =  ( wr_addr ) == ( bv_8_121_n311 )  ;
assign n17274 =  ( n17272 ) & (n17273 )  ;
assign n17275 =  ( n17274 ) & (wr )  ;
assign n17276 =  ( n17275 ) ? ( n5123 ) : ( iram_121 ) ;
assign n17277 = wr_addr[7:7] ;
assign n17278 =  ( n17277 ) == ( bv_1_0_n53 )  ;
assign n17279 =  ( wr_addr ) == ( bv_8_121_n311 )  ;
assign n17280 =  ( n17278 ) & (n17279 )  ;
assign n17281 =  ( n17280 ) & (wr )  ;
assign n17282 =  ( n17281 ) ? ( n5165 ) : ( iram_121 ) ;
assign n17283 = wr_addr[7:7] ;
assign n17284 =  ( n17283 ) == ( bv_1_0_n53 )  ;
assign n17285 =  ( wr_addr ) == ( bv_8_121_n311 )  ;
assign n17286 =  ( n17284 ) & (n17285 )  ;
assign n17287 =  ( n17286 ) & (wr )  ;
assign n17288 =  ( n17287 ) ? ( n5204 ) : ( iram_121 ) ;
assign n17289 = wr_addr[7:7] ;
assign n17290 =  ( n17289 ) == ( bv_1_0_n53 )  ;
assign n17291 =  ( wr_addr ) == ( bv_8_121_n311 )  ;
assign n17292 =  ( n17290 ) & (n17291 )  ;
assign n17293 =  ( n17292 ) & (wr )  ;
assign n17294 =  ( n17293 ) ? ( n5262 ) : ( iram_121 ) ;
assign n17295 = wr_addr[7:7] ;
assign n17296 =  ( n17295 ) == ( bv_1_0_n53 )  ;
assign n17297 =  ( wr_addr ) == ( bv_8_121_n311 )  ;
assign n17298 =  ( n17296 ) & (n17297 )  ;
assign n17299 =  ( n17298 ) & (wr )  ;
assign n17300 =  ( n17299 ) ? ( n5298 ) : ( iram_121 ) ;
assign n17301 = wr_addr[7:7] ;
assign n17302 =  ( n17301 ) == ( bv_1_0_n53 )  ;
assign n17303 =  ( wr_addr ) == ( bv_8_121_n311 )  ;
assign n17304 =  ( n17302 ) & (n17303 )  ;
assign n17305 =  ( n17304 ) & (wr )  ;
assign n17306 =  ( n17305 ) ? ( n5325 ) : ( iram_121 ) ;
assign n17307 = wr_addr[7:7] ;
assign n17308 =  ( n17307 ) == ( bv_1_0_n53 )  ;
assign n17309 =  ( wr_addr ) == ( bv_8_122_n313 )  ;
assign n17310 =  ( n17308 ) & (n17309 )  ;
assign n17311 =  ( n17310 ) & (wr )  ;
assign n17312 =  ( n17311 ) ? ( n4782 ) : ( iram_122 ) ;
assign n17313 = wr_addr[7:7] ;
assign n17314 =  ( n17313 ) == ( bv_1_0_n53 )  ;
assign n17315 =  ( wr_addr ) == ( bv_8_122_n313 )  ;
assign n17316 =  ( n17314 ) & (n17315 )  ;
assign n17317 =  ( n17316 ) & (wr )  ;
assign n17318 =  ( n17317 ) ? ( n4841 ) : ( iram_122 ) ;
assign n17319 = wr_addr[7:7] ;
assign n17320 =  ( n17319 ) == ( bv_1_0_n53 )  ;
assign n17321 =  ( wr_addr ) == ( bv_8_122_n313 )  ;
assign n17322 =  ( n17320 ) & (n17321 )  ;
assign n17323 =  ( n17322 ) & (wr )  ;
assign n17324 =  ( n17323 ) ? ( n5449 ) : ( iram_122 ) ;
assign n17325 = wr_addr[7:7] ;
assign n17326 =  ( n17325 ) == ( bv_1_0_n53 )  ;
assign n17327 =  ( wr_addr ) == ( bv_8_122_n313 )  ;
assign n17328 =  ( n17326 ) & (n17327 )  ;
assign n17329 =  ( n17328 ) & (wr )  ;
assign n17330 =  ( n17329 ) ? ( n4906 ) : ( iram_122 ) ;
assign n17331 = wr_addr[7:7] ;
assign n17332 =  ( n17331 ) == ( bv_1_0_n53 )  ;
assign n17333 =  ( wr_addr ) == ( bv_8_122_n313 )  ;
assign n17334 =  ( n17332 ) & (n17333 )  ;
assign n17335 =  ( n17334 ) & (wr )  ;
assign n17336 =  ( n17335 ) ? ( n5485 ) : ( iram_122 ) ;
assign n17337 = wr_addr[7:7] ;
assign n17338 =  ( n17337 ) == ( bv_1_0_n53 )  ;
assign n17339 =  ( wr_addr ) == ( bv_8_122_n313 )  ;
assign n17340 =  ( n17338 ) & (n17339 )  ;
assign n17341 =  ( n17340 ) & (wr )  ;
assign n17342 =  ( n17341 ) ? ( n5512 ) : ( iram_122 ) ;
assign n17343 = wr_addr[7:7] ;
assign n17344 =  ( n17343 ) == ( bv_1_0_n53 )  ;
assign n17345 =  ( wr_addr ) == ( bv_8_122_n313 )  ;
assign n17346 =  ( n17344 ) & (n17345 )  ;
assign n17347 =  ( n17346 ) & (wr )  ;
assign n17348 =  ( n17347 ) ? ( bv_8_0_n69 ) : ( iram_122 ) ;
assign n17349 = wr_addr[7:7] ;
assign n17350 =  ( n17349 ) == ( bv_1_0_n53 )  ;
assign n17351 =  ( wr_addr ) == ( bv_8_122_n313 )  ;
assign n17352 =  ( n17350 ) & (n17351 )  ;
assign n17353 =  ( n17352 ) & (wr )  ;
assign n17354 =  ( n17353 ) ? ( n5071 ) : ( iram_122 ) ;
assign n17355 = wr_addr[7:7] ;
assign n17356 =  ( n17355 ) == ( bv_1_0_n53 )  ;
assign n17357 =  ( wr_addr ) == ( bv_8_122_n313 )  ;
assign n17358 =  ( n17356 ) & (n17357 )  ;
assign n17359 =  ( n17358 ) & (wr )  ;
assign n17360 =  ( n17359 ) ? ( n5096 ) : ( iram_122 ) ;
assign n17361 = wr_addr[7:7] ;
assign n17362 =  ( n17361 ) == ( bv_1_0_n53 )  ;
assign n17363 =  ( wr_addr ) == ( bv_8_122_n313 )  ;
assign n17364 =  ( n17362 ) & (n17363 )  ;
assign n17365 =  ( n17364 ) & (wr )  ;
assign n17366 =  ( n17365 ) ? ( n5123 ) : ( iram_122 ) ;
assign n17367 = wr_addr[7:7] ;
assign n17368 =  ( n17367 ) == ( bv_1_0_n53 )  ;
assign n17369 =  ( wr_addr ) == ( bv_8_122_n313 )  ;
assign n17370 =  ( n17368 ) & (n17369 )  ;
assign n17371 =  ( n17370 ) & (wr )  ;
assign n17372 =  ( n17371 ) ? ( n5165 ) : ( iram_122 ) ;
assign n17373 = wr_addr[7:7] ;
assign n17374 =  ( n17373 ) == ( bv_1_0_n53 )  ;
assign n17375 =  ( wr_addr ) == ( bv_8_122_n313 )  ;
assign n17376 =  ( n17374 ) & (n17375 )  ;
assign n17377 =  ( n17376 ) & (wr )  ;
assign n17378 =  ( n17377 ) ? ( n5204 ) : ( iram_122 ) ;
assign n17379 = wr_addr[7:7] ;
assign n17380 =  ( n17379 ) == ( bv_1_0_n53 )  ;
assign n17381 =  ( wr_addr ) == ( bv_8_122_n313 )  ;
assign n17382 =  ( n17380 ) & (n17381 )  ;
assign n17383 =  ( n17382 ) & (wr )  ;
assign n17384 =  ( n17383 ) ? ( n5262 ) : ( iram_122 ) ;
assign n17385 = wr_addr[7:7] ;
assign n17386 =  ( n17385 ) == ( bv_1_0_n53 )  ;
assign n17387 =  ( wr_addr ) == ( bv_8_122_n313 )  ;
assign n17388 =  ( n17386 ) & (n17387 )  ;
assign n17389 =  ( n17388 ) & (wr )  ;
assign n17390 =  ( n17389 ) ? ( n5298 ) : ( iram_122 ) ;
assign n17391 = wr_addr[7:7] ;
assign n17392 =  ( n17391 ) == ( bv_1_0_n53 )  ;
assign n17393 =  ( wr_addr ) == ( bv_8_122_n313 )  ;
assign n17394 =  ( n17392 ) & (n17393 )  ;
assign n17395 =  ( n17394 ) & (wr )  ;
assign n17396 =  ( n17395 ) ? ( n5325 ) : ( iram_122 ) ;
assign n17397 = wr_addr[7:7] ;
assign n17398 =  ( n17397 ) == ( bv_1_0_n53 )  ;
assign n17399 =  ( wr_addr ) == ( bv_8_123_n315 )  ;
assign n17400 =  ( n17398 ) & (n17399 )  ;
assign n17401 =  ( n17400 ) & (wr )  ;
assign n17402 =  ( n17401 ) ? ( n4782 ) : ( iram_123 ) ;
assign n17403 = wr_addr[7:7] ;
assign n17404 =  ( n17403 ) == ( bv_1_0_n53 )  ;
assign n17405 =  ( wr_addr ) == ( bv_8_123_n315 )  ;
assign n17406 =  ( n17404 ) & (n17405 )  ;
assign n17407 =  ( n17406 ) & (wr )  ;
assign n17408 =  ( n17407 ) ? ( n4841 ) : ( iram_123 ) ;
assign n17409 = wr_addr[7:7] ;
assign n17410 =  ( n17409 ) == ( bv_1_0_n53 )  ;
assign n17411 =  ( wr_addr ) == ( bv_8_123_n315 )  ;
assign n17412 =  ( n17410 ) & (n17411 )  ;
assign n17413 =  ( n17412 ) & (wr )  ;
assign n17414 =  ( n17413 ) ? ( n5449 ) : ( iram_123 ) ;
assign n17415 = wr_addr[7:7] ;
assign n17416 =  ( n17415 ) == ( bv_1_0_n53 )  ;
assign n17417 =  ( wr_addr ) == ( bv_8_123_n315 )  ;
assign n17418 =  ( n17416 ) & (n17417 )  ;
assign n17419 =  ( n17418 ) & (wr )  ;
assign n17420 =  ( n17419 ) ? ( n4906 ) : ( iram_123 ) ;
assign n17421 = wr_addr[7:7] ;
assign n17422 =  ( n17421 ) == ( bv_1_0_n53 )  ;
assign n17423 =  ( wr_addr ) == ( bv_8_123_n315 )  ;
assign n17424 =  ( n17422 ) & (n17423 )  ;
assign n17425 =  ( n17424 ) & (wr )  ;
assign n17426 =  ( n17425 ) ? ( n5485 ) : ( iram_123 ) ;
assign n17427 = wr_addr[7:7] ;
assign n17428 =  ( n17427 ) == ( bv_1_0_n53 )  ;
assign n17429 =  ( wr_addr ) == ( bv_8_123_n315 )  ;
assign n17430 =  ( n17428 ) & (n17429 )  ;
assign n17431 =  ( n17430 ) & (wr )  ;
assign n17432 =  ( n17431 ) ? ( n5512 ) : ( iram_123 ) ;
assign n17433 = wr_addr[7:7] ;
assign n17434 =  ( n17433 ) == ( bv_1_0_n53 )  ;
assign n17435 =  ( wr_addr ) == ( bv_8_123_n315 )  ;
assign n17436 =  ( n17434 ) & (n17435 )  ;
assign n17437 =  ( n17436 ) & (wr )  ;
assign n17438 =  ( n17437 ) ? ( bv_8_0_n69 ) : ( iram_123 ) ;
assign n17439 = wr_addr[7:7] ;
assign n17440 =  ( n17439 ) == ( bv_1_0_n53 )  ;
assign n17441 =  ( wr_addr ) == ( bv_8_123_n315 )  ;
assign n17442 =  ( n17440 ) & (n17441 )  ;
assign n17443 =  ( n17442 ) & (wr )  ;
assign n17444 =  ( n17443 ) ? ( n5071 ) : ( iram_123 ) ;
assign n17445 = wr_addr[7:7] ;
assign n17446 =  ( n17445 ) == ( bv_1_0_n53 )  ;
assign n17447 =  ( wr_addr ) == ( bv_8_123_n315 )  ;
assign n17448 =  ( n17446 ) & (n17447 )  ;
assign n17449 =  ( n17448 ) & (wr )  ;
assign n17450 =  ( n17449 ) ? ( n5096 ) : ( iram_123 ) ;
assign n17451 = wr_addr[7:7] ;
assign n17452 =  ( n17451 ) == ( bv_1_0_n53 )  ;
assign n17453 =  ( wr_addr ) == ( bv_8_123_n315 )  ;
assign n17454 =  ( n17452 ) & (n17453 )  ;
assign n17455 =  ( n17454 ) & (wr )  ;
assign n17456 =  ( n17455 ) ? ( n5123 ) : ( iram_123 ) ;
assign n17457 = wr_addr[7:7] ;
assign n17458 =  ( n17457 ) == ( bv_1_0_n53 )  ;
assign n17459 =  ( wr_addr ) == ( bv_8_123_n315 )  ;
assign n17460 =  ( n17458 ) & (n17459 )  ;
assign n17461 =  ( n17460 ) & (wr )  ;
assign n17462 =  ( n17461 ) ? ( n5165 ) : ( iram_123 ) ;
assign n17463 = wr_addr[7:7] ;
assign n17464 =  ( n17463 ) == ( bv_1_0_n53 )  ;
assign n17465 =  ( wr_addr ) == ( bv_8_123_n315 )  ;
assign n17466 =  ( n17464 ) & (n17465 )  ;
assign n17467 =  ( n17466 ) & (wr )  ;
assign n17468 =  ( n17467 ) ? ( n5204 ) : ( iram_123 ) ;
assign n17469 = wr_addr[7:7] ;
assign n17470 =  ( n17469 ) == ( bv_1_0_n53 )  ;
assign n17471 =  ( wr_addr ) == ( bv_8_123_n315 )  ;
assign n17472 =  ( n17470 ) & (n17471 )  ;
assign n17473 =  ( n17472 ) & (wr )  ;
assign n17474 =  ( n17473 ) ? ( n5262 ) : ( iram_123 ) ;
assign n17475 = wr_addr[7:7] ;
assign n17476 =  ( n17475 ) == ( bv_1_0_n53 )  ;
assign n17477 =  ( wr_addr ) == ( bv_8_123_n315 )  ;
assign n17478 =  ( n17476 ) & (n17477 )  ;
assign n17479 =  ( n17478 ) & (wr )  ;
assign n17480 =  ( n17479 ) ? ( n5298 ) : ( iram_123 ) ;
assign n17481 = wr_addr[7:7] ;
assign n17482 =  ( n17481 ) == ( bv_1_0_n53 )  ;
assign n17483 =  ( wr_addr ) == ( bv_8_123_n315 )  ;
assign n17484 =  ( n17482 ) & (n17483 )  ;
assign n17485 =  ( n17484 ) & (wr )  ;
assign n17486 =  ( n17485 ) ? ( n5325 ) : ( iram_123 ) ;
assign n17487 = wr_addr[7:7] ;
assign n17488 =  ( n17487 ) == ( bv_1_0_n53 )  ;
assign n17489 =  ( wr_addr ) == ( bv_8_124_n317 )  ;
assign n17490 =  ( n17488 ) & (n17489 )  ;
assign n17491 =  ( n17490 ) & (wr )  ;
assign n17492 =  ( n17491 ) ? ( n4782 ) : ( iram_124 ) ;
assign n17493 = wr_addr[7:7] ;
assign n17494 =  ( n17493 ) == ( bv_1_0_n53 )  ;
assign n17495 =  ( wr_addr ) == ( bv_8_124_n317 )  ;
assign n17496 =  ( n17494 ) & (n17495 )  ;
assign n17497 =  ( n17496 ) & (wr )  ;
assign n17498 =  ( n17497 ) ? ( n4841 ) : ( iram_124 ) ;
assign n17499 = wr_addr[7:7] ;
assign n17500 =  ( n17499 ) == ( bv_1_0_n53 )  ;
assign n17501 =  ( wr_addr ) == ( bv_8_124_n317 )  ;
assign n17502 =  ( n17500 ) & (n17501 )  ;
assign n17503 =  ( n17502 ) & (wr )  ;
assign n17504 =  ( n17503 ) ? ( n5449 ) : ( iram_124 ) ;
assign n17505 = wr_addr[7:7] ;
assign n17506 =  ( n17505 ) == ( bv_1_0_n53 )  ;
assign n17507 =  ( wr_addr ) == ( bv_8_124_n317 )  ;
assign n17508 =  ( n17506 ) & (n17507 )  ;
assign n17509 =  ( n17508 ) & (wr )  ;
assign n17510 =  ( n17509 ) ? ( n4906 ) : ( iram_124 ) ;
assign n17511 = wr_addr[7:7] ;
assign n17512 =  ( n17511 ) == ( bv_1_0_n53 )  ;
assign n17513 =  ( wr_addr ) == ( bv_8_124_n317 )  ;
assign n17514 =  ( n17512 ) & (n17513 )  ;
assign n17515 =  ( n17514 ) & (wr )  ;
assign n17516 =  ( n17515 ) ? ( n5485 ) : ( iram_124 ) ;
assign n17517 = wr_addr[7:7] ;
assign n17518 =  ( n17517 ) == ( bv_1_0_n53 )  ;
assign n17519 =  ( wr_addr ) == ( bv_8_124_n317 )  ;
assign n17520 =  ( n17518 ) & (n17519 )  ;
assign n17521 =  ( n17520 ) & (wr )  ;
assign n17522 =  ( n17521 ) ? ( n5512 ) : ( iram_124 ) ;
assign n17523 = wr_addr[7:7] ;
assign n17524 =  ( n17523 ) == ( bv_1_0_n53 )  ;
assign n17525 =  ( wr_addr ) == ( bv_8_124_n317 )  ;
assign n17526 =  ( n17524 ) & (n17525 )  ;
assign n17527 =  ( n17526 ) & (wr )  ;
assign n17528 =  ( n17527 ) ? ( bv_8_0_n69 ) : ( iram_124 ) ;
assign n17529 = wr_addr[7:7] ;
assign n17530 =  ( n17529 ) == ( bv_1_0_n53 )  ;
assign n17531 =  ( wr_addr ) == ( bv_8_124_n317 )  ;
assign n17532 =  ( n17530 ) & (n17531 )  ;
assign n17533 =  ( n17532 ) & (wr )  ;
assign n17534 =  ( n17533 ) ? ( n5071 ) : ( iram_124 ) ;
assign n17535 = wr_addr[7:7] ;
assign n17536 =  ( n17535 ) == ( bv_1_0_n53 )  ;
assign n17537 =  ( wr_addr ) == ( bv_8_124_n317 )  ;
assign n17538 =  ( n17536 ) & (n17537 )  ;
assign n17539 =  ( n17538 ) & (wr )  ;
assign n17540 =  ( n17539 ) ? ( n5096 ) : ( iram_124 ) ;
assign n17541 = wr_addr[7:7] ;
assign n17542 =  ( n17541 ) == ( bv_1_0_n53 )  ;
assign n17543 =  ( wr_addr ) == ( bv_8_124_n317 )  ;
assign n17544 =  ( n17542 ) & (n17543 )  ;
assign n17545 =  ( n17544 ) & (wr )  ;
assign n17546 =  ( n17545 ) ? ( n5123 ) : ( iram_124 ) ;
assign n17547 = wr_addr[7:7] ;
assign n17548 =  ( n17547 ) == ( bv_1_0_n53 )  ;
assign n17549 =  ( wr_addr ) == ( bv_8_124_n317 )  ;
assign n17550 =  ( n17548 ) & (n17549 )  ;
assign n17551 =  ( n17550 ) & (wr )  ;
assign n17552 =  ( n17551 ) ? ( n5165 ) : ( iram_124 ) ;
assign n17553 = wr_addr[7:7] ;
assign n17554 =  ( n17553 ) == ( bv_1_0_n53 )  ;
assign n17555 =  ( wr_addr ) == ( bv_8_124_n317 )  ;
assign n17556 =  ( n17554 ) & (n17555 )  ;
assign n17557 =  ( n17556 ) & (wr )  ;
assign n17558 =  ( n17557 ) ? ( n5204 ) : ( iram_124 ) ;
assign n17559 = wr_addr[7:7] ;
assign n17560 =  ( n17559 ) == ( bv_1_0_n53 )  ;
assign n17561 =  ( wr_addr ) == ( bv_8_124_n317 )  ;
assign n17562 =  ( n17560 ) & (n17561 )  ;
assign n17563 =  ( n17562 ) & (wr )  ;
assign n17564 =  ( n17563 ) ? ( n5262 ) : ( iram_124 ) ;
assign n17565 = wr_addr[7:7] ;
assign n17566 =  ( n17565 ) == ( bv_1_0_n53 )  ;
assign n17567 =  ( wr_addr ) == ( bv_8_124_n317 )  ;
assign n17568 =  ( n17566 ) & (n17567 )  ;
assign n17569 =  ( n17568 ) & (wr )  ;
assign n17570 =  ( n17569 ) ? ( n5298 ) : ( iram_124 ) ;
assign n17571 = wr_addr[7:7] ;
assign n17572 =  ( n17571 ) == ( bv_1_0_n53 )  ;
assign n17573 =  ( wr_addr ) == ( bv_8_124_n317 )  ;
assign n17574 =  ( n17572 ) & (n17573 )  ;
assign n17575 =  ( n17574 ) & (wr )  ;
assign n17576 =  ( n17575 ) ? ( n5325 ) : ( iram_124 ) ;
assign n17577 = wr_addr[7:7] ;
assign n17578 =  ( n17577 ) == ( bv_1_0_n53 )  ;
assign n17579 =  ( wr_addr ) == ( bv_8_125_n319 )  ;
assign n17580 =  ( n17578 ) & (n17579 )  ;
assign n17581 =  ( n17580 ) & (wr )  ;
assign n17582 =  ( n17581 ) ? ( n4782 ) : ( iram_125 ) ;
assign n17583 = wr_addr[7:7] ;
assign n17584 =  ( n17583 ) == ( bv_1_0_n53 )  ;
assign n17585 =  ( wr_addr ) == ( bv_8_125_n319 )  ;
assign n17586 =  ( n17584 ) & (n17585 )  ;
assign n17587 =  ( n17586 ) & (wr )  ;
assign n17588 =  ( n17587 ) ? ( n4841 ) : ( iram_125 ) ;
assign n17589 = wr_addr[7:7] ;
assign n17590 =  ( n17589 ) == ( bv_1_0_n53 )  ;
assign n17591 =  ( wr_addr ) == ( bv_8_125_n319 )  ;
assign n17592 =  ( n17590 ) & (n17591 )  ;
assign n17593 =  ( n17592 ) & (wr )  ;
assign n17594 =  ( n17593 ) ? ( n5449 ) : ( iram_125 ) ;
assign n17595 = wr_addr[7:7] ;
assign n17596 =  ( n17595 ) == ( bv_1_0_n53 )  ;
assign n17597 =  ( wr_addr ) == ( bv_8_125_n319 )  ;
assign n17598 =  ( n17596 ) & (n17597 )  ;
assign n17599 =  ( n17598 ) & (wr )  ;
assign n17600 =  ( n17599 ) ? ( n4906 ) : ( iram_125 ) ;
assign n17601 = wr_addr[7:7] ;
assign n17602 =  ( n17601 ) == ( bv_1_0_n53 )  ;
assign n17603 =  ( wr_addr ) == ( bv_8_125_n319 )  ;
assign n17604 =  ( n17602 ) & (n17603 )  ;
assign n17605 =  ( n17604 ) & (wr )  ;
assign n17606 =  ( n17605 ) ? ( n5485 ) : ( iram_125 ) ;
assign n17607 = wr_addr[7:7] ;
assign n17608 =  ( n17607 ) == ( bv_1_0_n53 )  ;
assign n17609 =  ( wr_addr ) == ( bv_8_125_n319 )  ;
assign n17610 =  ( n17608 ) & (n17609 )  ;
assign n17611 =  ( n17610 ) & (wr )  ;
assign n17612 =  ( n17611 ) ? ( n5512 ) : ( iram_125 ) ;
assign n17613 = wr_addr[7:7] ;
assign n17614 =  ( n17613 ) == ( bv_1_0_n53 )  ;
assign n17615 =  ( wr_addr ) == ( bv_8_125_n319 )  ;
assign n17616 =  ( n17614 ) & (n17615 )  ;
assign n17617 =  ( n17616 ) & (wr )  ;
assign n17618 =  ( n17617 ) ? ( bv_8_0_n69 ) : ( iram_125 ) ;
assign n17619 = wr_addr[7:7] ;
assign n17620 =  ( n17619 ) == ( bv_1_0_n53 )  ;
assign n17621 =  ( wr_addr ) == ( bv_8_125_n319 )  ;
assign n17622 =  ( n17620 ) & (n17621 )  ;
assign n17623 =  ( n17622 ) & (wr )  ;
assign n17624 =  ( n17623 ) ? ( n5071 ) : ( iram_125 ) ;
assign n17625 = wr_addr[7:7] ;
assign n17626 =  ( n17625 ) == ( bv_1_0_n53 )  ;
assign n17627 =  ( wr_addr ) == ( bv_8_125_n319 )  ;
assign n17628 =  ( n17626 ) & (n17627 )  ;
assign n17629 =  ( n17628 ) & (wr )  ;
assign n17630 =  ( n17629 ) ? ( n5096 ) : ( iram_125 ) ;
assign n17631 = wr_addr[7:7] ;
assign n17632 =  ( n17631 ) == ( bv_1_0_n53 )  ;
assign n17633 =  ( wr_addr ) == ( bv_8_125_n319 )  ;
assign n17634 =  ( n17632 ) & (n17633 )  ;
assign n17635 =  ( n17634 ) & (wr )  ;
assign n17636 =  ( n17635 ) ? ( n5123 ) : ( iram_125 ) ;
assign n17637 = wr_addr[7:7] ;
assign n17638 =  ( n17637 ) == ( bv_1_0_n53 )  ;
assign n17639 =  ( wr_addr ) == ( bv_8_125_n319 )  ;
assign n17640 =  ( n17638 ) & (n17639 )  ;
assign n17641 =  ( n17640 ) & (wr )  ;
assign n17642 =  ( n17641 ) ? ( n5165 ) : ( iram_125 ) ;
assign n17643 = wr_addr[7:7] ;
assign n17644 =  ( n17643 ) == ( bv_1_0_n53 )  ;
assign n17645 =  ( wr_addr ) == ( bv_8_125_n319 )  ;
assign n17646 =  ( n17644 ) & (n17645 )  ;
assign n17647 =  ( n17646 ) & (wr )  ;
assign n17648 =  ( n17647 ) ? ( n5204 ) : ( iram_125 ) ;
assign n17649 = wr_addr[7:7] ;
assign n17650 =  ( n17649 ) == ( bv_1_0_n53 )  ;
assign n17651 =  ( wr_addr ) == ( bv_8_125_n319 )  ;
assign n17652 =  ( n17650 ) & (n17651 )  ;
assign n17653 =  ( n17652 ) & (wr )  ;
assign n17654 =  ( n17653 ) ? ( n5262 ) : ( iram_125 ) ;
assign n17655 = wr_addr[7:7] ;
assign n17656 =  ( n17655 ) == ( bv_1_0_n53 )  ;
assign n17657 =  ( wr_addr ) == ( bv_8_125_n319 )  ;
assign n17658 =  ( n17656 ) & (n17657 )  ;
assign n17659 =  ( n17658 ) & (wr )  ;
assign n17660 =  ( n17659 ) ? ( n5298 ) : ( iram_125 ) ;
assign n17661 = wr_addr[7:7] ;
assign n17662 =  ( n17661 ) == ( bv_1_0_n53 )  ;
assign n17663 =  ( wr_addr ) == ( bv_8_125_n319 )  ;
assign n17664 =  ( n17662 ) & (n17663 )  ;
assign n17665 =  ( n17664 ) & (wr )  ;
assign n17666 =  ( n17665 ) ? ( n5325 ) : ( iram_125 ) ;
assign n17667 = wr_addr[7:7] ;
assign n17668 =  ( n17667 ) == ( bv_1_0_n53 )  ;
assign n17669 =  ( wr_addr ) == ( bv_8_126_n321 )  ;
assign n17670 =  ( n17668 ) & (n17669 )  ;
assign n17671 =  ( n17670 ) & (wr )  ;
assign n17672 =  ( n17671 ) ? ( n4782 ) : ( iram_126 ) ;
assign n17673 = wr_addr[7:7] ;
assign n17674 =  ( n17673 ) == ( bv_1_0_n53 )  ;
assign n17675 =  ( wr_addr ) == ( bv_8_126_n321 )  ;
assign n17676 =  ( n17674 ) & (n17675 )  ;
assign n17677 =  ( n17676 ) & (wr )  ;
assign n17678 =  ( n17677 ) ? ( n4841 ) : ( iram_126 ) ;
assign n17679 = wr_addr[7:7] ;
assign n17680 =  ( n17679 ) == ( bv_1_0_n53 )  ;
assign n17681 =  ( wr_addr ) == ( bv_8_126_n321 )  ;
assign n17682 =  ( n17680 ) & (n17681 )  ;
assign n17683 =  ( n17682 ) & (wr )  ;
assign n17684 =  ( n17683 ) ? ( n5449 ) : ( iram_126 ) ;
assign n17685 = wr_addr[7:7] ;
assign n17686 =  ( n17685 ) == ( bv_1_0_n53 )  ;
assign n17687 =  ( wr_addr ) == ( bv_8_126_n321 )  ;
assign n17688 =  ( n17686 ) & (n17687 )  ;
assign n17689 =  ( n17688 ) & (wr )  ;
assign n17690 =  ( n17689 ) ? ( n4906 ) : ( iram_126 ) ;
assign n17691 = wr_addr[7:7] ;
assign n17692 =  ( n17691 ) == ( bv_1_0_n53 )  ;
assign n17693 =  ( wr_addr ) == ( bv_8_126_n321 )  ;
assign n17694 =  ( n17692 ) & (n17693 )  ;
assign n17695 =  ( n17694 ) & (wr )  ;
assign n17696 =  ( n17695 ) ? ( n5485 ) : ( iram_126 ) ;
assign n17697 = wr_addr[7:7] ;
assign n17698 =  ( n17697 ) == ( bv_1_0_n53 )  ;
assign n17699 =  ( wr_addr ) == ( bv_8_126_n321 )  ;
assign n17700 =  ( n17698 ) & (n17699 )  ;
assign n17701 =  ( n17700 ) & (wr )  ;
assign n17702 =  ( n17701 ) ? ( n5512 ) : ( iram_126 ) ;
assign n17703 = wr_addr[7:7] ;
assign n17704 =  ( n17703 ) == ( bv_1_0_n53 )  ;
assign n17705 =  ( wr_addr ) == ( bv_8_126_n321 )  ;
assign n17706 =  ( n17704 ) & (n17705 )  ;
assign n17707 =  ( n17706 ) & (wr )  ;
assign n17708 =  ( n17707 ) ? ( bv_8_0_n69 ) : ( iram_126 ) ;
assign n17709 = wr_addr[7:7] ;
assign n17710 =  ( n17709 ) == ( bv_1_0_n53 )  ;
assign n17711 =  ( wr_addr ) == ( bv_8_126_n321 )  ;
assign n17712 =  ( n17710 ) & (n17711 )  ;
assign n17713 =  ( n17712 ) & (wr )  ;
assign n17714 =  ( n17713 ) ? ( n5071 ) : ( iram_126 ) ;
assign n17715 = wr_addr[7:7] ;
assign n17716 =  ( n17715 ) == ( bv_1_0_n53 )  ;
assign n17717 =  ( wr_addr ) == ( bv_8_126_n321 )  ;
assign n17718 =  ( n17716 ) & (n17717 )  ;
assign n17719 =  ( n17718 ) & (wr )  ;
assign n17720 =  ( n17719 ) ? ( n5096 ) : ( iram_126 ) ;
assign n17721 = wr_addr[7:7] ;
assign n17722 =  ( n17721 ) == ( bv_1_0_n53 )  ;
assign n17723 =  ( wr_addr ) == ( bv_8_126_n321 )  ;
assign n17724 =  ( n17722 ) & (n17723 )  ;
assign n17725 =  ( n17724 ) & (wr )  ;
assign n17726 =  ( n17725 ) ? ( n5123 ) : ( iram_126 ) ;
assign n17727 = wr_addr[7:7] ;
assign n17728 =  ( n17727 ) == ( bv_1_0_n53 )  ;
assign n17729 =  ( wr_addr ) == ( bv_8_126_n321 )  ;
assign n17730 =  ( n17728 ) & (n17729 )  ;
assign n17731 =  ( n17730 ) & (wr )  ;
assign n17732 =  ( n17731 ) ? ( n5165 ) : ( iram_126 ) ;
assign n17733 = wr_addr[7:7] ;
assign n17734 =  ( n17733 ) == ( bv_1_0_n53 )  ;
assign n17735 =  ( wr_addr ) == ( bv_8_126_n321 )  ;
assign n17736 =  ( n17734 ) & (n17735 )  ;
assign n17737 =  ( n17736 ) & (wr )  ;
assign n17738 =  ( n17737 ) ? ( n5204 ) : ( iram_126 ) ;
assign n17739 = wr_addr[7:7] ;
assign n17740 =  ( n17739 ) == ( bv_1_0_n53 )  ;
assign n17741 =  ( wr_addr ) == ( bv_8_126_n321 )  ;
assign n17742 =  ( n17740 ) & (n17741 )  ;
assign n17743 =  ( n17742 ) & (wr )  ;
assign n17744 =  ( n17743 ) ? ( n5262 ) : ( iram_126 ) ;
assign n17745 = wr_addr[7:7] ;
assign n17746 =  ( n17745 ) == ( bv_1_0_n53 )  ;
assign n17747 =  ( wr_addr ) == ( bv_8_126_n321 )  ;
assign n17748 =  ( n17746 ) & (n17747 )  ;
assign n17749 =  ( n17748 ) & (wr )  ;
assign n17750 =  ( n17749 ) ? ( n5298 ) : ( iram_126 ) ;
assign n17751 = wr_addr[7:7] ;
assign n17752 =  ( n17751 ) == ( bv_1_0_n53 )  ;
assign n17753 =  ( wr_addr ) == ( bv_8_126_n321 )  ;
assign n17754 =  ( n17752 ) & (n17753 )  ;
assign n17755 =  ( n17754 ) & (wr )  ;
assign n17756 =  ( n17755 ) ? ( n5325 ) : ( iram_126 ) ;
assign n17757 = wr_addr[7:7] ;
assign n17758 =  ( n17757 ) == ( bv_1_0_n53 )  ;
assign n17759 =  ( wr_addr ) == ( bv_8_127_n323 )  ;
assign n17760 =  ( n17758 ) & (n17759 )  ;
assign n17761 =  ( n17760 ) & (wr )  ;
assign n17762 =  ( n17761 ) ? ( n4782 ) : ( iram_127 ) ;
assign n17763 = wr_addr[7:7] ;
assign n17764 =  ( n17763 ) == ( bv_1_0_n53 )  ;
assign n17765 =  ( wr_addr ) == ( bv_8_127_n323 )  ;
assign n17766 =  ( n17764 ) & (n17765 )  ;
assign n17767 =  ( n17766 ) & (wr )  ;
assign n17768 =  ( n17767 ) ? ( n4841 ) : ( iram_127 ) ;
assign n17769 = wr_addr[7:7] ;
assign n17770 =  ( n17769 ) == ( bv_1_0_n53 )  ;
assign n17771 =  ( wr_addr ) == ( bv_8_127_n323 )  ;
assign n17772 =  ( n17770 ) & (n17771 )  ;
assign n17773 =  ( n17772 ) & (wr )  ;
assign n17774 =  ( n17773 ) ? ( n5449 ) : ( iram_127 ) ;
assign n17775 = wr_addr[7:7] ;
assign n17776 =  ( n17775 ) == ( bv_1_0_n53 )  ;
assign n17777 =  ( wr_addr ) == ( bv_8_127_n323 )  ;
assign n17778 =  ( n17776 ) & (n17777 )  ;
assign n17779 =  ( n17778 ) & (wr )  ;
assign n17780 =  ( n17779 ) ? ( n4906 ) : ( iram_127 ) ;
assign n17781 = wr_addr[7:7] ;
assign n17782 =  ( n17781 ) == ( bv_1_0_n53 )  ;
assign n17783 =  ( wr_addr ) == ( bv_8_127_n323 )  ;
assign n17784 =  ( n17782 ) & (n17783 )  ;
assign n17785 =  ( n17784 ) & (wr )  ;
assign n17786 =  ( n17785 ) ? ( n5485 ) : ( iram_127 ) ;
assign n17787 = wr_addr[7:7] ;
assign n17788 =  ( n17787 ) == ( bv_1_0_n53 )  ;
assign n17789 =  ( wr_addr ) == ( bv_8_127_n323 )  ;
assign n17790 =  ( n17788 ) & (n17789 )  ;
assign n17791 =  ( n17790 ) & (wr )  ;
assign n17792 =  ( n17791 ) ? ( n5512 ) : ( iram_127 ) ;
assign n17793 = wr_addr[7:7] ;
assign n17794 =  ( n17793 ) == ( bv_1_0_n53 )  ;
assign n17795 =  ( wr_addr ) == ( bv_8_127_n323 )  ;
assign n17796 =  ( n17794 ) & (n17795 )  ;
assign n17797 =  ( n17796 ) & (wr )  ;
assign n17798 =  ( n17797 ) ? ( bv_8_0_n69 ) : ( iram_127 ) ;
assign n17799 = wr_addr[7:7] ;
assign n17800 =  ( n17799 ) == ( bv_1_0_n53 )  ;
assign n17801 =  ( wr_addr ) == ( bv_8_127_n323 )  ;
assign n17802 =  ( n17800 ) & (n17801 )  ;
assign n17803 =  ( n17802 ) & (wr )  ;
assign n17804 =  ( n17803 ) ? ( n5071 ) : ( iram_127 ) ;
assign n17805 = wr_addr[7:7] ;
assign n17806 =  ( n17805 ) == ( bv_1_0_n53 )  ;
assign n17807 =  ( wr_addr ) == ( bv_8_127_n323 )  ;
assign n17808 =  ( n17806 ) & (n17807 )  ;
assign n17809 =  ( n17808 ) & (wr )  ;
assign n17810 =  ( n17809 ) ? ( n5096 ) : ( iram_127 ) ;
assign n17811 = wr_addr[7:7] ;
assign n17812 =  ( n17811 ) == ( bv_1_0_n53 )  ;
assign n17813 =  ( wr_addr ) == ( bv_8_127_n323 )  ;
assign n17814 =  ( n17812 ) & (n17813 )  ;
assign n17815 =  ( n17814 ) & (wr )  ;
assign n17816 =  ( n17815 ) ? ( n5123 ) : ( iram_127 ) ;
assign n17817 = wr_addr[7:7] ;
assign n17818 =  ( n17817 ) == ( bv_1_0_n53 )  ;
assign n17819 =  ( wr_addr ) == ( bv_8_127_n323 )  ;
assign n17820 =  ( n17818 ) & (n17819 )  ;
assign n17821 =  ( n17820 ) & (wr )  ;
assign n17822 =  ( n17821 ) ? ( n5165 ) : ( iram_127 ) ;
assign n17823 = wr_addr[7:7] ;
assign n17824 =  ( n17823 ) == ( bv_1_0_n53 )  ;
assign n17825 =  ( wr_addr ) == ( bv_8_127_n323 )  ;
assign n17826 =  ( n17824 ) & (n17825 )  ;
assign n17827 =  ( n17826 ) & (wr )  ;
assign n17828 =  ( n17827 ) ? ( n5204 ) : ( iram_127 ) ;
assign n17829 = wr_addr[7:7] ;
assign n17830 =  ( n17829 ) == ( bv_1_0_n53 )  ;
assign n17831 =  ( wr_addr ) == ( bv_8_127_n323 )  ;
assign n17832 =  ( n17830 ) & (n17831 )  ;
assign n17833 =  ( n17832 ) & (wr )  ;
assign n17834 =  ( n17833 ) ? ( n5262 ) : ( iram_127 ) ;
assign n17835 = wr_addr[7:7] ;
assign n17836 =  ( n17835 ) == ( bv_1_0_n53 )  ;
assign n17837 =  ( wr_addr ) == ( bv_8_127_n323 )  ;
assign n17838 =  ( n17836 ) & (n17837 )  ;
assign n17839 =  ( n17838 ) & (wr )  ;
assign n17840 =  ( n17839 ) ? ( n5298 ) : ( iram_127 ) ;
assign n17841 = wr_addr[7:7] ;
assign n17842 =  ( n17841 ) == ( bv_1_0_n53 )  ;
assign n17843 =  ( wr_addr ) == ( bv_8_127_n323 )  ;
assign n17844 =  ( n17842 ) & (n17843 )  ;
assign n17845 =  ( n17844 ) & (wr )  ;
assign n17846 =  ( n17845 ) ? ( n5325 ) : ( iram_127 ) ;
assign n17847 = wr_addr[7:7] ;
assign n17848 =  ( n17847 ) == ( bv_1_0_n53 )  ;
assign n17849 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n17850 =  ( n17848 ) & (n17849 )  ;
assign n17851 =  ( n17850 ) & (wr )  ;
assign n17852 =  ( n17851 ) ? ( n4782 ) : ( iram_128 ) ;
assign n17853 = wr_addr[7:7] ;
assign n17854 =  ( n17853 ) == ( bv_1_0_n53 )  ;
assign n17855 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n17856 =  ( n17854 ) & (n17855 )  ;
assign n17857 =  ( n17856 ) & (wr )  ;
assign n17858 =  ( n17857 ) ? ( n4841 ) : ( iram_128 ) ;
assign n17859 = wr_addr[7:7] ;
assign n17860 =  ( n17859 ) == ( bv_1_0_n53 )  ;
assign n17861 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n17862 =  ( n17860 ) & (n17861 )  ;
assign n17863 =  ( n17862 ) & (wr )  ;
assign n17864 =  ( n17863 ) ? ( n5449 ) : ( iram_128 ) ;
assign n17865 = wr_addr[7:7] ;
assign n17866 =  ( n17865 ) == ( bv_1_0_n53 )  ;
assign n17867 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n17868 =  ( n17866 ) & (n17867 )  ;
assign n17869 =  ( n17868 ) & (wr )  ;
assign n17870 =  ( n17869 ) ? ( n4906 ) : ( iram_128 ) ;
assign n17871 = wr_addr[7:7] ;
assign n17872 =  ( n17871 ) == ( bv_1_0_n53 )  ;
assign n17873 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n17874 =  ( n17872 ) & (n17873 )  ;
assign n17875 =  ( n17874 ) & (wr )  ;
assign n17876 =  ( n17875 ) ? ( n5485 ) : ( iram_128 ) ;
assign n17877 = wr_addr[7:7] ;
assign n17878 =  ( n17877 ) == ( bv_1_0_n53 )  ;
assign n17879 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n17880 =  ( n17878 ) & (n17879 )  ;
assign n17881 =  ( n17880 ) & (wr )  ;
assign n17882 =  ( n17881 ) ? ( n5512 ) : ( iram_128 ) ;
assign n17883 = wr_addr[7:7] ;
assign n17884 =  ( n17883 ) == ( bv_1_0_n53 )  ;
assign n17885 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n17886 =  ( n17884 ) & (n17885 )  ;
assign n17887 =  ( n17886 ) & (wr )  ;
assign n17888 =  ( n17887 ) ? ( bv_8_0_n69 ) : ( iram_128 ) ;
assign n17889 = wr_addr[7:7] ;
assign n17890 =  ( n17889 ) == ( bv_1_0_n53 )  ;
assign n17891 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n17892 =  ( n17890 ) & (n17891 )  ;
assign n17893 =  ( n17892 ) & (wr )  ;
assign n17894 =  ( n17893 ) ? ( n5071 ) : ( iram_128 ) ;
assign n17895 = wr_addr[7:7] ;
assign n17896 =  ( n17895 ) == ( bv_1_0_n53 )  ;
assign n17897 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n17898 =  ( n17896 ) & (n17897 )  ;
assign n17899 =  ( n17898 ) & (wr )  ;
assign n17900 =  ( n17899 ) ? ( n5096 ) : ( iram_128 ) ;
assign n17901 = wr_addr[7:7] ;
assign n17902 =  ( n17901 ) == ( bv_1_0_n53 )  ;
assign n17903 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n17904 =  ( n17902 ) & (n17903 )  ;
assign n17905 =  ( n17904 ) & (wr )  ;
assign n17906 =  ( n17905 ) ? ( n5123 ) : ( iram_128 ) ;
assign n17907 = wr_addr[7:7] ;
assign n17908 =  ( n17907 ) == ( bv_1_0_n53 )  ;
assign n17909 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n17910 =  ( n17908 ) & (n17909 )  ;
assign n17911 =  ( n17910 ) & (wr )  ;
assign n17912 =  ( n17911 ) ? ( n5165 ) : ( iram_128 ) ;
assign n17913 = wr_addr[7:7] ;
assign n17914 =  ( n17913 ) == ( bv_1_0_n53 )  ;
assign n17915 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n17916 =  ( n17914 ) & (n17915 )  ;
assign n17917 =  ( n17916 ) & (wr )  ;
assign n17918 =  ( n17917 ) ? ( n5204 ) : ( iram_128 ) ;
assign n17919 = wr_addr[7:7] ;
assign n17920 =  ( n17919 ) == ( bv_1_0_n53 )  ;
assign n17921 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n17922 =  ( n17920 ) & (n17921 )  ;
assign n17923 =  ( n17922 ) & (wr )  ;
assign n17924 =  ( n17923 ) ? ( n5262 ) : ( iram_128 ) ;
assign n17925 = wr_addr[7:7] ;
assign n17926 =  ( n17925 ) == ( bv_1_0_n53 )  ;
assign n17927 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n17928 =  ( n17926 ) & (n17927 )  ;
assign n17929 =  ( n17928 ) & (wr )  ;
assign n17930 =  ( n17929 ) ? ( n5298 ) : ( iram_128 ) ;
assign n17931 = wr_addr[7:7] ;
assign n17932 =  ( n17931 ) == ( bv_1_0_n53 )  ;
assign n17933 =  ( wr_addr ) == ( bv_8_128_n325 )  ;
assign n17934 =  ( n17932 ) & (n17933 )  ;
assign n17935 =  ( n17934 ) & (wr )  ;
assign n17936 =  ( n17935 ) ? ( n5325 ) : ( iram_128 ) ;
assign n17937 = wr_addr[7:7] ;
assign n17938 =  ( n17937 ) == ( bv_1_0_n53 )  ;
assign n17939 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n17940 =  ( n17938 ) & (n17939 )  ;
assign n17941 =  ( n17940 ) & (wr )  ;
assign n17942 =  ( n17941 ) ? ( n4782 ) : ( iram_129 ) ;
assign n17943 = wr_addr[7:7] ;
assign n17944 =  ( n17943 ) == ( bv_1_0_n53 )  ;
assign n17945 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n17946 =  ( n17944 ) & (n17945 )  ;
assign n17947 =  ( n17946 ) & (wr )  ;
assign n17948 =  ( n17947 ) ? ( n4841 ) : ( iram_129 ) ;
assign n17949 = wr_addr[7:7] ;
assign n17950 =  ( n17949 ) == ( bv_1_0_n53 )  ;
assign n17951 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n17952 =  ( n17950 ) & (n17951 )  ;
assign n17953 =  ( n17952 ) & (wr )  ;
assign n17954 =  ( n17953 ) ? ( n5449 ) : ( iram_129 ) ;
assign n17955 = wr_addr[7:7] ;
assign n17956 =  ( n17955 ) == ( bv_1_0_n53 )  ;
assign n17957 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n17958 =  ( n17956 ) & (n17957 )  ;
assign n17959 =  ( n17958 ) & (wr )  ;
assign n17960 =  ( n17959 ) ? ( n4906 ) : ( iram_129 ) ;
assign n17961 = wr_addr[7:7] ;
assign n17962 =  ( n17961 ) == ( bv_1_0_n53 )  ;
assign n17963 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n17964 =  ( n17962 ) & (n17963 )  ;
assign n17965 =  ( n17964 ) & (wr )  ;
assign n17966 =  ( n17965 ) ? ( n5485 ) : ( iram_129 ) ;
assign n17967 = wr_addr[7:7] ;
assign n17968 =  ( n17967 ) == ( bv_1_0_n53 )  ;
assign n17969 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n17970 =  ( n17968 ) & (n17969 )  ;
assign n17971 =  ( n17970 ) & (wr )  ;
assign n17972 =  ( n17971 ) ? ( n5512 ) : ( iram_129 ) ;
assign n17973 = wr_addr[7:7] ;
assign n17974 =  ( n17973 ) == ( bv_1_0_n53 )  ;
assign n17975 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n17976 =  ( n17974 ) & (n17975 )  ;
assign n17977 =  ( n17976 ) & (wr )  ;
assign n17978 =  ( n17977 ) ? ( bv_8_0_n69 ) : ( iram_129 ) ;
assign n17979 = wr_addr[7:7] ;
assign n17980 =  ( n17979 ) == ( bv_1_0_n53 )  ;
assign n17981 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n17982 =  ( n17980 ) & (n17981 )  ;
assign n17983 =  ( n17982 ) & (wr )  ;
assign n17984 =  ( n17983 ) ? ( n5071 ) : ( iram_129 ) ;
assign n17985 = wr_addr[7:7] ;
assign n17986 =  ( n17985 ) == ( bv_1_0_n53 )  ;
assign n17987 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n17988 =  ( n17986 ) & (n17987 )  ;
assign n17989 =  ( n17988 ) & (wr )  ;
assign n17990 =  ( n17989 ) ? ( n5096 ) : ( iram_129 ) ;
assign n17991 = wr_addr[7:7] ;
assign n17992 =  ( n17991 ) == ( bv_1_0_n53 )  ;
assign n17993 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n17994 =  ( n17992 ) & (n17993 )  ;
assign n17995 =  ( n17994 ) & (wr )  ;
assign n17996 =  ( n17995 ) ? ( n5123 ) : ( iram_129 ) ;
assign n17997 = wr_addr[7:7] ;
assign n17998 =  ( n17997 ) == ( bv_1_0_n53 )  ;
assign n17999 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n18000 =  ( n17998 ) & (n17999 )  ;
assign n18001 =  ( n18000 ) & (wr )  ;
assign n18002 =  ( n18001 ) ? ( n5165 ) : ( iram_129 ) ;
assign n18003 = wr_addr[7:7] ;
assign n18004 =  ( n18003 ) == ( bv_1_0_n53 )  ;
assign n18005 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n18006 =  ( n18004 ) & (n18005 )  ;
assign n18007 =  ( n18006 ) & (wr )  ;
assign n18008 =  ( n18007 ) ? ( n5204 ) : ( iram_129 ) ;
assign n18009 = wr_addr[7:7] ;
assign n18010 =  ( n18009 ) == ( bv_1_0_n53 )  ;
assign n18011 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n18012 =  ( n18010 ) & (n18011 )  ;
assign n18013 =  ( n18012 ) & (wr )  ;
assign n18014 =  ( n18013 ) ? ( n5262 ) : ( iram_129 ) ;
assign n18015 = wr_addr[7:7] ;
assign n18016 =  ( n18015 ) == ( bv_1_0_n53 )  ;
assign n18017 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n18018 =  ( n18016 ) & (n18017 )  ;
assign n18019 =  ( n18018 ) & (wr )  ;
assign n18020 =  ( n18019 ) ? ( n5298 ) : ( iram_129 ) ;
assign n18021 = wr_addr[7:7] ;
assign n18022 =  ( n18021 ) == ( bv_1_0_n53 )  ;
assign n18023 =  ( wr_addr ) == ( bv_8_129_n327 )  ;
assign n18024 =  ( n18022 ) & (n18023 )  ;
assign n18025 =  ( n18024 ) & (wr )  ;
assign n18026 =  ( n18025 ) ? ( n5325 ) : ( iram_129 ) ;
assign n18027 = wr_addr[7:7] ;
assign n18028 =  ( n18027 ) == ( bv_1_0_n53 )  ;
assign n18029 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n18030 =  ( n18028 ) & (n18029 )  ;
assign n18031 =  ( n18030 ) & (wr )  ;
assign n18032 =  ( n18031 ) ? ( n4782 ) : ( iram_130 ) ;
assign n18033 = wr_addr[7:7] ;
assign n18034 =  ( n18033 ) == ( bv_1_0_n53 )  ;
assign n18035 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n18036 =  ( n18034 ) & (n18035 )  ;
assign n18037 =  ( n18036 ) & (wr )  ;
assign n18038 =  ( n18037 ) ? ( n4841 ) : ( iram_130 ) ;
assign n18039 = wr_addr[7:7] ;
assign n18040 =  ( n18039 ) == ( bv_1_0_n53 )  ;
assign n18041 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n18042 =  ( n18040 ) & (n18041 )  ;
assign n18043 =  ( n18042 ) & (wr )  ;
assign n18044 =  ( n18043 ) ? ( n5449 ) : ( iram_130 ) ;
assign n18045 = wr_addr[7:7] ;
assign n18046 =  ( n18045 ) == ( bv_1_0_n53 )  ;
assign n18047 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n18048 =  ( n18046 ) & (n18047 )  ;
assign n18049 =  ( n18048 ) & (wr )  ;
assign n18050 =  ( n18049 ) ? ( n4906 ) : ( iram_130 ) ;
assign n18051 = wr_addr[7:7] ;
assign n18052 =  ( n18051 ) == ( bv_1_0_n53 )  ;
assign n18053 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n18054 =  ( n18052 ) & (n18053 )  ;
assign n18055 =  ( n18054 ) & (wr )  ;
assign n18056 =  ( n18055 ) ? ( n5485 ) : ( iram_130 ) ;
assign n18057 = wr_addr[7:7] ;
assign n18058 =  ( n18057 ) == ( bv_1_0_n53 )  ;
assign n18059 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n18060 =  ( n18058 ) & (n18059 )  ;
assign n18061 =  ( n18060 ) & (wr )  ;
assign n18062 =  ( n18061 ) ? ( n5512 ) : ( iram_130 ) ;
assign n18063 = wr_addr[7:7] ;
assign n18064 =  ( n18063 ) == ( bv_1_0_n53 )  ;
assign n18065 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n18066 =  ( n18064 ) & (n18065 )  ;
assign n18067 =  ( n18066 ) & (wr )  ;
assign n18068 =  ( n18067 ) ? ( bv_8_0_n69 ) : ( iram_130 ) ;
assign n18069 = wr_addr[7:7] ;
assign n18070 =  ( n18069 ) == ( bv_1_0_n53 )  ;
assign n18071 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n18072 =  ( n18070 ) & (n18071 )  ;
assign n18073 =  ( n18072 ) & (wr )  ;
assign n18074 =  ( n18073 ) ? ( n5071 ) : ( iram_130 ) ;
assign n18075 = wr_addr[7:7] ;
assign n18076 =  ( n18075 ) == ( bv_1_0_n53 )  ;
assign n18077 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n18078 =  ( n18076 ) & (n18077 )  ;
assign n18079 =  ( n18078 ) & (wr )  ;
assign n18080 =  ( n18079 ) ? ( n5096 ) : ( iram_130 ) ;
assign n18081 = wr_addr[7:7] ;
assign n18082 =  ( n18081 ) == ( bv_1_0_n53 )  ;
assign n18083 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n18084 =  ( n18082 ) & (n18083 )  ;
assign n18085 =  ( n18084 ) & (wr )  ;
assign n18086 =  ( n18085 ) ? ( n5123 ) : ( iram_130 ) ;
assign n18087 = wr_addr[7:7] ;
assign n18088 =  ( n18087 ) == ( bv_1_0_n53 )  ;
assign n18089 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n18090 =  ( n18088 ) & (n18089 )  ;
assign n18091 =  ( n18090 ) & (wr )  ;
assign n18092 =  ( n18091 ) ? ( n5165 ) : ( iram_130 ) ;
assign n18093 = wr_addr[7:7] ;
assign n18094 =  ( n18093 ) == ( bv_1_0_n53 )  ;
assign n18095 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n18096 =  ( n18094 ) & (n18095 )  ;
assign n18097 =  ( n18096 ) & (wr )  ;
assign n18098 =  ( n18097 ) ? ( n5204 ) : ( iram_130 ) ;
assign n18099 = wr_addr[7:7] ;
assign n18100 =  ( n18099 ) == ( bv_1_0_n53 )  ;
assign n18101 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n18102 =  ( n18100 ) & (n18101 )  ;
assign n18103 =  ( n18102 ) & (wr )  ;
assign n18104 =  ( n18103 ) ? ( n5262 ) : ( iram_130 ) ;
assign n18105 = wr_addr[7:7] ;
assign n18106 =  ( n18105 ) == ( bv_1_0_n53 )  ;
assign n18107 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n18108 =  ( n18106 ) & (n18107 )  ;
assign n18109 =  ( n18108 ) & (wr )  ;
assign n18110 =  ( n18109 ) ? ( n5298 ) : ( iram_130 ) ;
assign n18111 = wr_addr[7:7] ;
assign n18112 =  ( n18111 ) == ( bv_1_0_n53 )  ;
assign n18113 =  ( wr_addr ) == ( bv_8_130_n329 )  ;
assign n18114 =  ( n18112 ) & (n18113 )  ;
assign n18115 =  ( n18114 ) & (wr )  ;
assign n18116 =  ( n18115 ) ? ( n5325 ) : ( iram_130 ) ;
assign n18117 = wr_addr[7:7] ;
assign n18118 =  ( n18117 ) == ( bv_1_0_n53 )  ;
assign n18119 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n18120 =  ( n18118 ) & (n18119 )  ;
assign n18121 =  ( n18120 ) & (wr )  ;
assign n18122 =  ( n18121 ) ? ( n4782 ) : ( iram_131 ) ;
assign n18123 = wr_addr[7:7] ;
assign n18124 =  ( n18123 ) == ( bv_1_0_n53 )  ;
assign n18125 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n18126 =  ( n18124 ) & (n18125 )  ;
assign n18127 =  ( n18126 ) & (wr )  ;
assign n18128 =  ( n18127 ) ? ( n4841 ) : ( iram_131 ) ;
assign n18129 = wr_addr[7:7] ;
assign n18130 =  ( n18129 ) == ( bv_1_0_n53 )  ;
assign n18131 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n18132 =  ( n18130 ) & (n18131 )  ;
assign n18133 =  ( n18132 ) & (wr )  ;
assign n18134 =  ( n18133 ) ? ( n5449 ) : ( iram_131 ) ;
assign n18135 = wr_addr[7:7] ;
assign n18136 =  ( n18135 ) == ( bv_1_0_n53 )  ;
assign n18137 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n18138 =  ( n18136 ) & (n18137 )  ;
assign n18139 =  ( n18138 ) & (wr )  ;
assign n18140 =  ( n18139 ) ? ( n4906 ) : ( iram_131 ) ;
assign n18141 = wr_addr[7:7] ;
assign n18142 =  ( n18141 ) == ( bv_1_0_n53 )  ;
assign n18143 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n18144 =  ( n18142 ) & (n18143 )  ;
assign n18145 =  ( n18144 ) & (wr )  ;
assign n18146 =  ( n18145 ) ? ( n5485 ) : ( iram_131 ) ;
assign n18147 = wr_addr[7:7] ;
assign n18148 =  ( n18147 ) == ( bv_1_0_n53 )  ;
assign n18149 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n18150 =  ( n18148 ) & (n18149 )  ;
assign n18151 =  ( n18150 ) & (wr )  ;
assign n18152 =  ( n18151 ) ? ( n5512 ) : ( iram_131 ) ;
assign n18153 = wr_addr[7:7] ;
assign n18154 =  ( n18153 ) == ( bv_1_0_n53 )  ;
assign n18155 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n18156 =  ( n18154 ) & (n18155 )  ;
assign n18157 =  ( n18156 ) & (wr )  ;
assign n18158 =  ( n18157 ) ? ( bv_8_0_n69 ) : ( iram_131 ) ;
assign n18159 = wr_addr[7:7] ;
assign n18160 =  ( n18159 ) == ( bv_1_0_n53 )  ;
assign n18161 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n18162 =  ( n18160 ) & (n18161 )  ;
assign n18163 =  ( n18162 ) & (wr )  ;
assign n18164 =  ( n18163 ) ? ( n5071 ) : ( iram_131 ) ;
assign n18165 = wr_addr[7:7] ;
assign n18166 =  ( n18165 ) == ( bv_1_0_n53 )  ;
assign n18167 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n18168 =  ( n18166 ) & (n18167 )  ;
assign n18169 =  ( n18168 ) & (wr )  ;
assign n18170 =  ( n18169 ) ? ( n5096 ) : ( iram_131 ) ;
assign n18171 = wr_addr[7:7] ;
assign n18172 =  ( n18171 ) == ( bv_1_0_n53 )  ;
assign n18173 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n18174 =  ( n18172 ) & (n18173 )  ;
assign n18175 =  ( n18174 ) & (wr )  ;
assign n18176 =  ( n18175 ) ? ( n5123 ) : ( iram_131 ) ;
assign n18177 = wr_addr[7:7] ;
assign n18178 =  ( n18177 ) == ( bv_1_0_n53 )  ;
assign n18179 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n18180 =  ( n18178 ) & (n18179 )  ;
assign n18181 =  ( n18180 ) & (wr )  ;
assign n18182 =  ( n18181 ) ? ( n5165 ) : ( iram_131 ) ;
assign n18183 = wr_addr[7:7] ;
assign n18184 =  ( n18183 ) == ( bv_1_0_n53 )  ;
assign n18185 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n18186 =  ( n18184 ) & (n18185 )  ;
assign n18187 =  ( n18186 ) & (wr )  ;
assign n18188 =  ( n18187 ) ? ( n5204 ) : ( iram_131 ) ;
assign n18189 = wr_addr[7:7] ;
assign n18190 =  ( n18189 ) == ( bv_1_0_n53 )  ;
assign n18191 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n18192 =  ( n18190 ) & (n18191 )  ;
assign n18193 =  ( n18192 ) & (wr )  ;
assign n18194 =  ( n18193 ) ? ( n5262 ) : ( iram_131 ) ;
assign n18195 = wr_addr[7:7] ;
assign n18196 =  ( n18195 ) == ( bv_1_0_n53 )  ;
assign n18197 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n18198 =  ( n18196 ) & (n18197 )  ;
assign n18199 =  ( n18198 ) & (wr )  ;
assign n18200 =  ( n18199 ) ? ( n5298 ) : ( iram_131 ) ;
assign n18201 = wr_addr[7:7] ;
assign n18202 =  ( n18201 ) == ( bv_1_0_n53 )  ;
assign n18203 =  ( wr_addr ) == ( bv_8_131_n331 )  ;
assign n18204 =  ( n18202 ) & (n18203 )  ;
assign n18205 =  ( n18204 ) & (wr )  ;
assign n18206 =  ( n18205 ) ? ( n5325 ) : ( iram_131 ) ;
assign n18207 = wr_addr[7:7] ;
assign n18208 =  ( n18207 ) == ( bv_1_0_n53 )  ;
assign n18209 =  ( wr_addr ) == ( bv_8_132_n333 )  ;
assign n18210 =  ( n18208 ) & (n18209 )  ;
assign n18211 =  ( n18210 ) & (wr )  ;
assign n18212 =  ( n18211 ) ? ( n4782 ) : ( iram_132 ) ;
assign n18213 = wr_addr[7:7] ;
assign n18214 =  ( n18213 ) == ( bv_1_0_n53 )  ;
assign n18215 =  ( wr_addr ) == ( bv_8_132_n333 )  ;
assign n18216 =  ( n18214 ) & (n18215 )  ;
assign n18217 =  ( n18216 ) & (wr )  ;
assign n18218 =  ( n18217 ) ? ( n4841 ) : ( iram_132 ) ;
assign n18219 = wr_addr[7:7] ;
assign n18220 =  ( n18219 ) == ( bv_1_0_n53 )  ;
assign n18221 =  ( wr_addr ) == ( bv_8_132_n333 )  ;
assign n18222 =  ( n18220 ) & (n18221 )  ;
assign n18223 =  ( n18222 ) & (wr )  ;
assign n18224 =  ( n18223 ) ? ( n5449 ) : ( iram_132 ) ;
assign n18225 = wr_addr[7:7] ;
assign n18226 =  ( n18225 ) == ( bv_1_0_n53 )  ;
assign n18227 =  ( wr_addr ) == ( bv_8_132_n333 )  ;
assign n18228 =  ( n18226 ) & (n18227 )  ;
assign n18229 =  ( n18228 ) & (wr )  ;
assign n18230 =  ( n18229 ) ? ( n4906 ) : ( iram_132 ) ;
assign n18231 = wr_addr[7:7] ;
assign n18232 =  ( n18231 ) == ( bv_1_0_n53 )  ;
assign n18233 =  ( wr_addr ) == ( bv_8_132_n333 )  ;
assign n18234 =  ( n18232 ) & (n18233 )  ;
assign n18235 =  ( n18234 ) & (wr )  ;
assign n18236 =  ( n18235 ) ? ( n5485 ) : ( iram_132 ) ;
assign n18237 = wr_addr[7:7] ;
assign n18238 =  ( n18237 ) == ( bv_1_0_n53 )  ;
assign n18239 =  ( wr_addr ) == ( bv_8_132_n333 )  ;
assign n18240 =  ( n18238 ) & (n18239 )  ;
assign n18241 =  ( n18240 ) & (wr )  ;
assign n18242 =  ( n18241 ) ? ( n5512 ) : ( iram_132 ) ;
assign n18243 = wr_addr[7:7] ;
assign n18244 =  ( n18243 ) == ( bv_1_0_n53 )  ;
assign n18245 =  ( wr_addr ) == ( bv_8_132_n333 )  ;
assign n18246 =  ( n18244 ) & (n18245 )  ;
assign n18247 =  ( n18246 ) & (wr )  ;
assign n18248 =  ( n18247 ) ? ( bv_8_0_n69 ) : ( iram_132 ) ;
assign n18249 = wr_addr[7:7] ;
assign n18250 =  ( n18249 ) == ( bv_1_0_n53 )  ;
assign n18251 =  ( wr_addr ) == ( bv_8_132_n333 )  ;
assign n18252 =  ( n18250 ) & (n18251 )  ;
assign n18253 =  ( n18252 ) & (wr )  ;
assign n18254 =  ( n18253 ) ? ( n5071 ) : ( iram_132 ) ;
assign n18255 = wr_addr[7:7] ;
assign n18256 =  ( n18255 ) == ( bv_1_0_n53 )  ;
assign n18257 =  ( wr_addr ) == ( bv_8_132_n333 )  ;
assign n18258 =  ( n18256 ) & (n18257 )  ;
assign n18259 =  ( n18258 ) & (wr )  ;
assign n18260 =  ( n18259 ) ? ( n5096 ) : ( iram_132 ) ;
assign n18261 = wr_addr[7:7] ;
assign n18262 =  ( n18261 ) == ( bv_1_0_n53 )  ;
assign n18263 =  ( wr_addr ) == ( bv_8_132_n333 )  ;
assign n18264 =  ( n18262 ) & (n18263 )  ;
assign n18265 =  ( n18264 ) & (wr )  ;
assign n18266 =  ( n18265 ) ? ( n5123 ) : ( iram_132 ) ;
assign n18267 = wr_addr[7:7] ;
assign n18268 =  ( n18267 ) == ( bv_1_0_n53 )  ;
assign n18269 =  ( wr_addr ) == ( bv_8_132_n333 )  ;
assign n18270 =  ( n18268 ) & (n18269 )  ;
assign n18271 =  ( n18270 ) & (wr )  ;
assign n18272 =  ( n18271 ) ? ( n5165 ) : ( iram_132 ) ;
assign n18273 = wr_addr[7:7] ;
assign n18274 =  ( n18273 ) == ( bv_1_0_n53 )  ;
assign n18275 =  ( wr_addr ) == ( bv_8_132_n333 )  ;
assign n18276 =  ( n18274 ) & (n18275 )  ;
assign n18277 =  ( n18276 ) & (wr )  ;
assign n18278 =  ( n18277 ) ? ( n5204 ) : ( iram_132 ) ;
assign n18279 = wr_addr[7:7] ;
assign n18280 =  ( n18279 ) == ( bv_1_0_n53 )  ;
assign n18281 =  ( wr_addr ) == ( bv_8_132_n333 )  ;
assign n18282 =  ( n18280 ) & (n18281 )  ;
assign n18283 =  ( n18282 ) & (wr )  ;
assign n18284 =  ( n18283 ) ? ( n5262 ) : ( iram_132 ) ;
assign n18285 = wr_addr[7:7] ;
assign n18286 =  ( n18285 ) == ( bv_1_0_n53 )  ;
assign n18287 =  ( wr_addr ) == ( bv_8_132_n333 )  ;
assign n18288 =  ( n18286 ) & (n18287 )  ;
assign n18289 =  ( n18288 ) & (wr )  ;
assign n18290 =  ( n18289 ) ? ( n5298 ) : ( iram_132 ) ;
assign n18291 = wr_addr[7:7] ;
assign n18292 =  ( n18291 ) == ( bv_1_0_n53 )  ;
assign n18293 =  ( wr_addr ) == ( bv_8_132_n333 )  ;
assign n18294 =  ( n18292 ) & (n18293 )  ;
assign n18295 =  ( n18294 ) & (wr )  ;
assign n18296 =  ( n18295 ) ? ( n5325 ) : ( iram_132 ) ;
assign n18297 = wr_addr[7:7] ;
assign n18298 =  ( n18297 ) == ( bv_1_0_n53 )  ;
assign n18299 =  ( wr_addr ) == ( bv_8_133_n335 )  ;
assign n18300 =  ( n18298 ) & (n18299 )  ;
assign n18301 =  ( n18300 ) & (wr )  ;
assign n18302 =  ( n18301 ) ? ( n4782 ) : ( iram_133 ) ;
assign n18303 = wr_addr[7:7] ;
assign n18304 =  ( n18303 ) == ( bv_1_0_n53 )  ;
assign n18305 =  ( wr_addr ) == ( bv_8_133_n335 )  ;
assign n18306 =  ( n18304 ) & (n18305 )  ;
assign n18307 =  ( n18306 ) & (wr )  ;
assign n18308 =  ( n18307 ) ? ( n4841 ) : ( iram_133 ) ;
assign n18309 = wr_addr[7:7] ;
assign n18310 =  ( n18309 ) == ( bv_1_0_n53 )  ;
assign n18311 =  ( wr_addr ) == ( bv_8_133_n335 )  ;
assign n18312 =  ( n18310 ) & (n18311 )  ;
assign n18313 =  ( n18312 ) & (wr )  ;
assign n18314 =  ( n18313 ) ? ( n5449 ) : ( iram_133 ) ;
assign n18315 = wr_addr[7:7] ;
assign n18316 =  ( n18315 ) == ( bv_1_0_n53 )  ;
assign n18317 =  ( wr_addr ) == ( bv_8_133_n335 )  ;
assign n18318 =  ( n18316 ) & (n18317 )  ;
assign n18319 =  ( n18318 ) & (wr )  ;
assign n18320 =  ( n18319 ) ? ( n4906 ) : ( iram_133 ) ;
assign n18321 = wr_addr[7:7] ;
assign n18322 =  ( n18321 ) == ( bv_1_0_n53 )  ;
assign n18323 =  ( wr_addr ) == ( bv_8_133_n335 )  ;
assign n18324 =  ( n18322 ) & (n18323 )  ;
assign n18325 =  ( n18324 ) & (wr )  ;
assign n18326 =  ( n18325 ) ? ( n5485 ) : ( iram_133 ) ;
assign n18327 = wr_addr[7:7] ;
assign n18328 =  ( n18327 ) == ( bv_1_0_n53 )  ;
assign n18329 =  ( wr_addr ) == ( bv_8_133_n335 )  ;
assign n18330 =  ( n18328 ) & (n18329 )  ;
assign n18331 =  ( n18330 ) & (wr )  ;
assign n18332 =  ( n18331 ) ? ( n5512 ) : ( iram_133 ) ;
assign n18333 = wr_addr[7:7] ;
assign n18334 =  ( n18333 ) == ( bv_1_0_n53 )  ;
assign n18335 =  ( wr_addr ) == ( bv_8_133_n335 )  ;
assign n18336 =  ( n18334 ) & (n18335 )  ;
assign n18337 =  ( n18336 ) & (wr )  ;
assign n18338 =  ( n18337 ) ? ( bv_8_0_n69 ) : ( iram_133 ) ;
assign n18339 = wr_addr[7:7] ;
assign n18340 =  ( n18339 ) == ( bv_1_0_n53 )  ;
assign n18341 =  ( wr_addr ) == ( bv_8_133_n335 )  ;
assign n18342 =  ( n18340 ) & (n18341 )  ;
assign n18343 =  ( n18342 ) & (wr )  ;
assign n18344 =  ( n18343 ) ? ( n5071 ) : ( iram_133 ) ;
assign n18345 = wr_addr[7:7] ;
assign n18346 =  ( n18345 ) == ( bv_1_0_n53 )  ;
assign n18347 =  ( wr_addr ) == ( bv_8_133_n335 )  ;
assign n18348 =  ( n18346 ) & (n18347 )  ;
assign n18349 =  ( n18348 ) & (wr )  ;
assign n18350 =  ( n18349 ) ? ( n5096 ) : ( iram_133 ) ;
assign n18351 = wr_addr[7:7] ;
assign n18352 =  ( n18351 ) == ( bv_1_0_n53 )  ;
assign n18353 =  ( wr_addr ) == ( bv_8_133_n335 )  ;
assign n18354 =  ( n18352 ) & (n18353 )  ;
assign n18355 =  ( n18354 ) & (wr )  ;
assign n18356 =  ( n18355 ) ? ( n5123 ) : ( iram_133 ) ;
assign n18357 = wr_addr[7:7] ;
assign n18358 =  ( n18357 ) == ( bv_1_0_n53 )  ;
assign n18359 =  ( wr_addr ) == ( bv_8_133_n335 )  ;
assign n18360 =  ( n18358 ) & (n18359 )  ;
assign n18361 =  ( n18360 ) & (wr )  ;
assign n18362 =  ( n18361 ) ? ( n5165 ) : ( iram_133 ) ;
assign n18363 = wr_addr[7:7] ;
assign n18364 =  ( n18363 ) == ( bv_1_0_n53 )  ;
assign n18365 =  ( wr_addr ) == ( bv_8_133_n335 )  ;
assign n18366 =  ( n18364 ) & (n18365 )  ;
assign n18367 =  ( n18366 ) & (wr )  ;
assign n18368 =  ( n18367 ) ? ( n5204 ) : ( iram_133 ) ;
assign n18369 = wr_addr[7:7] ;
assign n18370 =  ( n18369 ) == ( bv_1_0_n53 )  ;
assign n18371 =  ( wr_addr ) == ( bv_8_133_n335 )  ;
assign n18372 =  ( n18370 ) & (n18371 )  ;
assign n18373 =  ( n18372 ) & (wr )  ;
assign n18374 =  ( n18373 ) ? ( n5262 ) : ( iram_133 ) ;
assign n18375 = wr_addr[7:7] ;
assign n18376 =  ( n18375 ) == ( bv_1_0_n53 )  ;
assign n18377 =  ( wr_addr ) == ( bv_8_133_n335 )  ;
assign n18378 =  ( n18376 ) & (n18377 )  ;
assign n18379 =  ( n18378 ) & (wr )  ;
assign n18380 =  ( n18379 ) ? ( n5298 ) : ( iram_133 ) ;
assign n18381 = wr_addr[7:7] ;
assign n18382 =  ( n18381 ) == ( bv_1_0_n53 )  ;
assign n18383 =  ( wr_addr ) == ( bv_8_133_n335 )  ;
assign n18384 =  ( n18382 ) & (n18383 )  ;
assign n18385 =  ( n18384 ) & (wr )  ;
assign n18386 =  ( n18385 ) ? ( n5325 ) : ( iram_133 ) ;
assign n18387 = wr_addr[7:7] ;
assign n18388 =  ( n18387 ) == ( bv_1_0_n53 )  ;
assign n18389 =  ( wr_addr ) == ( bv_8_134_n337 )  ;
assign n18390 =  ( n18388 ) & (n18389 )  ;
assign n18391 =  ( n18390 ) & (wr )  ;
assign n18392 =  ( n18391 ) ? ( n4782 ) : ( iram_134 ) ;
assign n18393 = wr_addr[7:7] ;
assign n18394 =  ( n18393 ) == ( bv_1_0_n53 )  ;
assign n18395 =  ( wr_addr ) == ( bv_8_134_n337 )  ;
assign n18396 =  ( n18394 ) & (n18395 )  ;
assign n18397 =  ( n18396 ) & (wr )  ;
assign n18398 =  ( n18397 ) ? ( n4841 ) : ( iram_134 ) ;
assign n18399 = wr_addr[7:7] ;
assign n18400 =  ( n18399 ) == ( bv_1_0_n53 )  ;
assign n18401 =  ( wr_addr ) == ( bv_8_134_n337 )  ;
assign n18402 =  ( n18400 ) & (n18401 )  ;
assign n18403 =  ( n18402 ) & (wr )  ;
assign n18404 =  ( n18403 ) ? ( n5449 ) : ( iram_134 ) ;
assign n18405 = wr_addr[7:7] ;
assign n18406 =  ( n18405 ) == ( bv_1_0_n53 )  ;
assign n18407 =  ( wr_addr ) == ( bv_8_134_n337 )  ;
assign n18408 =  ( n18406 ) & (n18407 )  ;
assign n18409 =  ( n18408 ) & (wr )  ;
assign n18410 =  ( n18409 ) ? ( n4906 ) : ( iram_134 ) ;
assign n18411 = wr_addr[7:7] ;
assign n18412 =  ( n18411 ) == ( bv_1_0_n53 )  ;
assign n18413 =  ( wr_addr ) == ( bv_8_134_n337 )  ;
assign n18414 =  ( n18412 ) & (n18413 )  ;
assign n18415 =  ( n18414 ) & (wr )  ;
assign n18416 =  ( n18415 ) ? ( n5485 ) : ( iram_134 ) ;
assign n18417 = wr_addr[7:7] ;
assign n18418 =  ( n18417 ) == ( bv_1_0_n53 )  ;
assign n18419 =  ( wr_addr ) == ( bv_8_134_n337 )  ;
assign n18420 =  ( n18418 ) & (n18419 )  ;
assign n18421 =  ( n18420 ) & (wr )  ;
assign n18422 =  ( n18421 ) ? ( n5512 ) : ( iram_134 ) ;
assign n18423 = wr_addr[7:7] ;
assign n18424 =  ( n18423 ) == ( bv_1_0_n53 )  ;
assign n18425 =  ( wr_addr ) == ( bv_8_134_n337 )  ;
assign n18426 =  ( n18424 ) & (n18425 )  ;
assign n18427 =  ( n18426 ) & (wr )  ;
assign n18428 =  ( n18427 ) ? ( bv_8_0_n69 ) : ( iram_134 ) ;
assign n18429 = wr_addr[7:7] ;
assign n18430 =  ( n18429 ) == ( bv_1_0_n53 )  ;
assign n18431 =  ( wr_addr ) == ( bv_8_134_n337 )  ;
assign n18432 =  ( n18430 ) & (n18431 )  ;
assign n18433 =  ( n18432 ) & (wr )  ;
assign n18434 =  ( n18433 ) ? ( n5071 ) : ( iram_134 ) ;
assign n18435 = wr_addr[7:7] ;
assign n18436 =  ( n18435 ) == ( bv_1_0_n53 )  ;
assign n18437 =  ( wr_addr ) == ( bv_8_134_n337 )  ;
assign n18438 =  ( n18436 ) & (n18437 )  ;
assign n18439 =  ( n18438 ) & (wr )  ;
assign n18440 =  ( n18439 ) ? ( n5096 ) : ( iram_134 ) ;
assign n18441 = wr_addr[7:7] ;
assign n18442 =  ( n18441 ) == ( bv_1_0_n53 )  ;
assign n18443 =  ( wr_addr ) == ( bv_8_134_n337 )  ;
assign n18444 =  ( n18442 ) & (n18443 )  ;
assign n18445 =  ( n18444 ) & (wr )  ;
assign n18446 =  ( n18445 ) ? ( n5123 ) : ( iram_134 ) ;
assign n18447 = wr_addr[7:7] ;
assign n18448 =  ( n18447 ) == ( bv_1_0_n53 )  ;
assign n18449 =  ( wr_addr ) == ( bv_8_134_n337 )  ;
assign n18450 =  ( n18448 ) & (n18449 )  ;
assign n18451 =  ( n18450 ) & (wr )  ;
assign n18452 =  ( n18451 ) ? ( n5165 ) : ( iram_134 ) ;
assign n18453 = wr_addr[7:7] ;
assign n18454 =  ( n18453 ) == ( bv_1_0_n53 )  ;
assign n18455 =  ( wr_addr ) == ( bv_8_134_n337 )  ;
assign n18456 =  ( n18454 ) & (n18455 )  ;
assign n18457 =  ( n18456 ) & (wr )  ;
assign n18458 =  ( n18457 ) ? ( n5204 ) : ( iram_134 ) ;
assign n18459 = wr_addr[7:7] ;
assign n18460 =  ( n18459 ) == ( bv_1_0_n53 )  ;
assign n18461 =  ( wr_addr ) == ( bv_8_134_n337 )  ;
assign n18462 =  ( n18460 ) & (n18461 )  ;
assign n18463 =  ( n18462 ) & (wr )  ;
assign n18464 =  ( n18463 ) ? ( n5262 ) : ( iram_134 ) ;
assign n18465 = wr_addr[7:7] ;
assign n18466 =  ( n18465 ) == ( bv_1_0_n53 )  ;
assign n18467 =  ( wr_addr ) == ( bv_8_134_n337 )  ;
assign n18468 =  ( n18466 ) & (n18467 )  ;
assign n18469 =  ( n18468 ) & (wr )  ;
assign n18470 =  ( n18469 ) ? ( n5298 ) : ( iram_134 ) ;
assign n18471 = wr_addr[7:7] ;
assign n18472 =  ( n18471 ) == ( bv_1_0_n53 )  ;
assign n18473 =  ( wr_addr ) == ( bv_8_134_n337 )  ;
assign n18474 =  ( n18472 ) & (n18473 )  ;
assign n18475 =  ( n18474 ) & (wr )  ;
assign n18476 =  ( n18475 ) ? ( n5325 ) : ( iram_134 ) ;
assign n18477 = wr_addr[7:7] ;
assign n18478 =  ( n18477 ) == ( bv_1_0_n53 )  ;
assign n18479 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n18480 =  ( n18478 ) & (n18479 )  ;
assign n18481 =  ( n18480 ) & (wr )  ;
assign n18482 =  ( n18481 ) ? ( n4782 ) : ( iram_135 ) ;
assign n18483 = wr_addr[7:7] ;
assign n18484 =  ( n18483 ) == ( bv_1_0_n53 )  ;
assign n18485 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n18486 =  ( n18484 ) & (n18485 )  ;
assign n18487 =  ( n18486 ) & (wr )  ;
assign n18488 =  ( n18487 ) ? ( n4841 ) : ( iram_135 ) ;
assign n18489 = wr_addr[7:7] ;
assign n18490 =  ( n18489 ) == ( bv_1_0_n53 )  ;
assign n18491 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n18492 =  ( n18490 ) & (n18491 )  ;
assign n18493 =  ( n18492 ) & (wr )  ;
assign n18494 =  ( n18493 ) ? ( n5449 ) : ( iram_135 ) ;
assign n18495 = wr_addr[7:7] ;
assign n18496 =  ( n18495 ) == ( bv_1_0_n53 )  ;
assign n18497 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n18498 =  ( n18496 ) & (n18497 )  ;
assign n18499 =  ( n18498 ) & (wr )  ;
assign n18500 =  ( n18499 ) ? ( n4906 ) : ( iram_135 ) ;
assign n18501 = wr_addr[7:7] ;
assign n18502 =  ( n18501 ) == ( bv_1_0_n53 )  ;
assign n18503 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n18504 =  ( n18502 ) & (n18503 )  ;
assign n18505 =  ( n18504 ) & (wr )  ;
assign n18506 =  ( n18505 ) ? ( n5485 ) : ( iram_135 ) ;
assign n18507 = wr_addr[7:7] ;
assign n18508 =  ( n18507 ) == ( bv_1_0_n53 )  ;
assign n18509 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n18510 =  ( n18508 ) & (n18509 )  ;
assign n18511 =  ( n18510 ) & (wr )  ;
assign n18512 =  ( n18511 ) ? ( n5512 ) : ( iram_135 ) ;
assign n18513 = wr_addr[7:7] ;
assign n18514 =  ( n18513 ) == ( bv_1_0_n53 )  ;
assign n18515 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n18516 =  ( n18514 ) & (n18515 )  ;
assign n18517 =  ( n18516 ) & (wr )  ;
assign n18518 =  ( n18517 ) ? ( bv_8_0_n69 ) : ( iram_135 ) ;
assign n18519 = wr_addr[7:7] ;
assign n18520 =  ( n18519 ) == ( bv_1_0_n53 )  ;
assign n18521 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n18522 =  ( n18520 ) & (n18521 )  ;
assign n18523 =  ( n18522 ) & (wr )  ;
assign n18524 =  ( n18523 ) ? ( n5071 ) : ( iram_135 ) ;
assign n18525 = wr_addr[7:7] ;
assign n18526 =  ( n18525 ) == ( bv_1_0_n53 )  ;
assign n18527 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n18528 =  ( n18526 ) & (n18527 )  ;
assign n18529 =  ( n18528 ) & (wr )  ;
assign n18530 =  ( n18529 ) ? ( n5096 ) : ( iram_135 ) ;
assign n18531 = wr_addr[7:7] ;
assign n18532 =  ( n18531 ) == ( bv_1_0_n53 )  ;
assign n18533 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n18534 =  ( n18532 ) & (n18533 )  ;
assign n18535 =  ( n18534 ) & (wr )  ;
assign n18536 =  ( n18535 ) ? ( n5123 ) : ( iram_135 ) ;
assign n18537 = wr_addr[7:7] ;
assign n18538 =  ( n18537 ) == ( bv_1_0_n53 )  ;
assign n18539 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n18540 =  ( n18538 ) & (n18539 )  ;
assign n18541 =  ( n18540 ) & (wr )  ;
assign n18542 =  ( n18541 ) ? ( n5165 ) : ( iram_135 ) ;
assign n18543 = wr_addr[7:7] ;
assign n18544 =  ( n18543 ) == ( bv_1_0_n53 )  ;
assign n18545 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n18546 =  ( n18544 ) & (n18545 )  ;
assign n18547 =  ( n18546 ) & (wr )  ;
assign n18548 =  ( n18547 ) ? ( n5204 ) : ( iram_135 ) ;
assign n18549 = wr_addr[7:7] ;
assign n18550 =  ( n18549 ) == ( bv_1_0_n53 )  ;
assign n18551 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n18552 =  ( n18550 ) & (n18551 )  ;
assign n18553 =  ( n18552 ) & (wr )  ;
assign n18554 =  ( n18553 ) ? ( n5262 ) : ( iram_135 ) ;
assign n18555 = wr_addr[7:7] ;
assign n18556 =  ( n18555 ) == ( bv_1_0_n53 )  ;
assign n18557 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n18558 =  ( n18556 ) & (n18557 )  ;
assign n18559 =  ( n18558 ) & (wr )  ;
assign n18560 =  ( n18559 ) ? ( n5298 ) : ( iram_135 ) ;
assign n18561 = wr_addr[7:7] ;
assign n18562 =  ( n18561 ) == ( bv_1_0_n53 )  ;
assign n18563 =  ( wr_addr ) == ( bv_8_135_n339 )  ;
assign n18564 =  ( n18562 ) & (n18563 )  ;
assign n18565 =  ( n18564 ) & (wr )  ;
assign n18566 =  ( n18565 ) ? ( n5325 ) : ( iram_135 ) ;
assign n18567 = wr_addr[7:7] ;
assign n18568 =  ( n18567 ) == ( bv_1_0_n53 )  ;
assign n18569 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n18570 =  ( n18568 ) & (n18569 )  ;
assign n18571 =  ( n18570 ) & (wr )  ;
assign n18572 =  ( n18571 ) ? ( n4782 ) : ( iram_136 ) ;
assign n18573 = wr_addr[7:7] ;
assign n18574 =  ( n18573 ) == ( bv_1_0_n53 )  ;
assign n18575 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n18576 =  ( n18574 ) & (n18575 )  ;
assign n18577 =  ( n18576 ) & (wr )  ;
assign n18578 =  ( n18577 ) ? ( n4841 ) : ( iram_136 ) ;
assign n18579 = wr_addr[7:7] ;
assign n18580 =  ( n18579 ) == ( bv_1_0_n53 )  ;
assign n18581 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n18582 =  ( n18580 ) & (n18581 )  ;
assign n18583 =  ( n18582 ) & (wr )  ;
assign n18584 =  ( n18583 ) ? ( n5449 ) : ( iram_136 ) ;
assign n18585 = wr_addr[7:7] ;
assign n18586 =  ( n18585 ) == ( bv_1_0_n53 )  ;
assign n18587 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n18588 =  ( n18586 ) & (n18587 )  ;
assign n18589 =  ( n18588 ) & (wr )  ;
assign n18590 =  ( n18589 ) ? ( n4906 ) : ( iram_136 ) ;
assign n18591 = wr_addr[7:7] ;
assign n18592 =  ( n18591 ) == ( bv_1_0_n53 )  ;
assign n18593 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n18594 =  ( n18592 ) & (n18593 )  ;
assign n18595 =  ( n18594 ) & (wr )  ;
assign n18596 =  ( n18595 ) ? ( n5485 ) : ( iram_136 ) ;
assign n18597 = wr_addr[7:7] ;
assign n18598 =  ( n18597 ) == ( bv_1_0_n53 )  ;
assign n18599 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n18600 =  ( n18598 ) & (n18599 )  ;
assign n18601 =  ( n18600 ) & (wr )  ;
assign n18602 =  ( n18601 ) ? ( n5512 ) : ( iram_136 ) ;
assign n18603 = wr_addr[7:7] ;
assign n18604 =  ( n18603 ) == ( bv_1_0_n53 )  ;
assign n18605 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n18606 =  ( n18604 ) & (n18605 )  ;
assign n18607 =  ( n18606 ) & (wr )  ;
assign n18608 =  ( n18607 ) ? ( bv_8_0_n69 ) : ( iram_136 ) ;
assign n18609 = wr_addr[7:7] ;
assign n18610 =  ( n18609 ) == ( bv_1_0_n53 )  ;
assign n18611 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n18612 =  ( n18610 ) & (n18611 )  ;
assign n18613 =  ( n18612 ) & (wr )  ;
assign n18614 =  ( n18613 ) ? ( n5071 ) : ( iram_136 ) ;
assign n18615 = wr_addr[7:7] ;
assign n18616 =  ( n18615 ) == ( bv_1_0_n53 )  ;
assign n18617 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n18618 =  ( n18616 ) & (n18617 )  ;
assign n18619 =  ( n18618 ) & (wr )  ;
assign n18620 =  ( n18619 ) ? ( n5096 ) : ( iram_136 ) ;
assign n18621 = wr_addr[7:7] ;
assign n18622 =  ( n18621 ) == ( bv_1_0_n53 )  ;
assign n18623 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n18624 =  ( n18622 ) & (n18623 )  ;
assign n18625 =  ( n18624 ) & (wr )  ;
assign n18626 =  ( n18625 ) ? ( n5123 ) : ( iram_136 ) ;
assign n18627 = wr_addr[7:7] ;
assign n18628 =  ( n18627 ) == ( bv_1_0_n53 )  ;
assign n18629 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n18630 =  ( n18628 ) & (n18629 )  ;
assign n18631 =  ( n18630 ) & (wr )  ;
assign n18632 =  ( n18631 ) ? ( n5165 ) : ( iram_136 ) ;
assign n18633 = wr_addr[7:7] ;
assign n18634 =  ( n18633 ) == ( bv_1_0_n53 )  ;
assign n18635 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n18636 =  ( n18634 ) & (n18635 )  ;
assign n18637 =  ( n18636 ) & (wr )  ;
assign n18638 =  ( n18637 ) ? ( n5204 ) : ( iram_136 ) ;
assign n18639 = wr_addr[7:7] ;
assign n18640 =  ( n18639 ) == ( bv_1_0_n53 )  ;
assign n18641 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n18642 =  ( n18640 ) & (n18641 )  ;
assign n18643 =  ( n18642 ) & (wr )  ;
assign n18644 =  ( n18643 ) ? ( n5262 ) : ( iram_136 ) ;
assign n18645 = wr_addr[7:7] ;
assign n18646 =  ( n18645 ) == ( bv_1_0_n53 )  ;
assign n18647 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n18648 =  ( n18646 ) & (n18647 )  ;
assign n18649 =  ( n18648 ) & (wr )  ;
assign n18650 =  ( n18649 ) ? ( n5298 ) : ( iram_136 ) ;
assign n18651 = wr_addr[7:7] ;
assign n18652 =  ( n18651 ) == ( bv_1_0_n53 )  ;
assign n18653 =  ( wr_addr ) == ( bv_8_136_n341 )  ;
assign n18654 =  ( n18652 ) & (n18653 )  ;
assign n18655 =  ( n18654 ) & (wr )  ;
assign n18656 =  ( n18655 ) ? ( n5325 ) : ( iram_136 ) ;
assign n18657 = wr_addr[7:7] ;
assign n18658 =  ( n18657 ) == ( bv_1_0_n53 )  ;
assign n18659 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n18660 =  ( n18658 ) & (n18659 )  ;
assign n18661 =  ( n18660 ) & (wr )  ;
assign n18662 =  ( n18661 ) ? ( n4782 ) : ( iram_137 ) ;
assign n18663 = wr_addr[7:7] ;
assign n18664 =  ( n18663 ) == ( bv_1_0_n53 )  ;
assign n18665 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n18666 =  ( n18664 ) & (n18665 )  ;
assign n18667 =  ( n18666 ) & (wr )  ;
assign n18668 =  ( n18667 ) ? ( n4841 ) : ( iram_137 ) ;
assign n18669 = wr_addr[7:7] ;
assign n18670 =  ( n18669 ) == ( bv_1_0_n53 )  ;
assign n18671 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n18672 =  ( n18670 ) & (n18671 )  ;
assign n18673 =  ( n18672 ) & (wr )  ;
assign n18674 =  ( n18673 ) ? ( n5449 ) : ( iram_137 ) ;
assign n18675 = wr_addr[7:7] ;
assign n18676 =  ( n18675 ) == ( bv_1_0_n53 )  ;
assign n18677 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n18678 =  ( n18676 ) & (n18677 )  ;
assign n18679 =  ( n18678 ) & (wr )  ;
assign n18680 =  ( n18679 ) ? ( n4906 ) : ( iram_137 ) ;
assign n18681 = wr_addr[7:7] ;
assign n18682 =  ( n18681 ) == ( bv_1_0_n53 )  ;
assign n18683 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n18684 =  ( n18682 ) & (n18683 )  ;
assign n18685 =  ( n18684 ) & (wr )  ;
assign n18686 =  ( n18685 ) ? ( n5485 ) : ( iram_137 ) ;
assign n18687 = wr_addr[7:7] ;
assign n18688 =  ( n18687 ) == ( bv_1_0_n53 )  ;
assign n18689 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n18690 =  ( n18688 ) & (n18689 )  ;
assign n18691 =  ( n18690 ) & (wr )  ;
assign n18692 =  ( n18691 ) ? ( n5512 ) : ( iram_137 ) ;
assign n18693 = wr_addr[7:7] ;
assign n18694 =  ( n18693 ) == ( bv_1_0_n53 )  ;
assign n18695 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n18696 =  ( n18694 ) & (n18695 )  ;
assign n18697 =  ( n18696 ) & (wr )  ;
assign n18698 =  ( n18697 ) ? ( bv_8_0_n69 ) : ( iram_137 ) ;
assign n18699 = wr_addr[7:7] ;
assign n18700 =  ( n18699 ) == ( bv_1_0_n53 )  ;
assign n18701 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n18702 =  ( n18700 ) & (n18701 )  ;
assign n18703 =  ( n18702 ) & (wr )  ;
assign n18704 =  ( n18703 ) ? ( n5071 ) : ( iram_137 ) ;
assign n18705 = wr_addr[7:7] ;
assign n18706 =  ( n18705 ) == ( bv_1_0_n53 )  ;
assign n18707 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n18708 =  ( n18706 ) & (n18707 )  ;
assign n18709 =  ( n18708 ) & (wr )  ;
assign n18710 =  ( n18709 ) ? ( n5096 ) : ( iram_137 ) ;
assign n18711 = wr_addr[7:7] ;
assign n18712 =  ( n18711 ) == ( bv_1_0_n53 )  ;
assign n18713 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n18714 =  ( n18712 ) & (n18713 )  ;
assign n18715 =  ( n18714 ) & (wr )  ;
assign n18716 =  ( n18715 ) ? ( n5123 ) : ( iram_137 ) ;
assign n18717 = wr_addr[7:7] ;
assign n18718 =  ( n18717 ) == ( bv_1_0_n53 )  ;
assign n18719 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n18720 =  ( n18718 ) & (n18719 )  ;
assign n18721 =  ( n18720 ) & (wr )  ;
assign n18722 =  ( n18721 ) ? ( n5165 ) : ( iram_137 ) ;
assign n18723 = wr_addr[7:7] ;
assign n18724 =  ( n18723 ) == ( bv_1_0_n53 )  ;
assign n18725 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n18726 =  ( n18724 ) & (n18725 )  ;
assign n18727 =  ( n18726 ) & (wr )  ;
assign n18728 =  ( n18727 ) ? ( n5204 ) : ( iram_137 ) ;
assign n18729 = wr_addr[7:7] ;
assign n18730 =  ( n18729 ) == ( bv_1_0_n53 )  ;
assign n18731 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n18732 =  ( n18730 ) & (n18731 )  ;
assign n18733 =  ( n18732 ) & (wr )  ;
assign n18734 =  ( n18733 ) ? ( n5262 ) : ( iram_137 ) ;
assign n18735 = wr_addr[7:7] ;
assign n18736 =  ( n18735 ) == ( bv_1_0_n53 )  ;
assign n18737 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n18738 =  ( n18736 ) & (n18737 )  ;
assign n18739 =  ( n18738 ) & (wr )  ;
assign n18740 =  ( n18739 ) ? ( n5298 ) : ( iram_137 ) ;
assign n18741 = wr_addr[7:7] ;
assign n18742 =  ( n18741 ) == ( bv_1_0_n53 )  ;
assign n18743 =  ( wr_addr ) == ( bv_8_137_n343 )  ;
assign n18744 =  ( n18742 ) & (n18743 )  ;
assign n18745 =  ( n18744 ) & (wr )  ;
assign n18746 =  ( n18745 ) ? ( n5325 ) : ( iram_137 ) ;
assign n18747 = wr_addr[7:7] ;
assign n18748 =  ( n18747 ) == ( bv_1_0_n53 )  ;
assign n18749 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n18750 =  ( n18748 ) & (n18749 )  ;
assign n18751 =  ( n18750 ) & (wr )  ;
assign n18752 =  ( n18751 ) ? ( n4782 ) : ( iram_138 ) ;
assign n18753 = wr_addr[7:7] ;
assign n18754 =  ( n18753 ) == ( bv_1_0_n53 )  ;
assign n18755 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n18756 =  ( n18754 ) & (n18755 )  ;
assign n18757 =  ( n18756 ) & (wr )  ;
assign n18758 =  ( n18757 ) ? ( n4841 ) : ( iram_138 ) ;
assign n18759 = wr_addr[7:7] ;
assign n18760 =  ( n18759 ) == ( bv_1_0_n53 )  ;
assign n18761 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n18762 =  ( n18760 ) & (n18761 )  ;
assign n18763 =  ( n18762 ) & (wr )  ;
assign n18764 =  ( n18763 ) ? ( n5449 ) : ( iram_138 ) ;
assign n18765 = wr_addr[7:7] ;
assign n18766 =  ( n18765 ) == ( bv_1_0_n53 )  ;
assign n18767 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n18768 =  ( n18766 ) & (n18767 )  ;
assign n18769 =  ( n18768 ) & (wr )  ;
assign n18770 =  ( n18769 ) ? ( n4906 ) : ( iram_138 ) ;
assign n18771 = wr_addr[7:7] ;
assign n18772 =  ( n18771 ) == ( bv_1_0_n53 )  ;
assign n18773 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n18774 =  ( n18772 ) & (n18773 )  ;
assign n18775 =  ( n18774 ) & (wr )  ;
assign n18776 =  ( n18775 ) ? ( n5485 ) : ( iram_138 ) ;
assign n18777 = wr_addr[7:7] ;
assign n18778 =  ( n18777 ) == ( bv_1_0_n53 )  ;
assign n18779 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n18780 =  ( n18778 ) & (n18779 )  ;
assign n18781 =  ( n18780 ) & (wr )  ;
assign n18782 =  ( n18781 ) ? ( n5512 ) : ( iram_138 ) ;
assign n18783 = wr_addr[7:7] ;
assign n18784 =  ( n18783 ) == ( bv_1_0_n53 )  ;
assign n18785 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n18786 =  ( n18784 ) & (n18785 )  ;
assign n18787 =  ( n18786 ) & (wr )  ;
assign n18788 =  ( n18787 ) ? ( bv_8_0_n69 ) : ( iram_138 ) ;
assign n18789 = wr_addr[7:7] ;
assign n18790 =  ( n18789 ) == ( bv_1_0_n53 )  ;
assign n18791 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n18792 =  ( n18790 ) & (n18791 )  ;
assign n18793 =  ( n18792 ) & (wr )  ;
assign n18794 =  ( n18793 ) ? ( n5071 ) : ( iram_138 ) ;
assign n18795 = wr_addr[7:7] ;
assign n18796 =  ( n18795 ) == ( bv_1_0_n53 )  ;
assign n18797 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n18798 =  ( n18796 ) & (n18797 )  ;
assign n18799 =  ( n18798 ) & (wr )  ;
assign n18800 =  ( n18799 ) ? ( n5096 ) : ( iram_138 ) ;
assign n18801 = wr_addr[7:7] ;
assign n18802 =  ( n18801 ) == ( bv_1_0_n53 )  ;
assign n18803 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n18804 =  ( n18802 ) & (n18803 )  ;
assign n18805 =  ( n18804 ) & (wr )  ;
assign n18806 =  ( n18805 ) ? ( n5123 ) : ( iram_138 ) ;
assign n18807 = wr_addr[7:7] ;
assign n18808 =  ( n18807 ) == ( bv_1_0_n53 )  ;
assign n18809 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n18810 =  ( n18808 ) & (n18809 )  ;
assign n18811 =  ( n18810 ) & (wr )  ;
assign n18812 =  ( n18811 ) ? ( n5165 ) : ( iram_138 ) ;
assign n18813 = wr_addr[7:7] ;
assign n18814 =  ( n18813 ) == ( bv_1_0_n53 )  ;
assign n18815 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n18816 =  ( n18814 ) & (n18815 )  ;
assign n18817 =  ( n18816 ) & (wr )  ;
assign n18818 =  ( n18817 ) ? ( n5204 ) : ( iram_138 ) ;
assign n18819 = wr_addr[7:7] ;
assign n18820 =  ( n18819 ) == ( bv_1_0_n53 )  ;
assign n18821 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n18822 =  ( n18820 ) & (n18821 )  ;
assign n18823 =  ( n18822 ) & (wr )  ;
assign n18824 =  ( n18823 ) ? ( n5262 ) : ( iram_138 ) ;
assign n18825 = wr_addr[7:7] ;
assign n18826 =  ( n18825 ) == ( bv_1_0_n53 )  ;
assign n18827 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n18828 =  ( n18826 ) & (n18827 )  ;
assign n18829 =  ( n18828 ) & (wr )  ;
assign n18830 =  ( n18829 ) ? ( n5298 ) : ( iram_138 ) ;
assign n18831 = wr_addr[7:7] ;
assign n18832 =  ( n18831 ) == ( bv_1_0_n53 )  ;
assign n18833 =  ( wr_addr ) == ( bv_8_138_n345 )  ;
assign n18834 =  ( n18832 ) & (n18833 )  ;
assign n18835 =  ( n18834 ) & (wr )  ;
assign n18836 =  ( n18835 ) ? ( n5325 ) : ( iram_138 ) ;
assign n18837 = wr_addr[7:7] ;
assign n18838 =  ( n18837 ) == ( bv_1_0_n53 )  ;
assign n18839 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n18840 =  ( n18838 ) & (n18839 )  ;
assign n18841 =  ( n18840 ) & (wr )  ;
assign n18842 =  ( n18841 ) ? ( n4782 ) : ( iram_139 ) ;
assign n18843 = wr_addr[7:7] ;
assign n18844 =  ( n18843 ) == ( bv_1_0_n53 )  ;
assign n18845 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n18846 =  ( n18844 ) & (n18845 )  ;
assign n18847 =  ( n18846 ) & (wr )  ;
assign n18848 =  ( n18847 ) ? ( n4841 ) : ( iram_139 ) ;
assign n18849 = wr_addr[7:7] ;
assign n18850 =  ( n18849 ) == ( bv_1_0_n53 )  ;
assign n18851 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n18852 =  ( n18850 ) & (n18851 )  ;
assign n18853 =  ( n18852 ) & (wr )  ;
assign n18854 =  ( n18853 ) ? ( n5449 ) : ( iram_139 ) ;
assign n18855 = wr_addr[7:7] ;
assign n18856 =  ( n18855 ) == ( bv_1_0_n53 )  ;
assign n18857 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n18858 =  ( n18856 ) & (n18857 )  ;
assign n18859 =  ( n18858 ) & (wr )  ;
assign n18860 =  ( n18859 ) ? ( n4906 ) : ( iram_139 ) ;
assign n18861 = wr_addr[7:7] ;
assign n18862 =  ( n18861 ) == ( bv_1_0_n53 )  ;
assign n18863 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n18864 =  ( n18862 ) & (n18863 )  ;
assign n18865 =  ( n18864 ) & (wr )  ;
assign n18866 =  ( n18865 ) ? ( n5485 ) : ( iram_139 ) ;
assign n18867 = wr_addr[7:7] ;
assign n18868 =  ( n18867 ) == ( bv_1_0_n53 )  ;
assign n18869 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n18870 =  ( n18868 ) & (n18869 )  ;
assign n18871 =  ( n18870 ) & (wr )  ;
assign n18872 =  ( n18871 ) ? ( n5512 ) : ( iram_139 ) ;
assign n18873 = wr_addr[7:7] ;
assign n18874 =  ( n18873 ) == ( bv_1_0_n53 )  ;
assign n18875 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n18876 =  ( n18874 ) & (n18875 )  ;
assign n18877 =  ( n18876 ) & (wr )  ;
assign n18878 =  ( n18877 ) ? ( bv_8_0_n69 ) : ( iram_139 ) ;
assign n18879 = wr_addr[7:7] ;
assign n18880 =  ( n18879 ) == ( bv_1_0_n53 )  ;
assign n18881 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n18882 =  ( n18880 ) & (n18881 )  ;
assign n18883 =  ( n18882 ) & (wr )  ;
assign n18884 =  ( n18883 ) ? ( n5071 ) : ( iram_139 ) ;
assign n18885 = wr_addr[7:7] ;
assign n18886 =  ( n18885 ) == ( bv_1_0_n53 )  ;
assign n18887 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n18888 =  ( n18886 ) & (n18887 )  ;
assign n18889 =  ( n18888 ) & (wr )  ;
assign n18890 =  ( n18889 ) ? ( n5096 ) : ( iram_139 ) ;
assign n18891 = wr_addr[7:7] ;
assign n18892 =  ( n18891 ) == ( bv_1_0_n53 )  ;
assign n18893 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n18894 =  ( n18892 ) & (n18893 )  ;
assign n18895 =  ( n18894 ) & (wr )  ;
assign n18896 =  ( n18895 ) ? ( n5123 ) : ( iram_139 ) ;
assign n18897 = wr_addr[7:7] ;
assign n18898 =  ( n18897 ) == ( bv_1_0_n53 )  ;
assign n18899 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n18900 =  ( n18898 ) & (n18899 )  ;
assign n18901 =  ( n18900 ) & (wr )  ;
assign n18902 =  ( n18901 ) ? ( n5165 ) : ( iram_139 ) ;
assign n18903 = wr_addr[7:7] ;
assign n18904 =  ( n18903 ) == ( bv_1_0_n53 )  ;
assign n18905 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n18906 =  ( n18904 ) & (n18905 )  ;
assign n18907 =  ( n18906 ) & (wr )  ;
assign n18908 =  ( n18907 ) ? ( n5204 ) : ( iram_139 ) ;
assign n18909 = wr_addr[7:7] ;
assign n18910 =  ( n18909 ) == ( bv_1_0_n53 )  ;
assign n18911 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n18912 =  ( n18910 ) & (n18911 )  ;
assign n18913 =  ( n18912 ) & (wr )  ;
assign n18914 =  ( n18913 ) ? ( n5262 ) : ( iram_139 ) ;
assign n18915 = wr_addr[7:7] ;
assign n18916 =  ( n18915 ) == ( bv_1_0_n53 )  ;
assign n18917 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n18918 =  ( n18916 ) & (n18917 )  ;
assign n18919 =  ( n18918 ) & (wr )  ;
assign n18920 =  ( n18919 ) ? ( n5298 ) : ( iram_139 ) ;
assign n18921 = wr_addr[7:7] ;
assign n18922 =  ( n18921 ) == ( bv_1_0_n53 )  ;
assign n18923 =  ( wr_addr ) == ( bv_8_139_n347 )  ;
assign n18924 =  ( n18922 ) & (n18923 )  ;
assign n18925 =  ( n18924 ) & (wr )  ;
assign n18926 =  ( n18925 ) ? ( n5325 ) : ( iram_139 ) ;
assign n18927 = wr_addr[7:7] ;
assign n18928 =  ( n18927 ) == ( bv_1_0_n53 )  ;
assign n18929 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n18930 =  ( n18928 ) & (n18929 )  ;
assign n18931 =  ( n18930 ) & (wr )  ;
assign n18932 =  ( n18931 ) ? ( n4782 ) : ( iram_140 ) ;
assign n18933 = wr_addr[7:7] ;
assign n18934 =  ( n18933 ) == ( bv_1_0_n53 )  ;
assign n18935 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n18936 =  ( n18934 ) & (n18935 )  ;
assign n18937 =  ( n18936 ) & (wr )  ;
assign n18938 =  ( n18937 ) ? ( n4841 ) : ( iram_140 ) ;
assign n18939 = wr_addr[7:7] ;
assign n18940 =  ( n18939 ) == ( bv_1_0_n53 )  ;
assign n18941 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n18942 =  ( n18940 ) & (n18941 )  ;
assign n18943 =  ( n18942 ) & (wr )  ;
assign n18944 =  ( n18943 ) ? ( n5449 ) : ( iram_140 ) ;
assign n18945 = wr_addr[7:7] ;
assign n18946 =  ( n18945 ) == ( bv_1_0_n53 )  ;
assign n18947 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n18948 =  ( n18946 ) & (n18947 )  ;
assign n18949 =  ( n18948 ) & (wr )  ;
assign n18950 =  ( n18949 ) ? ( n4906 ) : ( iram_140 ) ;
assign n18951 = wr_addr[7:7] ;
assign n18952 =  ( n18951 ) == ( bv_1_0_n53 )  ;
assign n18953 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n18954 =  ( n18952 ) & (n18953 )  ;
assign n18955 =  ( n18954 ) & (wr )  ;
assign n18956 =  ( n18955 ) ? ( n5485 ) : ( iram_140 ) ;
assign n18957 = wr_addr[7:7] ;
assign n18958 =  ( n18957 ) == ( bv_1_0_n53 )  ;
assign n18959 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n18960 =  ( n18958 ) & (n18959 )  ;
assign n18961 =  ( n18960 ) & (wr )  ;
assign n18962 =  ( n18961 ) ? ( n5512 ) : ( iram_140 ) ;
assign n18963 = wr_addr[7:7] ;
assign n18964 =  ( n18963 ) == ( bv_1_0_n53 )  ;
assign n18965 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n18966 =  ( n18964 ) & (n18965 )  ;
assign n18967 =  ( n18966 ) & (wr )  ;
assign n18968 =  ( n18967 ) ? ( bv_8_0_n69 ) : ( iram_140 ) ;
assign n18969 = wr_addr[7:7] ;
assign n18970 =  ( n18969 ) == ( bv_1_0_n53 )  ;
assign n18971 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n18972 =  ( n18970 ) & (n18971 )  ;
assign n18973 =  ( n18972 ) & (wr )  ;
assign n18974 =  ( n18973 ) ? ( n5071 ) : ( iram_140 ) ;
assign n18975 = wr_addr[7:7] ;
assign n18976 =  ( n18975 ) == ( bv_1_0_n53 )  ;
assign n18977 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n18978 =  ( n18976 ) & (n18977 )  ;
assign n18979 =  ( n18978 ) & (wr )  ;
assign n18980 =  ( n18979 ) ? ( n5096 ) : ( iram_140 ) ;
assign n18981 = wr_addr[7:7] ;
assign n18982 =  ( n18981 ) == ( bv_1_0_n53 )  ;
assign n18983 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n18984 =  ( n18982 ) & (n18983 )  ;
assign n18985 =  ( n18984 ) & (wr )  ;
assign n18986 =  ( n18985 ) ? ( n5123 ) : ( iram_140 ) ;
assign n18987 = wr_addr[7:7] ;
assign n18988 =  ( n18987 ) == ( bv_1_0_n53 )  ;
assign n18989 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n18990 =  ( n18988 ) & (n18989 )  ;
assign n18991 =  ( n18990 ) & (wr )  ;
assign n18992 =  ( n18991 ) ? ( n5165 ) : ( iram_140 ) ;
assign n18993 = wr_addr[7:7] ;
assign n18994 =  ( n18993 ) == ( bv_1_0_n53 )  ;
assign n18995 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n18996 =  ( n18994 ) & (n18995 )  ;
assign n18997 =  ( n18996 ) & (wr )  ;
assign n18998 =  ( n18997 ) ? ( n5204 ) : ( iram_140 ) ;
assign n18999 = wr_addr[7:7] ;
assign n19000 =  ( n18999 ) == ( bv_1_0_n53 )  ;
assign n19001 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n19002 =  ( n19000 ) & (n19001 )  ;
assign n19003 =  ( n19002 ) & (wr )  ;
assign n19004 =  ( n19003 ) ? ( n5262 ) : ( iram_140 ) ;
assign n19005 = wr_addr[7:7] ;
assign n19006 =  ( n19005 ) == ( bv_1_0_n53 )  ;
assign n19007 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n19008 =  ( n19006 ) & (n19007 )  ;
assign n19009 =  ( n19008 ) & (wr )  ;
assign n19010 =  ( n19009 ) ? ( n5298 ) : ( iram_140 ) ;
assign n19011 = wr_addr[7:7] ;
assign n19012 =  ( n19011 ) == ( bv_1_0_n53 )  ;
assign n19013 =  ( wr_addr ) == ( bv_8_140_n349 )  ;
assign n19014 =  ( n19012 ) & (n19013 )  ;
assign n19015 =  ( n19014 ) & (wr )  ;
assign n19016 =  ( n19015 ) ? ( n5325 ) : ( iram_140 ) ;
assign n19017 = wr_addr[7:7] ;
assign n19018 =  ( n19017 ) == ( bv_1_0_n53 )  ;
assign n19019 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n19020 =  ( n19018 ) & (n19019 )  ;
assign n19021 =  ( n19020 ) & (wr )  ;
assign n19022 =  ( n19021 ) ? ( n4782 ) : ( iram_141 ) ;
assign n19023 = wr_addr[7:7] ;
assign n19024 =  ( n19023 ) == ( bv_1_0_n53 )  ;
assign n19025 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n19026 =  ( n19024 ) & (n19025 )  ;
assign n19027 =  ( n19026 ) & (wr )  ;
assign n19028 =  ( n19027 ) ? ( n4841 ) : ( iram_141 ) ;
assign n19029 = wr_addr[7:7] ;
assign n19030 =  ( n19029 ) == ( bv_1_0_n53 )  ;
assign n19031 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n19032 =  ( n19030 ) & (n19031 )  ;
assign n19033 =  ( n19032 ) & (wr )  ;
assign n19034 =  ( n19033 ) ? ( n5449 ) : ( iram_141 ) ;
assign n19035 = wr_addr[7:7] ;
assign n19036 =  ( n19035 ) == ( bv_1_0_n53 )  ;
assign n19037 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n19038 =  ( n19036 ) & (n19037 )  ;
assign n19039 =  ( n19038 ) & (wr )  ;
assign n19040 =  ( n19039 ) ? ( n4906 ) : ( iram_141 ) ;
assign n19041 = wr_addr[7:7] ;
assign n19042 =  ( n19041 ) == ( bv_1_0_n53 )  ;
assign n19043 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n19044 =  ( n19042 ) & (n19043 )  ;
assign n19045 =  ( n19044 ) & (wr )  ;
assign n19046 =  ( n19045 ) ? ( n5485 ) : ( iram_141 ) ;
assign n19047 = wr_addr[7:7] ;
assign n19048 =  ( n19047 ) == ( bv_1_0_n53 )  ;
assign n19049 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n19050 =  ( n19048 ) & (n19049 )  ;
assign n19051 =  ( n19050 ) & (wr )  ;
assign n19052 =  ( n19051 ) ? ( n5512 ) : ( iram_141 ) ;
assign n19053 = wr_addr[7:7] ;
assign n19054 =  ( n19053 ) == ( bv_1_0_n53 )  ;
assign n19055 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n19056 =  ( n19054 ) & (n19055 )  ;
assign n19057 =  ( n19056 ) & (wr )  ;
assign n19058 =  ( n19057 ) ? ( bv_8_0_n69 ) : ( iram_141 ) ;
assign n19059 = wr_addr[7:7] ;
assign n19060 =  ( n19059 ) == ( bv_1_0_n53 )  ;
assign n19061 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n19062 =  ( n19060 ) & (n19061 )  ;
assign n19063 =  ( n19062 ) & (wr )  ;
assign n19064 =  ( n19063 ) ? ( n5071 ) : ( iram_141 ) ;
assign n19065 = wr_addr[7:7] ;
assign n19066 =  ( n19065 ) == ( bv_1_0_n53 )  ;
assign n19067 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n19068 =  ( n19066 ) & (n19067 )  ;
assign n19069 =  ( n19068 ) & (wr )  ;
assign n19070 =  ( n19069 ) ? ( n5096 ) : ( iram_141 ) ;
assign n19071 = wr_addr[7:7] ;
assign n19072 =  ( n19071 ) == ( bv_1_0_n53 )  ;
assign n19073 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n19074 =  ( n19072 ) & (n19073 )  ;
assign n19075 =  ( n19074 ) & (wr )  ;
assign n19076 =  ( n19075 ) ? ( n5123 ) : ( iram_141 ) ;
assign n19077 = wr_addr[7:7] ;
assign n19078 =  ( n19077 ) == ( bv_1_0_n53 )  ;
assign n19079 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n19080 =  ( n19078 ) & (n19079 )  ;
assign n19081 =  ( n19080 ) & (wr )  ;
assign n19082 =  ( n19081 ) ? ( n5165 ) : ( iram_141 ) ;
assign n19083 = wr_addr[7:7] ;
assign n19084 =  ( n19083 ) == ( bv_1_0_n53 )  ;
assign n19085 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n19086 =  ( n19084 ) & (n19085 )  ;
assign n19087 =  ( n19086 ) & (wr )  ;
assign n19088 =  ( n19087 ) ? ( n5204 ) : ( iram_141 ) ;
assign n19089 = wr_addr[7:7] ;
assign n19090 =  ( n19089 ) == ( bv_1_0_n53 )  ;
assign n19091 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n19092 =  ( n19090 ) & (n19091 )  ;
assign n19093 =  ( n19092 ) & (wr )  ;
assign n19094 =  ( n19093 ) ? ( n5262 ) : ( iram_141 ) ;
assign n19095 = wr_addr[7:7] ;
assign n19096 =  ( n19095 ) == ( bv_1_0_n53 )  ;
assign n19097 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n19098 =  ( n19096 ) & (n19097 )  ;
assign n19099 =  ( n19098 ) & (wr )  ;
assign n19100 =  ( n19099 ) ? ( n5298 ) : ( iram_141 ) ;
assign n19101 = wr_addr[7:7] ;
assign n19102 =  ( n19101 ) == ( bv_1_0_n53 )  ;
assign n19103 =  ( wr_addr ) == ( bv_8_141_n351 )  ;
assign n19104 =  ( n19102 ) & (n19103 )  ;
assign n19105 =  ( n19104 ) & (wr )  ;
assign n19106 =  ( n19105 ) ? ( n5325 ) : ( iram_141 ) ;
assign n19107 = wr_addr[7:7] ;
assign n19108 =  ( n19107 ) == ( bv_1_0_n53 )  ;
assign n19109 =  ( wr_addr ) == ( bv_8_142_n353 )  ;
assign n19110 =  ( n19108 ) & (n19109 )  ;
assign n19111 =  ( n19110 ) & (wr )  ;
assign n19112 =  ( n19111 ) ? ( n4782 ) : ( iram_142 ) ;
assign n19113 = wr_addr[7:7] ;
assign n19114 =  ( n19113 ) == ( bv_1_0_n53 )  ;
assign n19115 =  ( wr_addr ) == ( bv_8_142_n353 )  ;
assign n19116 =  ( n19114 ) & (n19115 )  ;
assign n19117 =  ( n19116 ) & (wr )  ;
assign n19118 =  ( n19117 ) ? ( n4841 ) : ( iram_142 ) ;
assign n19119 = wr_addr[7:7] ;
assign n19120 =  ( n19119 ) == ( bv_1_0_n53 )  ;
assign n19121 =  ( wr_addr ) == ( bv_8_142_n353 )  ;
assign n19122 =  ( n19120 ) & (n19121 )  ;
assign n19123 =  ( n19122 ) & (wr )  ;
assign n19124 =  ( n19123 ) ? ( n5449 ) : ( iram_142 ) ;
assign n19125 = wr_addr[7:7] ;
assign n19126 =  ( n19125 ) == ( bv_1_0_n53 )  ;
assign n19127 =  ( wr_addr ) == ( bv_8_142_n353 )  ;
assign n19128 =  ( n19126 ) & (n19127 )  ;
assign n19129 =  ( n19128 ) & (wr )  ;
assign n19130 =  ( n19129 ) ? ( n4906 ) : ( iram_142 ) ;
assign n19131 = wr_addr[7:7] ;
assign n19132 =  ( n19131 ) == ( bv_1_0_n53 )  ;
assign n19133 =  ( wr_addr ) == ( bv_8_142_n353 )  ;
assign n19134 =  ( n19132 ) & (n19133 )  ;
assign n19135 =  ( n19134 ) & (wr )  ;
assign n19136 =  ( n19135 ) ? ( n5485 ) : ( iram_142 ) ;
assign n19137 = wr_addr[7:7] ;
assign n19138 =  ( n19137 ) == ( bv_1_0_n53 )  ;
assign n19139 =  ( wr_addr ) == ( bv_8_142_n353 )  ;
assign n19140 =  ( n19138 ) & (n19139 )  ;
assign n19141 =  ( n19140 ) & (wr )  ;
assign n19142 =  ( n19141 ) ? ( n5512 ) : ( iram_142 ) ;
assign n19143 = wr_addr[7:7] ;
assign n19144 =  ( n19143 ) == ( bv_1_0_n53 )  ;
assign n19145 =  ( wr_addr ) == ( bv_8_142_n353 )  ;
assign n19146 =  ( n19144 ) & (n19145 )  ;
assign n19147 =  ( n19146 ) & (wr )  ;
assign n19148 =  ( n19147 ) ? ( bv_8_0_n69 ) : ( iram_142 ) ;
assign n19149 = wr_addr[7:7] ;
assign n19150 =  ( n19149 ) == ( bv_1_0_n53 )  ;
assign n19151 =  ( wr_addr ) == ( bv_8_142_n353 )  ;
assign n19152 =  ( n19150 ) & (n19151 )  ;
assign n19153 =  ( n19152 ) & (wr )  ;
assign n19154 =  ( n19153 ) ? ( n5071 ) : ( iram_142 ) ;
assign n19155 = wr_addr[7:7] ;
assign n19156 =  ( n19155 ) == ( bv_1_0_n53 )  ;
assign n19157 =  ( wr_addr ) == ( bv_8_142_n353 )  ;
assign n19158 =  ( n19156 ) & (n19157 )  ;
assign n19159 =  ( n19158 ) & (wr )  ;
assign n19160 =  ( n19159 ) ? ( n5096 ) : ( iram_142 ) ;
assign n19161 = wr_addr[7:7] ;
assign n19162 =  ( n19161 ) == ( bv_1_0_n53 )  ;
assign n19163 =  ( wr_addr ) == ( bv_8_142_n353 )  ;
assign n19164 =  ( n19162 ) & (n19163 )  ;
assign n19165 =  ( n19164 ) & (wr )  ;
assign n19166 =  ( n19165 ) ? ( n5123 ) : ( iram_142 ) ;
assign n19167 = wr_addr[7:7] ;
assign n19168 =  ( n19167 ) == ( bv_1_0_n53 )  ;
assign n19169 =  ( wr_addr ) == ( bv_8_142_n353 )  ;
assign n19170 =  ( n19168 ) & (n19169 )  ;
assign n19171 =  ( n19170 ) & (wr )  ;
assign n19172 =  ( n19171 ) ? ( n5165 ) : ( iram_142 ) ;
assign n19173 = wr_addr[7:7] ;
assign n19174 =  ( n19173 ) == ( bv_1_0_n53 )  ;
assign n19175 =  ( wr_addr ) == ( bv_8_142_n353 )  ;
assign n19176 =  ( n19174 ) & (n19175 )  ;
assign n19177 =  ( n19176 ) & (wr )  ;
assign n19178 =  ( n19177 ) ? ( n5204 ) : ( iram_142 ) ;
assign n19179 = wr_addr[7:7] ;
assign n19180 =  ( n19179 ) == ( bv_1_0_n53 )  ;
assign n19181 =  ( wr_addr ) == ( bv_8_142_n353 )  ;
assign n19182 =  ( n19180 ) & (n19181 )  ;
assign n19183 =  ( n19182 ) & (wr )  ;
assign n19184 =  ( n19183 ) ? ( n5262 ) : ( iram_142 ) ;
assign n19185 = wr_addr[7:7] ;
assign n19186 =  ( n19185 ) == ( bv_1_0_n53 )  ;
assign n19187 =  ( wr_addr ) == ( bv_8_142_n353 )  ;
assign n19188 =  ( n19186 ) & (n19187 )  ;
assign n19189 =  ( n19188 ) & (wr )  ;
assign n19190 =  ( n19189 ) ? ( n5298 ) : ( iram_142 ) ;
assign n19191 = wr_addr[7:7] ;
assign n19192 =  ( n19191 ) == ( bv_1_0_n53 )  ;
assign n19193 =  ( wr_addr ) == ( bv_8_142_n353 )  ;
assign n19194 =  ( n19192 ) & (n19193 )  ;
assign n19195 =  ( n19194 ) & (wr )  ;
assign n19196 =  ( n19195 ) ? ( n5325 ) : ( iram_142 ) ;
assign n19197 = wr_addr[7:7] ;
assign n19198 =  ( n19197 ) == ( bv_1_0_n53 )  ;
assign n19199 =  ( wr_addr ) == ( bv_8_143_n355 )  ;
assign n19200 =  ( n19198 ) & (n19199 )  ;
assign n19201 =  ( n19200 ) & (wr )  ;
assign n19202 =  ( n19201 ) ? ( n4782 ) : ( iram_143 ) ;
assign n19203 = wr_addr[7:7] ;
assign n19204 =  ( n19203 ) == ( bv_1_0_n53 )  ;
assign n19205 =  ( wr_addr ) == ( bv_8_143_n355 )  ;
assign n19206 =  ( n19204 ) & (n19205 )  ;
assign n19207 =  ( n19206 ) & (wr )  ;
assign n19208 =  ( n19207 ) ? ( n4841 ) : ( iram_143 ) ;
assign n19209 = wr_addr[7:7] ;
assign n19210 =  ( n19209 ) == ( bv_1_0_n53 )  ;
assign n19211 =  ( wr_addr ) == ( bv_8_143_n355 )  ;
assign n19212 =  ( n19210 ) & (n19211 )  ;
assign n19213 =  ( n19212 ) & (wr )  ;
assign n19214 =  ( n19213 ) ? ( n5449 ) : ( iram_143 ) ;
assign n19215 = wr_addr[7:7] ;
assign n19216 =  ( n19215 ) == ( bv_1_0_n53 )  ;
assign n19217 =  ( wr_addr ) == ( bv_8_143_n355 )  ;
assign n19218 =  ( n19216 ) & (n19217 )  ;
assign n19219 =  ( n19218 ) & (wr )  ;
assign n19220 =  ( n19219 ) ? ( n4906 ) : ( iram_143 ) ;
assign n19221 = wr_addr[7:7] ;
assign n19222 =  ( n19221 ) == ( bv_1_0_n53 )  ;
assign n19223 =  ( wr_addr ) == ( bv_8_143_n355 )  ;
assign n19224 =  ( n19222 ) & (n19223 )  ;
assign n19225 =  ( n19224 ) & (wr )  ;
assign n19226 =  ( n19225 ) ? ( n5485 ) : ( iram_143 ) ;
assign n19227 = wr_addr[7:7] ;
assign n19228 =  ( n19227 ) == ( bv_1_0_n53 )  ;
assign n19229 =  ( wr_addr ) == ( bv_8_143_n355 )  ;
assign n19230 =  ( n19228 ) & (n19229 )  ;
assign n19231 =  ( n19230 ) & (wr )  ;
assign n19232 =  ( n19231 ) ? ( n5512 ) : ( iram_143 ) ;
assign n19233 = wr_addr[7:7] ;
assign n19234 =  ( n19233 ) == ( bv_1_0_n53 )  ;
assign n19235 =  ( wr_addr ) == ( bv_8_143_n355 )  ;
assign n19236 =  ( n19234 ) & (n19235 )  ;
assign n19237 =  ( n19236 ) & (wr )  ;
assign n19238 =  ( n19237 ) ? ( bv_8_0_n69 ) : ( iram_143 ) ;
assign n19239 = wr_addr[7:7] ;
assign n19240 =  ( n19239 ) == ( bv_1_0_n53 )  ;
assign n19241 =  ( wr_addr ) == ( bv_8_143_n355 )  ;
assign n19242 =  ( n19240 ) & (n19241 )  ;
assign n19243 =  ( n19242 ) & (wr )  ;
assign n19244 =  ( n19243 ) ? ( n5071 ) : ( iram_143 ) ;
assign n19245 = wr_addr[7:7] ;
assign n19246 =  ( n19245 ) == ( bv_1_0_n53 )  ;
assign n19247 =  ( wr_addr ) == ( bv_8_143_n355 )  ;
assign n19248 =  ( n19246 ) & (n19247 )  ;
assign n19249 =  ( n19248 ) & (wr )  ;
assign n19250 =  ( n19249 ) ? ( n5096 ) : ( iram_143 ) ;
assign n19251 = wr_addr[7:7] ;
assign n19252 =  ( n19251 ) == ( bv_1_0_n53 )  ;
assign n19253 =  ( wr_addr ) == ( bv_8_143_n355 )  ;
assign n19254 =  ( n19252 ) & (n19253 )  ;
assign n19255 =  ( n19254 ) & (wr )  ;
assign n19256 =  ( n19255 ) ? ( n5123 ) : ( iram_143 ) ;
assign n19257 = wr_addr[7:7] ;
assign n19258 =  ( n19257 ) == ( bv_1_0_n53 )  ;
assign n19259 =  ( wr_addr ) == ( bv_8_143_n355 )  ;
assign n19260 =  ( n19258 ) & (n19259 )  ;
assign n19261 =  ( n19260 ) & (wr )  ;
assign n19262 =  ( n19261 ) ? ( n5165 ) : ( iram_143 ) ;
assign n19263 = wr_addr[7:7] ;
assign n19264 =  ( n19263 ) == ( bv_1_0_n53 )  ;
assign n19265 =  ( wr_addr ) == ( bv_8_143_n355 )  ;
assign n19266 =  ( n19264 ) & (n19265 )  ;
assign n19267 =  ( n19266 ) & (wr )  ;
assign n19268 =  ( n19267 ) ? ( n5204 ) : ( iram_143 ) ;
assign n19269 = wr_addr[7:7] ;
assign n19270 =  ( n19269 ) == ( bv_1_0_n53 )  ;
assign n19271 =  ( wr_addr ) == ( bv_8_143_n355 )  ;
assign n19272 =  ( n19270 ) & (n19271 )  ;
assign n19273 =  ( n19272 ) & (wr )  ;
assign n19274 =  ( n19273 ) ? ( n5262 ) : ( iram_143 ) ;
assign n19275 = wr_addr[7:7] ;
assign n19276 =  ( n19275 ) == ( bv_1_0_n53 )  ;
assign n19277 =  ( wr_addr ) == ( bv_8_143_n355 )  ;
assign n19278 =  ( n19276 ) & (n19277 )  ;
assign n19279 =  ( n19278 ) & (wr )  ;
assign n19280 =  ( n19279 ) ? ( n5298 ) : ( iram_143 ) ;
assign n19281 = wr_addr[7:7] ;
assign n19282 =  ( n19281 ) == ( bv_1_0_n53 )  ;
assign n19283 =  ( wr_addr ) == ( bv_8_143_n355 )  ;
assign n19284 =  ( n19282 ) & (n19283 )  ;
assign n19285 =  ( n19284 ) & (wr )  ;
assign n19286 =  ( n19285 ) ? ( n5325 ) : ( iram_143 ) ;
assign n19287 = wr_addr[7:7] ;
assign n19288 =  ( n19287 ) == ( bv_1_0_n53 )  ;
assign n19289 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n19290 =  ( n19288 ) & (n19289 )  ;
assign n19291 =  ( n19290 ) & (wr )  ;
assign n19292 =  ( n19291 ) ? ( n4782 ) : ( iram_144 ) ;
assign n19293 = wr_addr[7:7] ;
assign n19294 =  ( n19293 ) == ( bv_1_0_n53 )  ;
assign n19295 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n19296 =  ( n19294 ) & (n19295 )  ;
assign n19297 =  ( n19296 ) & (wr )  ;
assign n19298 =  ( n19297 ) ? ( n4841 ) : ( iram_144 ) ;
assign n19299 = wr_addr[7:7] ;
assign n19300 =  ( n19299 ) == ( bv_1_0_n53 )  ;
assign n19301 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n19302 =  ( n19300 ) & (n19301 )  ;
assign n19303 =  ( n19302 ) & (wr )  ;
assign n19304 =  ( n19303 ) ? ( n5449 ) : ( iram_144 ) ;
assign n19305 = wr_addr[7:7] ;
assign n19306 =  ( n19305 ) == ( bv_1_0_n53 )  ;
assign n19307 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n19308 =  ( n19306 ) & (n19307 )  ;
assign n19309 =  ( n19308 ) & (wr )  ;
assign n19310 =  ( n19309 ) ? ( n4906 ) : ( iram_144 ) ;
assign n19311 = wr_addr[7:7] ;
assign n19312 =  ( n19311 ) == ( bv_1_0_n53 )  ;
assign n19313 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n19314 =  ( n19312 ) & (n19313 )  ;
assign n19315 =  ( n19314 ) & (wr )  ;
assign n19316 =  ( n19315 ) ? ( n5485 ) : ( iram_144 ) ;
assign n19317 = wr_addr[7:7] ;
assign n19318 =  ( n19317 ) == ( bv_1_0_n53 )  ;
assign n19319 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n19320 =  ( n19318 ) & (n19319 )  ;
assign n19321 =  ( n19320 ) & (wr )  ;
assign n19322 =  ( n19321 ) ? ( n5512 ) : ( iram_144 ) ;
assign n19323 = wr_addr[7:7] ;
assign n19324 =  ( n19323 ) == ( bv_1_0_n53 )  ;
assign n19325 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n19326 =  ( n19324 ) & (n19325 )  ;
assign n19327 =  ( n19326 ) & (wr )  ;
assign n19328 =  ( n19327 ) ? ( bv_8_0_n69 ) : ( iram_144 ) ;
assign n19329 = wr_addr[7:7] ;
assign n19330 =  ( n19329 ) == ( bv_1_0_n53 )  ;
assign n19331 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n19332 =  ( n19330 ) & (n19331 )  ;
assign n19333 =  ( n19332 ) & (wr )  ;
assign n19334 =  ( n19333 ) ? ( n5071 ) : ( iram_144 ) ;
assign n19335 = wr_addr[7:7] ;
assign n19336 =  ( n19335 ) == ( bv_1_0_n53 )  ;
assign n19337 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n19338 =  ( n19336 ) & (n19337 )  ;
assign n19339 =  ( n19338 ) & (wr )  ;
assign n19340 =  ( n19339 ) ? ( n5096 ) : ( iram_144 ) ;
assign n19341 = wr_addr[7:7] ;
assign n19342 =  ( n19341 ) == ( bv_1_0_n53 )  ;
assign n19343 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n19344 =  ( n19342 ) & (n19343 )  ;
assign n19345 =  ( n19344 ) & (wr )  ;
assign n19346 =  ( n19345 ) ? ( n5123 ) : ( iram_144 ) ;
assign n19347 = wr_addr[7:7] ;
assign n19348 =  ( n19347 ) == ( bv_1_0_n53 )  ;
assign n19349 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n19350 =  ( n19348 ) & (n19349 )  ;
assign n19351 =  ( n19350 ) & (wr )  ;
assign n19352 =  ( n19351 ) ? ( n5165 ) : ( iram_144 ) ;
assign n19353 = wr_addr[7:7] ;
assign n19354 =  ( n19353 ) == ( bv_1_0_n53 )  ;
assign n19355 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n19356 =  ( n19354 ) & (n19355 )  ;
assign n19357 =  ( n19356 ) & (wr )  ;
assign n19358 =  ( n19357 ) ? ( n5204 ) : ( iram_144 ) ;
assign n19359 = wr_addr[7:7] ;
assign n19360 =  ( n19359 ) == ( bv_1_0_n53 )  ;
assign n19361 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n19362 =  ( n19360 ) & (n19361 )  ;
assign n19363 =  ( n19362 ) & (wr )  ;
assign n19364 =  ( n19363 ) ? ( n5262 ) : ( iram_144 ) ;
assign n19365 = wr_addr[7:7] ;
assign n19366 =  ( n19365 ) == ( bv_1_0_n53 )  ;
assign n19367 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n19368 =  ( n19366 ) & (n19367 )  ;
assign n19369 =  ( n19368 ) & (wr )  ;
assign n19370 =  ( n19369 ) ? ( n5298 ) : ( iram_144 ) ;
assign n19371 = wr_addr[7:7] ;
assign n19372 =  ( n19371 ) == ( bv_1_0_n53 )  ;
assign n19373 =  ( wr_addr ) == ( bv_8_144_n357 )  ;
assign n19374 =  ( n19372 ) & (n19373 )  ;
assign n19375 =  ( n19374 ) & (wr )  ;
assign n19376 =  ( n19375 ) ? ( n5325 ) : ( iram_144 ) ;
assign n19377 = wr_addr[7:7] ;
assign n19378 =  ( n19377 ) == ( bv_1_0_n53 )  ;
assign n19379 =  ( wr_addr ) == ( bv_8_145_n359 )  ;
assign n19380 =  ( n19378 ) & (n19379 )  ;
assign n19381 =  ( n19380 ) & (wr )  ;
assign n19382 =  ( n19381 ) ? ( n4782 ) : ( iram_145 ) ;
assign n19383 = wr_addr[7:7] ;
assign n19384 =  ( n19383 ) == ( bv_1_0_n53 )  ;
assign n19385 =  ( wr_addr ) == ( bv_8_145_n359 )  ;
assign n19386 =  ( n19384 ) & (n19385 )  ;
assign n19387 =  ( n19386 ) & (wr )  ;
assign n19388 =  ( n19387 ) ? ( n4841 ) : ( iram_145 ) ;
assign n19389 = wr_addr[7:7] ;
assign n19390 =  ( n19389 ) == ( bv_1_0_n53 )  ;
assign n19391 =  ( wr_addr ) == ( bv_8_145_n359 )  ;
assign n19392 =  ( n19390 ) & (n19391 )  ;
assign n19393 =  ( n19392 ) & (wr )  ;
assign n19394 =  ( n19393 ) ? ( n5449 ) : ( iram_145 ) ;
assign n19395 = wr_addr[7:7] ;
assign n19396 =  ( n19395 ) == ( bv_1_0_n53 )  ;
assign n19397 =  ( wr_addr ) == ( bv_8_145_n359 )  ;
assign n19398 =  ( n19396 ) & (n19397 )  ;
assign n19399 =  ( n19398 ) & (wr )  ;
assign n19400 =  ( n19399 ) ? ( n4906 ) : ( iram_145 ) ;
assign n19401 = wr_addr[7:7] ;
assign n19402 =  ( n19401 ) == ( bv_1_0_n53 )  ;
assign n19403 =  ( wr_addr ) == ( bv_8_145_n359 )  ;
assign n19404 =  ( n19402 ) & (n19403 )  ;
assign n19405 =  ( n19404 ) & (wr )  ;
assign n19406 =  ( n19405 ) ? ( n5485 ) : ( iram_145 ) ;
assign n19407 = wr_addr[7:7] ;
assign n19408 =  ( n19407 ) == ( bv_1_0_n53 )  ;
assign n19409 =  ( wr_addr ) == ( bv_8_145_n359 )  ;
assign n19410 =  ( n19408 ) & (n19409 )  ;
assign n19411 =  ( n19410 ) & (wr )  ;
assign n19412 =  ( n19411 ) ? ( n5512 ) : ( iram_145 ) ;
assign n19413 = wr_addr[7:7] ;
assign n19414 =  ( n19413 ) == ( bv_1_0_n53 )  ;
assign n19415 =  ( wr_addr ) == ( bv_8_145_n359 )  ;
assign n19416 =  ( n19414 ) & (n19415 )  ;
assign n19417 =  ( n19416 ) & (wr )  ;
assign n19418 =  ( n19417 ) ? ( bv_8_0_n69 ) : ( iram_145 ) ;
assign n19419 = wr_addr[7:7] ;
assign n19420 =  ( n19419 ) == ( bv_1_0_n53 )  ;
assign n19421 =  ( wr_addr ) == ( bv_8_145_n359 )  ;
assign n19422 =  ( n19420 ) & (n19421 )  ;
assign n19423 =  ( n19422 ) & (wr )  ;
assign n19424 =  ( n19423 ) ? ( n5071 ) : ( iram_145 ) ;
assign n19425 = wr_addr[7:7] ;
assign n19426 =  ( n19425 ) == ( bv_1_0_n53 )  ;
assign n19427 =  ( wr_addr ) == ( bv_8_145_n359 )  ;
assign n19428 =  ( n19426 ) & (n19427 )  ;
assign n19429 =  ( n19428 ) & (wr )  ;
assign n19430 =  ( n19429 ) ? ( n5096 ) : ( iram_145 ) ;
assign n19431 = wr_addr[7:7] ;
assign n19432 =  ( n19431 ) == ( bv_1_0_n53 )  ;
assign n19433 =  ( wr_addr ) == ( bv_8_145_n359 )  ;
assign n19434 =  ( n19432 ) & (n19433 )  ;
assign n19435 =  ( n19434 ) & (wr )  ;
assign n19436 =  ( n19435 ) ? ( n5123 ) : ( iram_145 ) ;
assign n19437 = wr_addr[7:7] ;
assign n19438 =  ( n19437 ) == ( bv_1_0_n53 )  ;
assign n19439 =  ( wr_addr ) == ( bv_8_145_n359 )  ;
assign n19440 =  ( n19438 ) & (n19439 )  ;
assign n19441 =  ( n19440 ) & (wr )  ;
assign n19442 =  ( n19441 ) ? ( n5165 ) : ( iram_145 ) ;
assign n19443 = wr_addr[7:7] ;
assign n19444 =  ( n19443 ) == ( bv_1_0_n53 )  ;
assign n19445 =  ( wr_addr ) == ( bv_8_145_n359 )  ;
assign n19446 =  ( n19444 ) & (n19445 )  ;
assign n19447 =  ( n19446 ) & (wr )  ;
assign n19448 =  ( n19447 ) ? ( n5204 ) : ( iram_145 ) ;
assign n19449 = wr_addr[7:7] ;
assign n19450 =  ( n19449 ) == ( bv_1_0_n53 )  ;
assign n19451 =  ( wr_addr ) == ( bv_8_145_n359 )  ;
assign n19452 =  ( n19450 ) & (n19451 )  ;
assign n19453 =  ( n19452 ) & (wr )  ;
assign n19454 =  ( n19453 ) ? ( n5262 ) : ( iram_145 ) ;
assign n19455 = wr_addr[7:7] ;
assign n19456 =  ( n19455 ) == ( bv_1_0_n53 )  ;
assign n19457 =  ( wr_addr ) == ( bv_8_145_n359 )  ;
assign n19458 =  ( n19456 ) & (n19457 )  ;
assign n19459 =  ( n19458 ) & (wr )  ;
assign n19460 =  ( n19459 ) ? ( n5298 ) : ( iram_145 ) ;
assign n19461 = wr_addr[7:7] ;
assign n19462 =  ( n19461 ) == ( bv_1_0_n53 )  ;
assign n19463 =  ( wr_addr ) == ( bv_8_145_n359 )  ;
assign n19464 =  ( n19462 ) & (n19463 )  ;
assign n19465 =  ( n19464 ) & (wr )  ;
assign n19466 =  ( n19465 ) ? ( n5325 ) : ( iram_145 ) ;
assign n19467 = wr_addr[7:7] ;
assign n19468 =  ( n19467 ) == ( bv_1_0_n53 )  ;
assign n19469 =  ( wr_addr ) == ( bv_8_146_n361 )  ;
assign n19470 =  ( n19468 ) & (n19469 )  ;
assign n19471 =  ( n19470 ) & (wr )  ;
assign n19472 =  ( n19471 ) ? ( n4782 ) : ( iram_146 ) ;
assign n19473 = wr_addr[7:7] ;
assign n19474 =  ( n19473 ) == ( bv_1_0_n53 )  ;
assign n19475 =  ( wr_addr ) == ( bv_8_146_n361 )  ;
assign n19476 =  ( n19474 ) & (n19475 )  ;
assign n19477 =  ( n19476 ) & (wr )  ;
assign n19478 =  ( n19477 ) ? ( n4841 ) : ( iram_146 ) ;
assign n19479 = wr_addr[7:7] ;
assign n19480 =  ( n19479 ) == ( bv_1_0_n53 )  ;
assign n19481 =  ( wr_addr ) == ( bv_8_146_n361 )  ;
assign n19482 =  ( n19480 ) & (n19481 )  ;
assign n19483 =  ( n19482 ) & (wr )  ;
assign n19484 =  ( n19483 ) ? ( n5449 ) : ( iram_146 ) ;
assign n19485 = wr_addr[7:7] ;
assign n19486 =  ( n19485 ) == ( bv_1_0_n53 )  ;
assign n19487 =  ( wr_addr ) == ( bv_8_146_n361 )  ;
assign n19488 =  ( n19486 ) & (n19487 )  ;
assign n19489 =  ( n19488 ) & (wr )  ;
assign n19490 =  ( n19489 ) ? ( n4906 ) : ( iram_146 ) ;
assign n19491 = wr_addr[7:7] ;
assign n19492 =  ( n19491 ) == ( bv_1_0_n53 )  ;
assign n19493 =  ( wr_addr ) == ( bv_8_146_n361 )  ;
assign n19494 =  ( n19492 ) & (n19493 )  ;
assign n19495 =  ( n19494 ) & (wr )  ;
assign n19496 =  ( n19495 ) ? ( n5485 ) : ( iram_146 ) ;
assign n19497 = wr_addr[7:7] ;
assign n19498 =  ( n19497 ) == ( bv_1_0_n53 )  ;
assign n19499 =  ( wr_addr ) == ( bv_8_146_n361 )  ;
assign n19500 =  ( n19498 ) & (n19499 )  ;
assign n19501 =  ( n19500 ) & (wr )  ;
assign n19502 =  ( n19501 ) ? ( n5512 ) : ( iram_146 ) ;
assign n19503 = wr_addr[7:7] ;
assign n19504 =  ( n19503 ) == ( bv_1_0_n53 )  ;
assign n19505 =  ( wr_addr ) == ( bv_8_146_n361 )  ;
assign n19506 =  ( n19504 ) & (n19505 )  ;
assign n19507 =  ( n19506 ) & (wr )  ;
assign n19508 =  ( n19507 ) ? ( bv_8_0_n69 ) : ( iram_146 ) ;
assign n19509 = wr_addr[7:7] ;
assign n19510 =  ( n19509 ) == ( bv_1_0_n53 )  ;
assign n19511 =  ( wr_addr ) == ( bv_8_146_n361 )  ;
assign n19512 =  ( n19510 ) & (n19511 )  ;
assign n19513 =  ( n19512 ) & (wr )  ;
assign n19514 =  ( n19513 ) ? ( n5071 ) : ( iram_146 ) ;
assign n19515 = wr_addr[7:7] ;
assign n19516 =  ( n19515 ) == ( bv_1_0_n53 )  ;
assign n19517 =  ( wr_addr ) == ( bv_8_146_n361 )  ;
assign n19518 =  ( n19516 ) & (n19517 )  ;
assign n19519 =  ( n19518 ) & (wr )  ;
assign n19520 =  ( n19519 ) ? ( n5096 ) : ( iram_146 ) ;
assign n19521 = wr_addr[7:7] ;
assign n19522 =  ( n19521 ) == ( bv_1_0_n53 )  ;
assign n19523 =  ( wr_addr ) == ( bv_8_146_n361 )  ;
assign n19524 =  ( n19522 ) & (n19523 )  ;
assign n19525 =  ( n19524 ) & (wr )  ;
assign n19526 =  ( n19525 ) ? ( n5123 ) : ( iram_146 ) ;
assign n19527 = wr_addr[7:7] ;
assign n19528 =  ( n19527 ) == ( bv_1_0_n53 )  ;
assign n19529 =  ( wr_addr ) == ( bv_8_146_n361 )  ;
assign n19530 =  ( n19528 ) & (n19529 )  ;
assign n19531 =  ( n19530 ) & (wr )  ;
assign n19532 =  ( n19531 ) ? ( n5165 ) : ( iram_146 ) ;
assign n19533 = wr_addr[7:7] ;
assign n19534 =  ( n19533 ) == ( bv_1_0_n53 )  ;
assign n19535 =  ( wr_addr ) == ( bv_8_146_n361 )  ;
assign n19536 =  ( n19534 ) & (n19535 )  ;
assign n19537 =  ( n19536 ) & (wr )  ;
assign n19538 =  ( n19537 ) ? ( n5204 ) : ( iram_146 ) ;
assign n19539 = wr_addr[7:7] ;
assign n19540 =  ( n19539 ) == ( bv_1_0_n53 )  ;
assign n19541 =  ( wr_addr ) == ( bv_8_146_n361 )  ;
assign n19542 =  ( n19540 ) & (n19541 )  ;
assign n19543 =  ( n19542 ) & (wr )  ;
assign n19544 =  ( n19543 ) ? ( n5262 ) : ( iram_146 ) ;
assign n19545 = wr_addr[7:7] ;
assign n19546 =  ( n19545 ) == ( bv_1_0_n53 )  ;
assign n19547 =  ( wr_addr ) == ( bv_8_146_n361 )  ;
assign n19548 =  ( n19546 ) & (n19547 )  ;
assign n19549 =  ( n19548 ) & (wr )  ;
assign n19550 =  ( n19549 ) ? ( n5298 ) : ( iram_146 ) ;
assign n19551 = wr_addr[7:7] ;
assign n19552 =  ( n19551 ) == ( bv_1_0_n53 )  ;
assign n19553 =  ( wr_addr ) == ( bv_8_146_n361 )  ;
assign n19554 =  ( n19552 ) & (n19553 )  ;
assign n19555 =  ( n19554 ) & (wr )  ;
assign n19556 =  ( n19555 ) ? ( n5325 ) : ( iram_146 ) ;
assign n19557 = wr_addr[7:7] ;
assign n19558 =  ( n19557 ) == ( bv_1_0_n53 )  ;
assign n19559 =  ( wr_addr ) == ( bv_8_147_n363 )  ;
assign n19560 =  ( n19558 ) & (n19559 )  ;
assign n19561 =  ( n19560 ) & (wr )  ;
assign n19562 =  ( n19561 ) ? ( n4782 ) : ( iram_147 ) ;
assign n19563 = wr_addr[7:7] ;
assign n19564 =  ( n19563 ) == ( bv_1_0_n53 )  ;
assign n19565 =  ( wr_addr ) == ( bv_8_147_n363 )  ;
assign n19566 =  ( n19564 ) & (n19565 )  ;
assign n19567 =  ( n19566 ) & (wr )  ;
assign n19568 =  ( n19567 ) ? ( n4841 ) : ( iram_147 ) ;
assign n19569 = wr_addr[7:7] ;
assign n19570 =  ( n19569 ) == ( bv_1_0_n53 )  ;
assign n19571 =  ( wr_addr ) == ( bv_8_147_n363 )  ;
assign n19572 =  ( n19570 ) & (n19571 )  ;
assign n19573 =  ( n19572 ) & (wr )  ;
assign n19574 =  ( n19573 ) ? ( n5449 ) : ( iram_147 ) ;
assign n19575 = wr_addr[7:7] ;
assign n19576 =  ( n19575 ) == ( bv_1_0_n53 )  ;
assign n19577 =  ( wr_addr ) == ( bv_8_147_n363 )  ;
assign n19578 =  ( n19576 ) & (n19577 )  ;
assign n19579 =  ( n19578 ) & (wr )  ;
assign n19580 =  ( n19579 ) ? ( n4906 ) : ( iram_147 ) ;
assign n19581 = wr_addr[7:7] ;
assign n19582 =  ( n19581 ) == ( bv_1_0_n53 )  ;
assign n19583 =  ( wr_addr ) == ( bv_8_147_n363 )  ;
assign n19584 =  ( n19582 ) & (n19583 )  ;
assign n19585 =  ( n19584 ) & (wr )  ;
assign n19586 =  ( n19585 ) ? ( n5485 ) : ( iram_147 ) ;
assign n19587 = wr_addr[7:7] ;
assign n19588 =  ( n19587 ) == ( bv_1_0_n53 )  ;
assign n19589 =  ( wr_addr ) == ( bv_8_147_n363 )  ;
assign n19590 =  ( n19588 ) & (n19589 )  ;
assign n19591 =  ( n19590 ) & (wr )  ;
assign n19592 =  ( n19591 ) ? ( n5512 ) : ( iram_147 ) ;
assign n19593 = wr_addr[7:7] ;
assign n19594 =  ( n19593 ) == ( bv_1_0_n53 )  ;
assign n19595 =  ( wr_addr ) == ( bv_8_147_n363 )  ;
assign n19596 =  ( n19594 ) & (n19595 )  ;
assign n19597 =  ( n19596 ) & (wr )  ;
assign n19598 =  ( n19597 ) ? ( bv_8_0_n69 ) : ( iram_147 ) ;
assign n19599 = wr_addr[7:7] ;
assign n19600 =  ( n19599 ) == ( bv_1_0_n53 )  ;
assign n19601 =  ( wr_addr ) == ( bv_8_147_n363 )  ;
assign n19602 =  ( n19600 ) & (n19601 )  ;
assign n19603 =  ( n19602 ) & (wr )  ;
assign n19604 =  ( n19603 ) ? ( n5071 ) : ( iram_147 ) ;
assign n19605 = wr_addr[7:7] ;
assign n19606 =  ( n19605 ) == ( bv_1_0_n53 )  ;
assign n19607 =  ( wr_addr ) == ( bv_8_147_n363 )  ;
assign n19608 =  ( n19606 ) & (n19607 )  ;
assign n19609 =  ( n19608 ) & (wr )  ;
assign n19610 =  ( n19609 ) ? ( n5096 ) : ( iram_147 ) ;
assign n19611 = wr_addr[7:7] ;
assign n19612 =  ( n19611 ) == ( bv_1_0_n53 )  ;
assign n19613 =  ( wr_addr ) == ( bv_8_147_n363 )  ;
assign n19614 =  ( n19612 ) & (n19613 )  ;
assign n19615 =  ( n19614 ) & (wr )  ;
assign n19616 =  ( n19615 ) ? ( n5123 ) : ( iram_147 ) ;
assign n19617 = wr_addr[7:7] ;
assign n19618 =  ( n19617 ) == ( bv_1_0_n53 )  ;
assign n19619 =  ( wr_addr ) == ( bv_8_147_n363 )  ;
assign n19620 =  ( n19618 ) & (n19619 )  ;
assign n19621 =  ( n19620 ) & (wr )  ;
assign n19622 =  ( n19621 ) ? ( n5165 ) : ( iram_147 ) ;
assign n19623 = wr_addr[7:7] ;
assign n19624 =  ( n19623 ) == ( bv_1_0_n53 )  ;
assign n19625 =  ( wr_addr ) == ( bv_8_147_n363 )  ;
assign n19626 =  ( n19624 ) & (n19625 )  ;
assign n19627 =  ( n19626 ) & (wr )  ;
assign n19628 =  ( n19627 ) ? ( n5204 ) : ( iram_147 ) ;
assign n19629 = wr_addr[7:7] ;
assign n19630 =  ( n19629 ) == ( bv_1_0_n53 )  ;
assign n19631 =  ( wr_addr ) == ( bv_8_147_n363 )  ;
assign n19632 =  ( n19630 ) & (n19631 )  ;
assign n19633 =  ( n19632 ) & (wr )  ;
assign n19634 =  ( n19633 ) ? ( n5262 ) : ( iram_147 ) ;
assign n19635 = wr_addr[7:7] ;
assign n19636 =  ( n19635 ) == ( bv_1_0_n53 )  ;
assign n19637 =  ( wr_addr ) == ( bv_8_147_n363 )  ;
assign n19638 =  ( n19636 ) & (n19637 )  ;
assign n19639 =  ( n19638 ) & (wr )  ;
assign n19640 =  ( n19639 ) ? ( n5298 ) : ( iram_147 ) ;
assign n19641 = wr_addr[7:7] ;
assign n19642 =  ( n19641 ) == ( bv_1_0_n53 )  ;
assign n19643 =  ( wr_addr ) == ( bv_8_147_n363 )  ;
assign n19644 =  ( n19642 ) & (n19643 )  ;
assign n19645 =  ( n19644 ) & (wr )  ;
assign n19646 =  ( n19645 ) ? ( n5325 ) : ( iram_147 ) ;
assign n19647 = wr_addr[7:7] ;
assign n19648 =  ( n19647 ) == ( bv_1_0_n53 )  ;
assign n19649 =  ( wr_addr ) == ( bv_8_148_n365 )  ;
assign n19650 =  ( n19648 ) & (n19649 )  ;
assign n19651 =  ( n19650 ) & (wr )  ;
assign n19652 =  ( n19651 ) ? ( n4782 ) : ( iram_148 ) ;
assign n19653 = wr_addr[7:7] ;
assign n19654 =  ( n19653 ) == ( bv_1_0_n53 )  ;
assign n19655 =  ( wr_addr ) == ( bv_8_148_n365 )  ;
assign n19656 =  ( n19654 ) & (n19655 )  ;
assign n19657 =  ( n19656 ) & (wr )  ;
assign n19658 =  ( n19657 ) ? ( n4841 ) : ( iram_148 ) ;
assign n19659 = wr_addr[7:7] ;
assign n19660 =  ( n19659 ) == ( bv_1_0_n53 )  ;
assign n19661 =  ( wr_addr ) == ( bv_8_148_n365 )  ;
assign n19662 =  ( n19660 ) & (n19661 )  ;
assign n19663 =  ( n19662 ) & (wr )  ;
assign n19664 =  ( n19663 ) ? ( n5449 ) : ( iram_148 ) ;
assign n19665 = wr_addr[7:7] ;
assign n19666 =  ( n19665 ) == ( bv_1_0_n53 )  ;
assign n19667 =  ( wr_addr ) == ( bv_8_148_n365 )  ;
assign n19668 =  ( n19666 ) & (n19667 )  ;
assign n19669 =  ( n19668 ) & (wr )  ;
assign n19670 =  ( n19669 ) ? ( n4906 ) : ( iram_148 ) ;
assign n19671 = wr_addr[7:7] ;
assign n19672 =  ( n19671 ) == ( bv_1_0_n53 )  ;
assign n19673 =  ( wr_addr ) == ( bv_8_148_n365 )  ;
assign n19674 =  ( n19672 ) & (n19673 )  ;
assign n19675 =  ( n19674 ) & (wr )  ;
assign n19676 =  ( n19675 ) ? ( n5485 ) : ( iram_148 ) ;
assign n19677 = wr_addr[7:7] ;
assign n19678 =  ( n19677 ) == ( bv_1_0_n53 )  ;
assign n19679 =  ( wr_addr ) == ( bv_8_148_n365 )  ;
assign n19680 =  ( n19678 ) & (n19679 )  ;
assign n19681 =  ( n19680 ) & (wr )  ;
assign n19682 =  ( n19681 ) ? ( n5512 ) : ( iram_148 ) ;
assign n19683 = wr_addr[7:7] ;
assign n19684 =  ( n19683 ) == ( bv_1_0_n53 )  ;
assign n19685 =  ( wr_addr ) == ( bv_8_148_n365 )  ;
assign n19686 =  ( n19684 ) & (n19685 )  ;
assign n19687 =  ( n19686 ) & (wr )  ;
assign n19688 =  ( n19687 ) ? ( bv_8_0_n69 ) : ( iram_148 ) ;
assign n19689 = wr_addr[7:7] ;
assign n19690 =  ( n19689 ) == ( bv_1_0_n53 )  ;
assign n19691 =  ( wr_addr ) == ( bv_8_148_n365 )  ;
assign n19692 =  ( n19690 ) & (n19691 )  ;
assign n19693 =  ( n19692 ) & (wr )  ;
assign n19694 =  ( n19693 ) ? ( n5071 ) : ( iram_148 ) ;
assign n19695 = wr_addr[7:7] ;
assign n19696 =  ( n19695 ) == ( bv_1_0_n53 )  ;
assign n19697 =  ( wr_addr ) == ( bv_8_148_n365 )  ;
assign n19698 =  ( n19696 ) & (n19697 )  ;
assign n19699 =  ( n19698 ) & (wr )  ;
assign n19700 =  ( n19699 ) ? ( n5096 ) : ( iram_148 ) ;
assign n19701 = wr_addr[7:7] ;
assign n19702 =  ( n19701 ) == ( bv_1_0_n53 )  ;
assign n19703 =  ( wr_addr ) == ( bv_8_148_n365 )  ;
assign n19704 =  ( n19702 ) & (n19703 )  ;
assign n19705 =  ( n19704 ) & (wr )  ;
assign n19706 =  ( n19705 ) ? ( n5123 ) : ( iram_148 ) ;
assign n19707 = wr_addr[7:7] ;
assign n19708 =  ( n19707 ) == ( bv_1_0_n53 )  ;
assign n19709 =  ( wr_addr ) == ( bv_8_148_n365 )  ;
assign n19710 =  ( n19708 ) & (n19709 )  ;
assign n19711 =  ( n19710 ) & (wr )  ;
assign n19712 =  ( n19711 ) ? ( n5165 ) : ( iram_148 ) ;
assign n19713 = wr_addr[7:7] ;
assign n19714 =  ( n19713 ) == ( bv_1_0_n53 )  ;
assign n19715 =  ( wr_addr ) == ( bv_8_148_n365 )  ;
assign n19716 =  ( n19714 ) & (n19715 )  ;
assign n19717 =  ( n19716 ) & (wr )  ;
assign n19718 =  ( n19717 ) ? ( n5204 ) : ( iram_148 ) ;
assign n19719 = wr_addr[7:7] ;
assign n19720 =  ( n19719 ) == ( bv_1_0_n53 )  ;
assign n19721 =  ( wr_addr ) == ( bv_8_148_n365 )  ;
assign n19722 =  ( n19720 ) & (n19721 )  ;
assign n19723 =  ( n19722 ) & (wr )  ;
assign n19724 =  ( n19723 ) ? ( n5262 ) : ( iram_148 ) ;
assign n19725 = wr_addr[7:7] ;
assign n19726 =  ( n19725 ) == ( bv_1_0_n53 )  ;
assign n19727 =  ( wr_addr ) == ( bv_8_148_n365 )  ;
assign n19728 =  ( n19726 ) & (n19727 )  ;
assign n19729 =  ( n19728 ) & (wr )  ;
assign n19730 =  ( n19729 ) ? ( n5298 ) : ( iram_148 ) ;
assign n19731 = wr_addr[7:7] ;
assign n19732 =  ( n19731 ) == ( bv_1_0_n53 )  ;
assign n19733 =  ( wr_addr ) == ( bv_8_148_n365 )  ;
assign n19734 =  ( n19732 ) & (n19733 )  ;
assign n19735 =  ( n19734 ) & (wr )  ;
assign n19736 =  ( n19735 ) ? ( n5325 ) : ( iram_148 ) ;
assign n19737 = wr_addr[7:7] ;
assign n19738 =  ( n19737 ) == ( bv_1_0_n53 )  ;
assign n19739 =  ( wr_addr ) == ( bv_8_149_n367 )  ;
assign n19740 =  ( n19738 ) & (n19739 )  ;
assign n19741 =  ( n19740 ) & (wr )  ;
assign n19742 =  ( n19741 ) ? ( n4782 ) : ( iram_149 ) ;
assign n19743 = wr_addr[7:7] ;
assign n19744 =  ( n19743 ) == ( bv_1_0_n53 )  ;
assign n19745 =  ( wr_addr ) == ( bv_8_149_n367 )  ;
assign n19746 =  ( n19744 ) & (n19745 )  ;
assign n19747 =  ( n19746 ) & (wr )  ;
assign n19748 =  ( n19747 ) ? ( n4841 ) : ( iram_149 ) ;
assign n19749 = wr_addr[7:7] ;
assign n19750 =  ( n19749 ) == ( bv_1_0_n53 )  ;
assign n19751 =  ( wr_addr ) == ( bv_8_149_n367 )  ;
assign n19752 =  ( n19750 ) & (n19751 )  ;
assign n19753 =  ( n19752 ) & (wr )  ;
assign n19754 =  ( n19753 ) ? ( n5449 ) : ( iram_149 ) ;
assign n19755 = wr_addr[7:7] ;
assign n19756 =  ( n19755 ) == ( bv_1_0_n53 )  ;
assign n19757 =  ( wr_addr ) == ( bv_8_149_n367 )  ;
assign n19758 =  ( n19756 ) & (n19757 )  ;
assign n19759 =  ( n19758 ) & (wr )  ;
assign n19760 =  ( n19759 ) ? ( n4906 ) : ( iram_149 ) ;
assign n19761 = wr_addr[7:7] ;
assign n19762 =  ( n19761 ) == ( bv_1_0_n53 )  ;
assign n19763 =  ( wr_addr ) == ( bv_8_149_n367 )  ;
assign n19764 =  ( n19762 ) & (n19763 )  ;
assign n19765 =  ( n19764 ) & (wr )  ;
assign n19766 =  ( n19765 ) ? ( n5485 ) : ( iram_149 ) ;
assign n19767 = wr_addr[7:7] ;
assign n19768 =  ( n19767 ) == ( bv_1_0_n53 )  ;
assign n19769 =  ( wr_addr ) == ( bv_8_149_n367 )  ;
assign n19770 =  ( n19768 ) & (n19769 )  ;
assign n19771 =  ( n19770 ) & (wr )  ;
assign n19772 =  ( n19771 ) ? ( n5512 ) : ( iram_149 ) ;
assign n19773 = wr_addr[7:7] ;
assign n19774 =  ( n19773 ) == ( bv_1_0_n53 )  ;
assign n19775 =  ( wr_addr ) == ( bv_8_149_n367 )  ;
assign n19776 =  ( n19774 ) & (n19775 )  ;
assign n19777 =  ( n19776 ) & (wr )  ;
assign n19778 =  ( n19777 ) ? ( bv_8_0_n69 ) : ( iram_149 ) ;
assign n19779 = wr_addr[7:7] ;
assign n19780 =  ( n19779 ) == ( bv_1_0_n53 )  ;
assign n19781 =  ( wr_addr ) == ( bv_8_149_n367 )  ;
assign n19782 =  ( n19780 ) & (n19781 )  ;
assign n19783 =  ( n19782 ) & (wr )  ;
assign n19784 =  ( n19783 ) ? ( n5071 ) : ( iram_149 ) ;
assign n19785 = wr_addr[7:7] ;
assign n19786 =  ( n19785 ) == ( bv_1_0_n53 )  ;
assign n19787 =  ( wr_addr ) == ( bv_8_149_n367 )  ;
assign n19788 =  ( n19786 ) & (n19787 )  ;
assign n19789 =  ( n19788 ) & (wr )  ;
assign n19790 =  ( n19789 ) ? ( n5096 ) : ( iram_149 ) ;
assign n19791 = wr_addr[7:7] ;
assign n19792 =  ( n19791 ) == ( bv_1_0_n53 )  ;
assign n19793 =  ( wr_addr ) == ( bv_8_149_n367 )  ;
assign n19794 =  ( n19792 ) & (n19793 )  ;
assign n19795 =  ( n19794 ) & (wr )  ;
assign n19796 =  ( n19795 ) ? ( n5123 ) : ( iram_149 ) ;
assign n19797 = wr_addr[7:7] ;
assign n19798 =  ( n19797 ) == ( bv_1_0_n53 )  ;
assign n19799 =  ( wr_addr ) == ( bv_8_149_n367 )  ;
assign n19800 =  ( n19798 ) & (n19799 )  ;
assign n19801 =  ( n19800 ) & (wr )  ;
assign n19802 =  ( n19801 ) ? ( n5165 ) : ( iram_149 ) ;
assign n19803 = wr_addr[7:7] ;
assign n19804 =  ( n19803 ) == ( bv_1_0_n53 )  ;
assign n19805 =  ( wr_addr ) == ( bv_8_149_n367 )  ;
assign n19806 =  ( n19804 ) & (n19805 )  ;
assign n19807 =  ( n19806 ) & (wr )  ;
assign n19808 =  ( n19807 ) ? ( n5204 ) : ( iram_149 ) ;
assign n19809 = wr_addr[7:7] ;
assign n19810 =  ( n19809 ) == ( bv_1_0_n53 )  ;
assign n19811 =  ( wr_addr ) == ( bv_8_149_n367 )  ;
assign n19812 =  ( n19810 ) & (n19811 )  ;
assign n19813 =  ( n19812 ) & (wr )  ;
assign n19814 =  ( n19813 ) ? ( n5262 ) : ( iram_149 ) ;
assign n19815 = wr_addr[7:7] ;
assign n19816 =  ( n19815 ) == ( bv_1_0_n53 )  ;
assign n19817 =  ( wr_addr ) == ( bv_8_149_n367 )  ;
assign n19818 =  ( n19816 ) & (n19817 )  ;
assign n19819 =  ( n19818 ) & (wr )  ;
assign n19820 =  ( n19819 ) ? ( n5298 ) : ( iram_149 ) ;
assign n19821 = wr_addr[7:7] ;
assign n19822 =  ( n19821 ) == ( bv_1_0_n53 )  ;
assign n19823 =  ( wr_addr ) == ( bv_8_149_n367 )  ;
assign n19824 =  ( n19822 ) & (n19823 )  ;
assign n19825 =  ( n19824 ) & (wr )  ;
assign n19826 =  ( n19825 ) ? ( n5325 ) : ( iram_149 ) ;
assign n19827 = wr_addr[7:7] ;
assign n19828 =  ( n19827 ) == ( bv_1_0_n53 )  ;
assign n19829 =  ( wr_addr ) == ( bv_8_150_n369 )  ;
assign n19830 =  ( n19828 ) & (n19829 )  ;
assign n19831 =  ( n19830 ) & (wr )  ;
assign n19832 =  ( n19831 ) ? ( n4782 ) : ( iram_150 ) ;
assign n19833 = wr_addr[7:7] ;
assign n19834 =  ( n19833 ) == ( bv_1_0_n53 )  ;
assign n19835 =  ( wr_addr ) == ( bv_8_150_n369 )  ;
assign n19836 =  ( n19834 ) & (n19835 )  ;
assign n19837 =  ( n19836 ) & (wr )  ;
assign n19838 =  ( n19837 ) ? ( n4841 ) : ( iram_150 ) ;
assign n19839 = wr_addr[7:7] ;
assign n19840 =  ( n19839 ) == ( bv_1_0_n53 )  ;
assign n19841 =  ( wr_addr ) == ( bv_8_150_n369 )  ;
assign n19842 =  ( n19840 ) & (n19841 )  ;
assign n19843 =  ( n19842 ) & (wr )  ;
assign n19844 =  ( n19843 ) ? ( n5449 ) : ( iram_150 ) ;
assign n19845 = wr_addr[7:7] ;
assign n19846 =  ( n19845 ) == ( bv_1_0_n53 )  ;
assign n19847 =  ( wr_addr ) == ( bv_8_150_n369 )  ;
assign n19848 =  ( n19846 ) & (n19847 )  ;
assign n19849 =  ( n19848 ) & (wr )  ;
assign n19850 =  ( n19849 ) ? ( n4906 ) : ( iram_150 ) ;
assign n19851 = wr_addr[7:7] ;
assign n19852 =  ( n19851 ) == ( bv_1_0_n53 )  ;
assign n19853 =  ( wr_addr ) == ( bv_8_150_n369 )  ;
assign n19854 =  ( n19852 ) & (n19853 )  ;
assign n19855 =  ( n19854 ) & (wr )  ;
assign n19856 =  ( n19855 ) ? ( n5485 ) : ( iram_150 ) ;
assign n19857 = wr_addr[7:7] ;
assign n19858 =  ( n19857 ) == ( bv_1_0_n53 )  ;
assign n19859 =  ( wr_addr ) == ( bv_8_150_n369 )  ;
assign n19860 =  ( n19858 ) & (n19859 )  ;
assign n19861 =  ( n19860 ) & (wr )  ;
assign n19862 =  ( n19861 ) ? ( n5512 ) : ( iram_150 ) ;
assign n19863 = wr_addr[7:7] ;
assign n19864 =  ( n19863 ) == ( bv_1_0_n53 )  ;
assign n19865 =  ( wr_addr ) == ( bv_8_150_n369 )  ;
assign n19866 =  ( n19864 ) & (n19865 )  ;
assign n19867 =  ( n19866 ) & (wr )  ;
assign n19868 =  ( n19867 ) ? ( bv_8_0_n69 ) : ( iram_150 ) ;
assign n19869 = wr_addr[7:7] ;
assign n19870 =  ( n19869 ) == ( bv_1_0_n53 )  ;
assign n19871 =  ( wr_addr ) == ( bv_8_150_n369 )  ;
assign n19872 =  ( n19870 ) & (n19871 )  ;
assign n19873 =  ( n19872 ) & (wr )  ;
assign n19874 =  ( n19873 ) ? ( n5071 ) : ( iram_150 ) ;
assign n19875 = wr_addr[7:7] ;
assign n19876 =  ( n19875 ) == ( bv_1_0_n53 )  ;
assign n19877 =  ( wr_addr ) == ( bv_8_150_n369 )  ;
assign n19878 =  ( n19876 ) & (n19877 )  ;
assign n19879 =  ( n19878 ) & (wr )  ;
assign n19880 =  ( n19879 ) ? ( n5096 ) : ( iram_150 ) ;
assign n19881 = wr_addr[7:7] ;
assign n19882 =  ( n19881 ) == ( bv_1_0_n53 )  ;
assign n19883 =  ( wr_addr ) == ( bv_8_150_n369 )  ;
assign n19884 =  ( n19882 ) & (n19883 )  ;
assign n19885 =  ( n19884 ) & (wr )  ;
assign n19886 =  ( n19885 ) ? ( n5123 ) : ( iram_150 ) ;
assign n19887 = wr_addr[7:7] ;
assign n19888 =  ( n19887 ) == ( bv_1_0_n53 )  ;
assign n19889 =  ( wr_addr ) == ( bv_8_150_n369 )  ;
assign n19890 =  ( n19888 ) & (n19889 )  ;
assign n19891 =  ( n19890 ) & (wr )  ;
assign n19892 =  ( n19891 ) ? ( n5165 ) : ( iram_150 ) ;
assign n19893 = wr_addr[7:7] ;
assign n19894 =  ( n19893 ) == ( bv_1_0_n53 )  ;
assign n19895 =  ( wr_addr ) == ( bv_8_150_n369 )  ;
assign n19896 =  ( n19894 ) & (n19895 )  ;
assign n19897 =  ( n19896 ) & (wr )  ;
assign n19898 =  ( n19897 ) ? ( n5204 ) : ( iram_150 ) ;
assign n19899 = wr_addr[7:7] ;
assign n19900 =  ( n19899 ) == ( bv_1_0_n53 )  ;
assign n19901 =  ( wr_addr ) == ( bv_8_150_n369 )  ;
assign n19902 =  ( n19900 ) & (n19901 )  ;
assign n19903 =  ( n19902 ) & (wr )  ;
assign n19904 =  ( n19903 ) ? ( n5262 ) : ( iram_150 ) ;
assign n19905 = wr_addr[7:7] ;
assign n19906 =  ( n19905 ) == ( bv_1_0_n53 )  ;
assign n19907 =  ( wr_addr ) == ( bv_8_150_n369 )  ;
assign n19908 =  ( n19906 ) & (n19907 )  ;
assign n19909 =  ( n19908 ) & (wr )  ;
assign n19910 =  ( n19909 ) ? ( n5298 ) : ( iram_150 ) ;
assign n19911 = wr_addr[7:7] ;
assign n19912 =  ( n19911 ) == ( bv_1_0_n53 )  ;
assign n19913 =  ( wr_addr ) == ( bv_8_150_n369 )  ;
assign n19914 =  ( n19912 ) & (n19913 )  ;
assign n19915 =  ( n19914 ) & (wr )  ;
assign n19916 =  ( n19915 ) ? ( n5325 ) : ( iram_150 ) ;
assign n19917 = wr_addr[7:7] ;
assign n19918 =  ( n19917 ) == ( bv_1_0_n53 )  ;
assign n19919 =  ( wr_addr ) == ( bv_8_151_n371 )  ;
assign n19920 =  ( n19918 ) & (n19919 )  ;
assign n19921 =  ( n19920 ) & (wr )  ;
assign n19922 =  ( n19921 ) ? ( n4782 ) : ( iram_151 ) ;
assign n19923 = wr_addr[7:7] ;
assign n19924 =  ( n19923 ) == ( bv_1_0_n53 )  ;
assign n19925 =  ( wr_addr ) == ( bv_8_151_n371 )  ;
assign n19926 =  ( n19924 ) & (n19925 )  ;
assign n19927 =  ( n19926 ) & (wr )  ;
assign n19928 =  ( n19927 ) ? ( n4841 ) : ( iram_151 ) ;
assign n19929 = wr_addr[7:7] ;
assign n19930 =  ( n19929 ) == ( bv_1_0_n53 )  ;
assign n19931 =  ( wr_addr ) == ( bv_8_151_n371 )  ;
assign n19932 =  ( n19930 ) & (n19931 )  ;
assign n19933 =  ( n19932 ) & (wr )  ;
assign n19934 =  ( n19933 ) ? ( n5449 ) : ( iram_151 ) ;
assign n19935 = wr_addr[7:7] ;
assign n19936 =  ( n19935 ) == ( bv_1_0_n53 )  ;
assign n19937 =  ( wr_addr ) == ( bv_8_151_n371 )  ;
assign n19938 =  ( n19936 ) & (n19937 )  ;
assign n19939 =  ( n19938 ) & (wr )  ;
assign n19940 =  ( n19939 ) ? ( n4906 ) : ( iram_151 ) ;
assign n19941 = wr_addr[7:7] ;
assign n19942 =  ( n19941 ) == ( bv_1_0_n53 )  ;
assign n19943 =  ( wr_addr ) == ( bv_8_151_n371 )  ;
assign n19944 =  ( n19942 ) & (n19943 )  ;
assign n19945 =  ( n19944 ) & (wr )  ;
assign n19946 =  ( n19945 ) ? ( n5485 ) : ( iram_151 ) ;
assign n19947 = wr_addr[7:7] ;
assign n19948 =  ( n19947 ) == ( bv_1_0_n53 )  ;
assign n19949 =  ( wr_addr ) == ( bv_8_151_n371 )  ;
assign n19950 =  ( n19948 ) & (n19949 )  ;
assign n19951 =  ( n19950 ) & (wr )  ;
assign n19952 =  ( n19951 ) ? ( n5512 ) : ( iram_151 ) ;
assign n19953 = wr_addr[7:7] ;
assign n19954 =  ( n19953 ) == ( bv_1_0_n53 )  ;
assign n19955 =  ( wr_addr ) == ( bv_8_151_n371 )  ;
assign n19956 =  ( n19954 ) & (n19955 )  ;
assign n19957 =  ( n19956 ) & (wr )  ;
assign n19958 =  ( n19957 ) ? ( bv_8_0_n69 ) : ( iram_151 ) ;
assign n19959 = wr_addr[7:7] ;
assign n19960 =  ( n19959 ) == ( bv_1_0_n53 )  ;
assign n19961 =  ( wr_addr ) == ( bv_8_151_n371 )  ;
assign n19962 =  ( n19960 ) & (n19961 )  ;
assign n19963 =  ( n19962 ) & (wr )  ;
assign n19964 =  ( n19963 ) ? ( n5071 ) : ( iram_151 ) ;
assign n19965 = wr_addr[7:7] ;
assign n19966 =  ( n19965 ) == ( bv_1_0_n53 )  ;
assign n19967 =  ( wr_addr ) == ( bv_8_151_n371 )  ;
assign n19968 =  ( n19966 ) & (n19967 )  ;
assign n19969 =  ( n19968 ) & (wr )  ;
assign n19970 =  ( n19969 ) ? ( n5096 ) : ( iram_151 ) ;
assign n19971 = wr_addr[7:7] ;
assign n19972 =  ( n19971 ) == ( bv_1_0_n53 )  ;
assign n19973 =  ( wr_addr ) == ( bv_8_151_n371 )  ;
assign n19974 =  ( n19972 ) & (n19973 )  ;
assign n19975 =  ( n19974 ) & (wr )  ;
assign n19976 =  ( n19975 ) ? ( n5123 ) : ( iram_151 ) ;
assign n19977 = wr_addr[7:7] ;
assign n19978 =  ( n19977 ) == ( bv_1_0_n53 )  ;
assign n19979 =  ( wr_addr ) == ( bv_8_151_n371 )  ;
assign n19980 =  ( n19978 ) & (n19979 )  ;
assign n19981 =  ( n19980 ) & (wr )  ;
assign n19982 =  ( n19981 ) ? ( n5165 ) : ( iram_151 ) ;
assign n19983 = wr_addr[7:7] ;
assign n19984 =  ( n19983 ) == ( bv_1_0_n53 )  ;
assign n19985 =  ( wr_addr ) == ( bv_8_151_n371 )  ;
assign n19986 =  ( n19984 ) & (n19985 )  ;
assign n19987 =  ( n19986 ) & (wr )  ;
assign n19988 =  ( n19987 ) ? ( n5204 ) : ( iram_151 ) ;
assign n19989 = wr_addr[7:7] ;
assign n19990 =  ( n19989 ) == ( bv_1_0_n53 )  ;
assign n19991 =  ( wr_addr ) == ( bv_8_151_n371 )  ;
assign n19992 =  ( n19990 ) & (n19991 )  ;
assign n19993 =  ( n19992 ) & (wr )  ;
assign n19994 =  ( n19993 ) ? ( n5262 ) : ( iram_151 ) ;
assign n19995 = wr_addr[7:7] ;
assign n19996 =  ( n19995 ) == ( bv_1_0_n53 )  ;
assign n19997 =  ( wr_addr ) == ( bv_8_151_n371 )  ;
assign n19998 =  ( n19996 ) & (n19997 )  ;
assign n19999 =  ( n19998 ) & (wr )  ;
assign n20000 =  ( n19999 ) ? ( n5298 ) : ( iram_151 ) ;
assign n20001 = wr_addr[7:7] ;
assign n20002 =  ( n20001 ) == ( bv_1_0_n53 )  ;
assign n20003 =  ( wr_addr ) == ( bv_8_151_n371 )  ;
assign n20004 =  ( n20002 ) & (n20003 )  ;
assign n20005 =  ( n20004 ) & (wr )  ;
assign n20006 =  ( n20005 ) ? ( n5325 ) : ( iram_151 ) ;
assign n20007 = wr_addr[7:7] ;
assign n20008 =  ( n20007 ) == ( bv_1_0_n53 )  ;
assign n20009 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n20010 =  ( n20008 ) & (n20009 )  ;
assign n20011 =  ( n20010 ) & (wr )  ;
assign n20012 =  ( n20011 ) ? ( n4782 ) : ( iram_152 ) ;
assign n20013 = wr_addr[7:7] ;
assign n20014 =  ( n20013 ) == ( bv_1_0_n53 )  ;
assign n20015 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n20016 =  ( n20014 ) & (n20015 )  ;
assign n20017 =  ( n20016 ) & (wr )  ;
assign n20018 =  ( n20017 ) ? ( n4841 ) : ( iram_152 ) ;
assign n20019 = wr_addr[7:7] ;
assign n20020 =  ( n20019 ) == ( bv_1_0_n53 )  ;
assign n20021 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n20022 =  ( n20020 ) & (n20021 )  ;
assign n20023 =  ( n20022 ) & (wr )  ;
assign n20024 =  ( n20023 ) ? ( n5449 ) : ( iram_152 ) ;
assign n20025 = wr_addr[7:7] ;
assign n20026 =  ( n20025 ) == ( bv_1_0_n53 )  ;
assign n20027 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n20028 =  ( n20026 ) & (n20027 )  ;
assign n20029 =  ( n20028 ) & (wr )  ;
assign n20030 =  ( n20029 ) ? ( n4906 ) : ( iram_152 ) ;
assign n20031 = wr_addr[7:7] ;
assign n20032 =  ( n20031 ) == ( bv_1_0_n53 )  ;
assign n20033 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n20034 =  ( n20032 ) & (n20033 )  ;
assign n20035 =  ( n20034 ) & (wr )  ;
assign n20036 =  ( n20035 ) ? ( n5485 ) : ( iram_152 ) ;
assign n20037 = wr_addr[7:7] ;
assign n20038 =  ( n20037 ) == ( bv_1_0_n53 )  ;
assign n20039 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n20040 =  ( n20038 ) & (n20039 )  ;
assign n20041 =  ( n20040 ) & (wr )  ;
assign n20042 =  ( n20041 ) ? ( n5512 ) : ( iram_152 ) ;
assign n20043 = wr_addr[7:7] ;
assign n20044 =  ( n20043 ) == ( bv_1_0_n53 )  ;
assign n20045 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n20046 =  ( n20044 ) & (n20045 )  ;
assign n20047 =  ( n20046 ) & (wr )  ;
assign n20048 =  ( n20047 ) ? ( bv_8_0_n69 ) : ( iram_152 ) ;
assign n20049 = wr_addr[7:7] ;
assign n20050 =  ( n20049 ) == ( bv_1_0_n53 )  ;
assign n20051 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n20052 =  ( n20050 ) & (n20051 )  ;
assign n20053 =  ( n20052 ) & (wr )  ;
assign n20054 =  ( n20053 ) ? ( n5071 ) : ( iram_152 ) ;
assign n20055 = wr_addr[7:7] ;
assign n20056 =  ( n20055 ) == ( bv_1_0_n53 )  ;
assign n20057 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n20058 =  ( n20056 ) & (n20057 )  ;
assign n20059 =  ( n20058 ) & (wr )  ;
assign n20060 =  ( n20059 ) ? ( n5096 ) : ( iram_152 ) ;
assign n20061 = wr_addr[7:7] ;
assign n20062 =  ( n20061 ) == ( bv_1_0_n53 )  ;
assign n20063 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n20064 =  ( n20062 ) & (n20063 )  ;
assign n20065 =  ( n20064 ) & (wr )  ;
assign n20066 =  ( n20065 ) ? ( n5123 ) : ( iram_152 ) ;
assign n20067 = wr_addr[7:7] ;
assign n20068 =  ( n20067 ) == ( bv_1_0_n53 )  ;
assign n20069 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n20070 =  ( n20068 ) & (n20069 )  ;
assign n20071 =  ( n20070 ) & (wr )  ;
assign n20072 =  ( n20071 ) ? ( n5165 ) : ( iram_152 ) ;
assign n20073 = wr_addr[7:7] ;
assign n20074 =  ( n20073 ) == ( bv_1_0_n53 )  ;
assign n20075 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n20076 =  ( n20074 ) & (n20075 )  ;
assign n20077 =  ( n20076 ) & (wr )  ;
assign n20078 =  ( n20077 ) ? ( n5204 ) : ( iram_152 ) ;
assign n20079 = wr_addr[7:7] ;
assign n20080 =  ( n20079 ) == ( bv_1_0_n53 )  ;
assign n20081 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n20082 =  ( n20080 ) & (n20081 )  ;
assign n20083 =  ( n20082 ) & (wr )  ;
assign n20084 =  ( n20083 ) ? ( n5262 ) : ( iram_152 ) ;
assign n20085 = wr_addr[7:7] ;
assign n20086 =  ( n20085 ) == ( bv_1_0_n53 )  ;
assign n20087 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n20088 =  ( n20086 ) & (n20087 )  ;
assign n20089 =  ( n20088 ) & (wr )  ;
assign n20090 =  ( n20089 ) ? ( n5298 ) : ( iram_152 ) ;
assign n20091 = wr_addr[7:7] ;
assign n20092 =  ( n20091 ) == ( bv_1_0_n53 )  ;
assign n20093 =  ( wr_addr ) == ( bv_8_152_n373 )  ;
assign n20094 =  ( n20092 ) & (n20093 )  ;
assign n20095 =  ( n20094 ) & (wr )  ;
assign n20096 =  ( n20095 ) ? ( n5325 ) : ( iram_152 ) ;
assign n20097 = wr_addr[7:7] ;
assign n20098 =  ( n20097 ) == ( bv_1_0_n53 )  ;
assign n20099 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n20100 =  ( n20098 ) & (n20099 )  ;
assign n20101 =  ( n20100 ) & (wr )  ;
assign n20102 =  ( n20101 ) ? ( n4782 ) : ( iram_153 ) ;
assign n20103 = wr_addr[7:7] ;
assign n20104 =  ( n20103 ) == ( bv_1_0_n53 )  ;
assign n20105 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n20106 =  ( n20104 ) & (n20105 )  ;
assign n20107 =  ( n20106 ) & (wr )  ;
assign n20108 =  ( n20107 ) ? ( n4841 ) : ( iram_153 ) ;
assign n20109 = wr_addr[7:7] ;
assign n20110 =  ( n20109 ) == ( bv_1_0_n53 )  ;
assign n20111 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n20112 =  ( n20110 ) & (n20111 )  ;
assign n20113 =  ( n20112 ) & (wr )  ;
assign n20114 =  ( n20113 ) ? ( n5449 ) : ( iram_153 ) ;
assign n20115 = wr_addr[7:7] ;
assign n20116 =  ( n20115 ) == ( bv_1_0_n53 )  ;
assign n20117 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n20118 =  ( n20116 ) & (n20117 )  ;
assign n20119 =  ( n20118 ) & (wr )  ;
assign n20120 =  ( n20119 ) ? ( n4906 ) : ( iram_153 ) ;
assign n20121 = wr_addr[7:7] ;
assign n20122 =  ( n20121 ) == ( bv_1_0_n53 )  ;
assign n20123 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n20124 =  ( n20122 ) & (n20123 )  ;
assign n20125 =  ( n20124 ) & (wr )  ;
assign n20126 =  ( n20125 ) ? ( n5485 ) : ( iram_153 ) ;
assign n20127 = wr_addr[7:7] ;
assign n20128 =  ( n20127 ) == ( bv_1_0_n53 )  ;
assign n20129 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n20130 =  ( n20128 ) & (n20129 )  ;
assign n20131 =  ( n20130 ) & (wr )  ;
assign n20132 =  ( n20131 ) ? ( n5512 ) : ( iram_153 ) ;
assign n20133 = wr_addr[7:7] ;
assign n20134 =  ( n20133 ) == ( bv_1_0_n53 )  ;
assign n20135 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n20136 =  ( n20134 ) & (n20135 )  ;
assign n20137 =  ( n20136 ) & (wr )  ;
assign n20138 =  ( n20137 ) ? ( bv_8_0_n69 ) : ( iram_153 ) ;
assign n20139 = wr_addr[7:7] ;
assign n20140 =  ( n20139 ) == ( bv_1_0_n53 )  ;
assign n20141 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n20142 =  ( n20140 ) & (n20141 )  ;
assign n20143 =  ( n20142 ) & (wr )  ;
assign n20144 =  ( n20143 ) ? ( n5071 ) : ( iram_153 ) ;
assign n20145 = wr_addr[7:7] ;
assign n20146 =  ( n20145 ) == ( bv_1_0_n53 )  ;
assign n20147 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n20148 =  ( n20146 ) & (n20147 )  ;
assign n20149 =  ( n20148 ) & (wr )  ;
assign n20150 =  ( n20149 ) ? ( n5096 ) : ( iram_153 ) ;
assign n20151 = wr_addr[7:7] ;
assign n20152 =  ( n20151 ) == ( bv_1_0_n53 )  ;
assign n20153 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n20154 =  ( n20152 ) & (n20153 )  ;
assign n20155 =  ( n20154 ) & (wr )  ;
assign n20156 =  ( n20155 ) ? ( n5123 ) : ( iram_153 ) ;
assign n20157 = wr_addr[7:7] ;
assign n20158 =  ( n20157 ) == ( bv_1_0_n53 )  ;
assign n20159 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n20160 =  ( n20158 ) & (n20159 )  ;
assign n20161 =  ( n20160 ) & (wr )  ;
assign n20162 =  ( n20161 ) ? ( n5165 ) : ( iram_153 ) ;
assign n20163 = wr_addr[7:7] ;
assign n20164 =  ( n20163 ) == ( bv_1_0_n53 )  ;
assign n20165 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n20166 =  ( n20164 ) & (n20165 )  ;
assign n20167 =  ( n20166 ) & (wr )  ;
assign n20168 =  ( n20167 ) ? ( n5204 ) : ( iram_153 ) ;
assign n20169 = wr_addr[7:7] ;
assign n20170 =  ( n20169 ) == ( bv_1_0_n53 )  ;
assign n20171 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n20172 =  ( n20170 ) & (n20171 )  ;
assign n20173 =  ( n20172 ) & (wr )  ;
assign n20174 =  ( n20173 ) ? ( n5262 ) : ( iram_153 ) ;
assign n20175 = wr_addr[7:7] ;
assign n20176 =  ( n20175 ) == ( bv_1_0_n53 )  ;
assign n20177 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n20178 =  ( n20176 ) & (n20177 )  ;
assign n20179 =  ( n20178 ) & (wr )  ;
assign n20180 =  ( n20179 ) ? ( n5298 ) : ( iram_153 ) ;
assign n20181 = wr_addr[7:7] ;
assign n20182 =  ( n20181 ) == ( bv_1_0_n53 )  ;
assign n20183 =  ( wr_addr ) == ( bv_8_153_n375 )  ;
assign n20184 =  ( n20182 ) & (n20183 )  ;
assign n20185 =  ( n20184 ) & (wr )  ;
assign n20186 =  ( n20185 ) ? ( n5325 ) : ( iram_153 ) ;
assign n20187 = wr_addr[7:7] ;
assign n20188 =  ( n20187 ) == ( bv_1_0_n53 )  ;
assign n20189 =  ( wr_addr ) == ( bv_8_154_n377 )  ;
assign n20190 =  ( n20188 ) & (n20189 )  ;
assign n20191 =  ( n20190 ) & (wr )  ;
assign n20192 =  ( n20191 ) ? ( n4782 ) : ( iram_154 ) ;
assign n20193 = wr_addr[7:7] ;
assign n20194 =  ( n20193 ) == ( bv_1_0_n53 )  ;
assign n20195 =  ( wr_addr ) == ( bv_8_154_n377 )  ;
assign n20196 =  ( n20194 ) & (n20195 )  ;
assign n20197 =  ( n20196 ) & (wr )  ;
assign n20198 =  ( n20197 ) ? ( n4841 ) : ( iram_154 ) ;
assign n20199 = wr_addr[7:7] ;
assign n20200 =  ( n20199 ) == ( bv_1_0_n53 )  ;
assign n20201 =  ( wr_addr ) == ( bv_8_154_n377 )  ;
assign n20202 =  ( n20200 ) & (n20201 )  ;
assign n20203 =  ( n20202 ) & (wr )  ;
assign n20204 =  ( n20203 ) ? ( n5449 ) : ( iram_154 ) ;
assign n20205 = wr_addr[7:7] ;
assign n20206 =  ( n20205 ) == ( bv_1_0_n53 )  ;
assign n20207 =  ( wr_addr ) == ( bv_8_154_n377 )  ;
assign n20208 =  ( n20206 ) & (n20207 )  ;
assign n20209 =  ( n20208 ) & (wr )  ;
assign n20210 =  ( n20209 ) ? ( n4906 ) : ( iram_154 ) ;
assign n20211 = wr_addr[7:7] ;
assign n20212 =  ( n20211 ) == ( bv_1_0_n53 )  ;
assign n20213 =  ( wr_addr ) == ( bv_8_154_n377 )  ;
assign n20214 =  ( n20212 ) & (n20213 )  ;
assign n20215 =  ( n20214 ) & (wr )  ;
assign n20216 =  ( n20215 ) ? ( n5485 ) : ( iram_154 ) ;
assign n20217 = wr_addr[7:7] ;
assign n20218 =  ( n20217 ) == ( bv_1_0_n53 )  ;
assign n20219 =  ( wr_addr ) == ( bv_8_154_n377 )  ;
assign n20220 =  ( n20218 ) & (n20219 )  ;
assign n20221 =  ( n20220 ) & (wr )  ;
assign n20222 =  ( n20221 ) ? ( n5512 ) : ( iram_154 ) ;
assign n20223 = wr_addr[7:7] ;
assign n20224 =  ( n20223 ) == ( bv_1_0_n53 )  ;
assign n20225 =  ( wr_addr ) == ( bv_8_154_n377 )  ;
assign n20226 =  ( n20224 ) & (n20225 )  ;
assign n20227 =  ( n20226 ) & (wr )  ;
assign n20228 =  ( n20227 ) ? ( bv_8_0_n69 ) : ( iram_154 ) ;
assign n20229 = wr_addr[7:7] ;
assign n20230 =  ( n20229 ) == ( bv_1_0_n53 )  ;
assign n20231 =  ( wr_addr ) == ( bv_8_154_n377 )  ;
assign n20232 =  ( n20230 ) & (n20231 )  ;
assign n20233 =  ( n20232 ) & (wr )  ;
assign n20234 =  ( n20233 ) ? ( n5071 ) : ( iram_154 ) ;
assign n20235 = wr_addr[7:7] ;
assign n20236 =  ( n20235 ) == ( bv_1_0_n53 )  ;
assign n20237 =  ( wr_addr ) == ( bv_8_154_n377 )  ;
assign n20238 =  ( n20236 ) & (n20237 )  ;
assign n20239 =  ( n20238 ) & (wr )  ;
assign n20240 =  ( n20239 ) ? ( n5096 ) : ( iram_154 ) ;
assign n20241 = wr_addr[7:7] ;
assign n20242 =  ( n20241 ) == ( bv_1_0_n53 )  ;
assign n20243 =  ( wr_addr ) == ( bv_8_154_n377 )  ;
assign n20244 =  ( n20242 ) & (n20243 )  ;
assign n20245 =  ( n20244 ) & (wr )  ;
assign n20246 =  ( n20245 ) ? ( n5123 ) : ( iram_154 ) ;
assign n20247 = wr_addr[7:7] ;
assign n20248 =  ( n20247 ) == ( bv_1_0_n53 )  ;
assign n20249 =  ( wr_addr ) == ( bv_8_154_n377 )  ;
assign n20250 =  ( n20248 ) & (n20249 )  ;
assign n20251 =  ( n20250 ) & (wr )  ;
assign n20252 =  ( n20251 ) ? ( n5165 ) : ( iram_154 ) ;
assign n20253 = wr_addr[7:7] ;
assign n20254 =  ( n20253 ) == ( bv_1_0_n53 )  ;
assign n20255 =  ( wr_addr ) == ( bv_8_154_n377 )  ;
assign n20256 =  ( n20254 ) & (n20255 )  ;
assign n20257 =  ( n20256 ) & (wr )  ;
assign n20258 =  ( n20257 ) ? ( n5204 ) : ( iram_154 ) ;
assign n20259 = wr_addr[7:7] ;
assign n20260 =  ( n20259 ) == ( bv_1_0_n53 )  ;
assign n20261 =  ( wr_addr ) == ( bv_8_154_n377 )  ;
assign n20262 =  ( n20260 ) & (n20261 )  ;
assign n20263 =  ( n20262 ) & (wr )  ;
assign n20264 =  ( n20263 ) ? ( n5262 ) : ( iram_154 ) ;
assign n20265 = wr_addr[7:7] ;
assign n20266 =  ( n20265 ) == ( bv_1_0_n53 )  ;
assign n20267 =  ( wr_addr ) == ( bv_8_154_n377 )  ;
assign n20268 =  ( n20266 ) & (n20267 )  ;
assign n20269 =  ( n20268 ) & (wr )  ;
assign n20270 =  ( n20269 ) ? ( n5298 ) : ( iram_154 ) ;
assign n20271 = wr_addr[7:7] ;
assign n20272 =  ( n20271 ) == ( bv_1_0_n53 )  ;
assign n20273 =  ( wr_addr ) == ( bv_8_154_n377 )  ;
assign n20274 =  ( n20272 ) & (n20273 )  ;
assign n20275 =  ( n20274 ) & (wr )  ;
assign n20276 =  ( n20275 ) ? ( n5325 ) : ( iram_154 ) ;
assign n20277 = wr_addr[7:7] ;
assign n20278 =  ( n20277 ) == ( bv_1_0_n53 )  ;
assign n20279 =  ( wr_addr ) == ( bv_8_155_n379 )  ;
assign n20280 =  ( n20278 ) & (n20279 )  ;
assign n20281 =  ( n20280 ) & (wr )  ;
assign n20282 =  ( n20281 ) ? ( n4782 ) : ( iram_155 ) ;
assign n20283 = wr_addr[7:7] ;
assign n20284 =  ( n20283 ) == ( bv_1_0_n53 )  ;
assign n20285 =  ( wr_addr ) == ( bv_8_155_n379 )  ;
assign n20286 =  ( n20284 ) & (n20285 )  ;
assign n20287 =  ( n20286 ) & (wr )  ;
assign n20288 =  ( n20287 ) ? ( n4841 ) : ( iram_155 ) ;
assign n20289 = wr_addr[7:7] ;
assign n20290 =  ( n20289 ) == ( bv_1_0_n53 )  ;
assign n20291 =  ( wr_addr ) == ( bv_8_155_n379 )  ;
assign n20292 =  ( n20290 ) & (n20291 )  ;
assign n20293 =  ( n20292 ) & (wr )  ;
assign n20294 =  ( n20293 ) ? ( n5449 ) : ( iram_155 ) ;
assign n20295 = wr_addr[7:7] ;
assign n20296 =  ( n20295 ) == ( bv_1_0_n53 )  ;
assign n20297 =  ( wr_addr ) == ( bv_8_155_n379 )  ;
assign n20298 =  ( n20296 ) & (n20297 )  ;
assign n20299 =  ( n20298 ) & (wr )  ;
assign n20300 =  ( n20299 ) ? ( n4906 ) : ( iram_155 ) ;
assign n20301 = wr_addr[7:7] ;
assign n20302 =  ( n20301 ) == ( bv_1_0_n53 )  ;
assign n20303 =  ( wr_addr ) == ( bv_8_155_n379 )  ;
assign n20304 =  ( n20302 ) & (n20303 )  ;
assign n20305 =  ( n20304 ) & (wr )  ;
assign n20306 =  ( n20305 ) ? ( n5485 ) : ( iram_155 ) ;
assign n20307 = wr_addr[7:7] ;
assign n20308 =  ( n20307 ) == ( bv_1_0_n53 )  ;
assign n20309 =  ( wr_addr ) == ( bv_8_155_n379 )  ;
assign n20310 =  ( n20308 ) & (n20309 )  ;
assign n20311 =  ( n20310 ) & (wr )  ;
assign n20312 =  ( n20311 ) ? ( n5512 ) : ( iram_155 ) ;
assign n20313 = wr_addr[7:7] ;
assign n20314 =  ( n20313 ) == ( bv_1_0_n53 )  ;
assign n20315 =  ( wr_addr ) == ( bv_8_155_n379 )  ;
assign n20316 =  ( n20314 ) & (n20315 )  ;
assign n20317 =  ( n20316 ) & (wr )  ;
assign n20318 =  ( n20317 ) ? ( bv_8_0_n69 ) : ( iram_155 ) ;
assign n20319 = wr_addr[7:7] ;
assign n20320 =  ( n20319 ) == ( bv_1_0_n53 )  ;
assign n20321 =  ( wr_addr ) == ( bv_8_155_n379 )  ;
assign n20322 =  ( n20320 ) & (n20321 )  ;
assign n20323 =  ( n20322 ) & (wr )  ;
assign n20324 =  ( n20323 ) ? ( n5071 ) : ( iram_155 ) ;
assign n20325 = wr_addr[7:7] ;
assign n20326 =  ( n20325 ) == ( bv_1_0_n53 )  ;
assign n20327 =  ( wr_addr ) == ( bv_8_155_n379 )  ;
assign n20328 =  ( n20326 ) & (n20327 )  ;
assign n20329 =  ( n20328 ) & (wr )  ;
assign n20330 =  ( n20329 ) ? ( n5096 ) : ( iram_155 ) ;
assign n20331 = wr_addr[7:7] ;
assign n20332 =  ( n20331 ) == ( bv_1_0_n53 )  ;
assign n20333 =  ( wr_addr ) == ( bv_8_155_n379 )  ;
assign n20334 =  ( n20332 ) & (n20333 )  ;
assign n20335 =  ( n20334 ) & (wr )  ;
assign n20336 =  ( n20335 ) ? ( n5123 ) : ( iram_155 ) ;
assign n20337 = wr_addr[7:7] ;
assign n20338 =  ( n20337 ) == ( bv_1_0_n53 )  ;
assign n20339 =  ( wr_addr ) == ( bv_8_155_n379 )  ;
assign n20340 =  ( n20338 ) & (n20339 )  ;
assign n20341 =  ( n20340 ) & (wr )  ;
assign n20342 =  ( n20341 ) ? ( n5165 ) : ( iram_155 ) ;
assign n20343 = wr_addr[7:7] ;
assign n20344 =  ( n20343 ) == ( bv_1_0_n53 )  ;
assign n20345 =  ( wr_addr ) == ( bv_8_155_n379 )  ;
assign n20346 =  ( n20344 ) & (n20345 )  ;
assign n20347 =  ( n20346 ) & (wr )  ;
assign n20348 =  ( n20347 ) ? ( n5204 ) : ( iram_155 ) ;
assign n20349 = wr_addr[7:7] ;
assign n20350 =  ( n20349 ) == ( bv_1_0_n53 )  ;
assign n20351 =  ( wr_addr ) == ( bv_8_155_n379 )  ;
assign n20352 =  ( n20350 ) & (n20351 )  ;
assign n20353 =  ( n20352 ) & (wr )  ;
assign n20354 =  ( n20353 ) ? ( n5262 ) : ( iram_155 ) ;
assign n20355 = wr_addr[7:7] ;
assign n20356 =  ( n20355 ) == ( bv_1_0_n53 )  ;
assign n20357 =  ( wr_addr ) == ( bv_8_155_n379 )  ;
assign n20358 =  ( n20356 ) & (n20357 )  ;
assign n20359 =  ( n20358 ) & (wr )  ;
assign n20360 =  ( n20359 ) ? ( n5298 ) : ( iram_155 ) ;
assign n20361 = wr_addr[7:7] ;
assign n20362 =  ( n20361 ) == ( bv_1_0_n53 )  ;
assign n20363 =  ( wr_addr ) == ( bv_8_155_n379 )  ;
assign n20364 =  ( n20362 ) & (n20363 )  ;
assign n20365 =  ( n20364 ) & (wr )  ;
assign n20366 =  ( n20365 ) ? ( n5325 ) : ( iram_155 ) ;
assign n20367 = wr_addr[7:7] ;
assign n20368 =  ( n20367 ) == ( bv_1_0_n53 )  ;
assign n20369 =  ( wr_addr ) == ( bv_8_156_n381 )  ;
assign n20370 =  ( n20368 ) & (n20369 )  ;
assign n20371 =  ( n20370 ) & (wr )  ;
assign n20372 =  ( n20371 ) ? ( n4782 ) : ( iram_156 ) ;
assign n20373 = wr_addr[7:7] ;
assign n20374 =  ( n20373 ) == ( bv_1_0_n53 )  ;
assign n20375 =  ( wr_addr ) == ( bv_8_156_n381 )  ;
assign n20376 =  ( n20374 ) & (n20375 )  ;
assign n20377 =  ( n20376 ) & (wr )  ;
assign n20378 =  ( n20377 ) ? ( n4841 ) : ( iram_156 ) ;
assign n20379 = wr_addr[7:7] ;
assign n20380 =  ( n20379 ) == ( bv_1_0_n53 )  ;
assign n20381 =  ( wr_addr ) == ( bv_8_156_n381 )  ;
assign n20382 =  ( n20380 ) & (n20381 )  ;
assign n20383 =  ( n20382 ) & (wr )  ;
assign n20384 =  ( n20383 ) ? ( n5449 ) : ( iram_156 ) ;
assign n20385 = wr_addr[7:7] ;
assign n20386 =  ( n20385 ) == ( bv_1_0_n53 )  ;
assign n20387 =  ( wr_addr ) == ( bv_8_156_n381 )  ;
assign n20388 =  ( n20386 ) & (n20387 )  ;
assign n20389 =  ( n20388 ) & (wr )  ;
assign n20390 =  ( n20389 ) ? ( n4906 ) : ( iram_156 ) ;
assign n20391 = wr_addr[7:7] ;
assign n20392 =  ( n20391 ) == ( bv_1_0_n53 )  ;
assign n20393 =  ( wr_addr ) == ( bv_8_156_n381 )  ;
assign n20394 =  ( n20392 ) & (n20393 )  ;
assign n20395 =  ( n20394 ) & (wr )  ;
assign n20396 =  ( n20395 ) ? ( n5485 ) : ( iram_156 ) ;
assign n20397 = wr_addr[7:7] ;
assign n20398 =  ( n20397 ) == ( bv_1_0_n53 )  ;
assign n20399 =  ( wr_addr ) == ( bv_8_156_n381 )  ;
assign n20400 =  ( n20398 ) & (n20399 )  ;
assign n20401 =  ( n20400 ) & (wr )  ;
assign n20402 =  ( n20401 ) ? ( n5512 ) : ( iram_156 ) ;
assign n20403 = wr_addr[7:7] ;
assign n20404 =  ( n20403 ) == ( bv_1_0_n53 )  ;
assign n20405 =  ( wr_addr ) == ( bv_8_156_n381 )  ;
assign n20406 =  ( n20404 ) & (n20405 )  ;
assign n20407 =  ( n20406 ) & (wr )  ;
assign n20408 =  ( n20407 ) ? ( bv_8_0_n69 ) : ( iram_156 ) ;
assign n20409 = wr_addr[7:7] ;
assign n20410 =  ( n20409 ) == ( bv_1_0_n53 )  ;
assign n20411 =  ( wr_addr ) == ( bv_8_156_n381 )  ;
assign n20412 =  ( n20410 ) & (n20411 )  ;
assign n20413 =  ( n20412 ) & (wr )  ;
assign n20414 =  ( n20413 ) ? ( n5071 ) : ( iram_156 ) ;
assign n20415 = wr_addr[7:7] ;
assign n20416 =  ( n20415 ) == ( bv_1_0_n53 )  ;
assign n20417 =  ( wr_addr ) == ( bv_8_156_n381 )  ;
assign n20418 =  ( n20416 ) & (n20417 )  ;
assign n20419 =  ( n20418 ) & (wr )  ;
assign n20420 =  ( n20419 ) ? ( n5096 ) : ( iram_156 ) ;
assign n20421 = wr_addr[7:7] ;
assign n20422 =  ( n20421 ) == ( bv_1_0_n53 )  ;
assign n20423 =  ( wr_addr ) == ( bv_8_156_n381 )  ;
assign n20424 =  ( n20422 ) & (n20423 )  ;
assign n20425 =  ( n20424 ) & (wr )  ;
assign n20426 =  ( n20425 ) ? ( n5123 ) : ( iram_156 ) ;
assign n20427 = wr_addr[7:7] ;
assign n20428 =  ( n20427 ) == ( bv_1_0_n53 )  ;
assign n20429 =  ( wr_addr ) == ( bv_8_156_n381 )  ;
assign n20430 =  ( n20428 ) & (n20429 )  ;
assign n20431 =  ( n20430 ) & (wr )  ;
assign n20432 =  ( n20431 ) ? ( n5165 ) : ( iram_156 ) ;
assign n20433 = wr_addr[7:7] ;
assign n20434 =  ( n20433 ) == ( bv_1_0_n53 )  ;
assign n20435 =  ( wr_addr ) == ( bv_8_156_n381 )  ;
assign n20436 =  ( n20434 ) & (n20435 )  ;
assign n20437 =  ( n20436 ) & (wr )  ;
assign n20438 =  ( n20437 ) ? ( n5204 ) : ( iram_156 ) ;
assign n20439 = wr_addr[7:7] ;
assign n20440 =  ( n20439 ) == ( bv_1_0_n53 )  ;
assign n20441 =  ( wr_addr ) == ( bv_8_156_n381 )  ;
assign n20442 =  ( n20440 ) & (n20441 )  ;
assign n20443 =  ( n20442 ) & (wr )  ;
assign n20444 =  ( n20443 ) ? ( n5262 ) : ( iram_156 ) ;
assign n20445 = wr_addr[7:7] ;
assign n20446 =  ( n20445 ) == ( bv_1_0_n53 )  ;
assign n20447 =  ( wr_addr ) == ( bv_8_156_n381 )  ;
assign n20448 =  ( n20446 ) & (n20447 )  ;
assign n20449 =  ( n20448 ) & (wr )  ;
assign n20450 =  ( n20449 ) ? ( n5298 ) : ( iram_156 ) ;
assign n20451 = wr_addr[7:7] ;
assign n20452 =  ( n20451 ) == ( bv_1_0_n53 )  ;
assign n20453 =  ( wr_addr ) == ( bv_8_156_n381 )  ;
assign n20454 =  ( n20452 ) & (n20453 )  ;
assign n20455 =  ( n20454 ) & (wr )  ;
assign n20456 =  ( n20455 ) ? ( n5325 ) : ( iram_156 ) ;
assign n20457 = wr_addr[7:7] ;
assign n20458 =  ( n20457 ) == ( bv_1_0_n53 )  ;
assign n20459 =  ( wr_addr ) == ( bv_8_157_n383 )  ;
assign n20460 =  ( n20458 ) & (n20459 )  ;
assign n20461 =  ( n20460 ) & (wr )  ;
assign n20462 =  ( n20461 ) ? ( n4782 ) : ( iram_157 ) ;
assign n20463 = wr_addr[7:7] ;
assign n20464 =  ( n20463 ) == ( bv_1_0_n53 )  ;
assign n20465 =  ( wr_addr ) == ( bv_8_157_n383 )  ;
assign n20466 =  ( n20464 ) & (n20465 )  ;
assign n20467 =  ( n20466 ) & (wr )  ;
assign n20468 =  ( n20467 ) ? ( n4841 ) : ( iram_157 ) ;
assign n20469 = wr_addr[7:7] ;
assign n20470 =  ( n20469 ) == ( bv_1_0_n53 )  ;
assign n20471 =  ( wr_addr ) == ( bv_8_157_n383 )  ;
assign n20472 =  ( n20470 ) & (n20471 )  ;
assign n20473 =  ( n20472 ) & (wr )  ;
assign n20474 =  ( n20473 ) ? ( n5449 ) : ( iram_157 ) ;
assign n20475 = wr_addr[7:7] ;
assign n20476 =  ( n20475 ) == ( bv_1_0_n53 )  ;
assign n20477 =  ( wr_addr ) == ( bv_8_157_n383 )  ;
assign n20478 =  ( n20476 ) & (n20477 )  ;
assign n20479 =  ( n20478 ) & (wr )  ;
assign n20480 =  ( n20479 ) ? ( n4906 ) : ( iram_157 ) ;
assign n20481 = wr_addr[7:7] ;
assign n20482 =  ( n20481 ) == ( bv_1_0_n53 )  ;
assign n20483 =  ( wr_addr ) == ( bv_8_157_n383 )  ;
assign n20484 =  ( n20482 ) & (n20483 )  ;
assign n20485 =  ( n20484 ) & (wr )  ;
assign n20486 =  ( n20485 ) ? ( n5485 ) : ( iram_157 ) ;
assign n20487 = wr_addr[7:7] ;
assign n20488 =  ( n20487 ) == ( bv_1_0_n53 )  ;
assign n20489 =  ( wr_addr ) == ( bv_8_157_n383 )  ;
assign n20490 =  ( n20488 ) & (n20489 )  ;
assign n20491 =  ( n20490 ) & (wr )  ;
assign n20492 =  ( n20491 ) ? ( n5512 ) : ( iram_157 ) ;
assign n20493 = wr_addr[7:7] ;
assign n20494 =  ( n20493 ) == ( bv_1_0_n53 )  ;
assign n20495 =  ( wr_addr ) == ( bv_8_157_n383 )  ;
assign n20496 =  ( n20494 ) & (n20495 )  ;
assign n20497 =  ( n20496 ) & (wr )  ;
assign n20498 =  ( n20497 ) ? ( bv_8_0_n69 ) : ( iram_157 ) ;
assign n20499 = wr_addr[7:7] ;
assign n20500 =  ( n20499 ) == ( bv_1_0_n53 )  ;
assign n20501 =  ( wr_addr ) == ( bv_8_157_n383 )  ;
assign n20502 =  ( n20500 ) & (n20501 )  ;
assign n20503 =  ( n20502 ) & (wr )  ;
assign n20504 =  ( n20503 ) ? ( n5071 ) : ( iram_157 ) ;
assign n20505 = wr_addr[7:7] ;
assign n20506 =  ( n20505 ) == ( bv_1_0_n53 )  ;
assign n20507 =  ( wr_addr ) == ( bv_8_157_n383 )  ;
assign n20508 =  ( n20506 ) & (n20507 )  ;
assign n20509 =  ( n20508 ) & (wr )  ;
assign n20510 =  ( n20509 ) ? ( n5096 ) : ( iram_157 ) ;
assign n20511 = wr_addr[7:7] ;
assign n20512 =  ( n20511 ) == ( bv_1_0_n53 )  ;
assign n20513 =  ( wr_addr ) == ( bv_8_157_n383 )  ;
assign n20514 =  ( n20512 ) & (n20513 )  ;
assign n20515 =  ( n20514 ) & (wr )  ;
assign n20516 =  ( n20515 ) ? ( n5123 ) : ( iram_157 ) ;
assign n20517 = wr_addr[7:7] ;
assign n20518 =  ( n20517 ) == ( bv_1_0_n53 )  ;
assign n20519 =  ( wr_addr ) == ( bv_8_157_n383 )  ;
assign n20520 =  ( n20518 ) & (n20519 )  ;
assign n20521 =  ( n20520 ) & (wr )  ;
assign n20522 =  ( n20521 ) ? ( n5165 ) : ( iram_157 ) ;
assign n20523 = wr_addr[7:7] ;
assign n20524 =  ( n20523 ) == ( bv_1_0_n53 )  ;
assign n20525 =  ( wr_addr ) == ( bv_8_157_n383 )  ;
assign n20526 =  ( n20524 ) & (n20525 )  ;
assign n20527 =  ( n20526 ) & (wr )  ;
assign n20528 =  ( n20527 ) ? ( n5204 ) : ( iram_157 ) ;
assign n20529 = wr_addr[7:7] ;
assign n20530 =  ( n20529 ) == ( bv_1_0_n53 )  ;
assign n20531 =  ( wr_addr ) == ( bv_8_157_n383 )  ;
assign n20532 =  ( n20530 ) & (n20531 )  ;
assign n20533 =  ( n20532 ) & (wr )  ;
assign n20534 =  ( n20533 ) ? ( n5262 ) : ( iram_157 ) ;
assign n20535 = wr_addr[7:7] ;
assign n20536 =  ( n20535 ) == ( bv_1_0_n53 )  ;
assign n20537 =  ( wr_addr ) == ( bv_8_157_n383 )  ;
assign n20538 =  ( n20536 ) & (n20537 )  ;
assign n20539 =  ( n20538 ) & (wr )  ;
assign n20540 =  ( n20539 ) ? ( n5298 ) : ( iram_157 ) ;
assign n20541 = wr_addr[7:7] ;
assign n20542 =  ( n20541 ) == ( bv_1_0_n53 )  ;
assign n20543 =  ( wr_addr ) == ( bv_8_157_n383 )  ;
assign n20544 =  ( n20542 ) & (n20543 )  ;
assign n20545 =  ( n20544 ) & (wr )  ;
assign n20546 =  ( n20545 ) ? ( n5325 ) : ( iram_157 ) ;
assign n20547 = wr_addr[7:7] ;
assign n20548 =  ( n20547 ) == ( bv_1_0_n53 )  ;
assign n20549 =  ( wr_addr ) == ( bv_8_158_n385 )  ;
assign n20550 =  ( n20548 ) & (n20549 )  ;
assign n20551 =  ( n20550 ) & (wr )  ;
assign n20552 =  ( n20551 ) ? ( n4782 ) : ( iram_158 ) ;
assign n20553 = wr_addr[7:7] ;
assign n20554 =  ( n20553 ) == ( bv_1_0_n53 )  ;
assign n20555 =  ( wr_addr ) == ( bv_8_158_n385 )  ;
assign n20556 =  ( n20554 ) & (n20555 )  ;
assign n20557 =  ( n20556 ) & (wr )  ;
assign n20558 =  ( n20557 ) ? ( n4841 ) : ( iram_158 ) ;
assign n20559 = wr_addr[7:7] ;
assign n20560 =  ( n20559 ) == ( bv_1_0_n53 )  ;
assign n20561 =  ( wr_addr ) == ( bv_8_158_n385 )  ;
assign n20562 =  ( n20560 ) & (n20561 )  ;
assign n20563 =  ( n20562 ) & (wr )  ;
assign n20564 =  ( n20563 ) ? ( n5449 ) : ( iram_158 ) ;
assign n20565 = wr_addr[7:7] ;
assign n20566 =  ( n20565 ) == ( bv_1_0_n53 )  ;
assign n20567 =  ( wr_addr ) == ( bv_8_158_n385 )  ;
assign n20568 =  ( n20566 ) & (n20567 )  ;
assign n20569 =  ( n20568 ) & (wr )  ;
assign n20570 =  ( n20569 ) ? ( n4906 ) : ( iram_158 ) ;
assign n20571 = wr_addr[7:7] ;
assign n20572 =  ( n20571 ) == ( bv_1_0_n53 )  ;
assign n20573 =  ( wr_addr ) == ( bv_8_158_n385 )  ;
assign n20574 =  ( n20572 ) & (n20573 )  ;
assign n20575 =  ( n20574 ) & (wr )  ;
assign n20576 =  ( n20575 ) ? ( n5485 ) : ( iram_158 ) ;
assign n20577 = wr_addr[7:7] ;
assign n20578 =  ( n20577 ) == ( bv_1_0_n53 )  ;
assign n20579 =  ( wr_addr ) == ( bv_8_158_n385 )  ;
assign n20580 =  ( n20578 ) & (n20579 )  ;
assign n20581 =  ( n20580 ) & (wr )  ;
assign n20582 =  ( n20581 ) ? ( n5512 ) : ( iram_158 ) ;
assign n20583 = wr_addr[7:7] ;
assign n20584 =  ( n20583 ) == ( bv_1_0_n53 )  ;
assign n20585 =  ( wr_addr ) == ( bv_8_158_n385 )  ;
assign n20586 =  ( n20584 ) & (n20585 )  ;
assign n20587 =  ( n20586 ) & (wr )  ;
assign n20588 =  ( n20587 ) ? ( bv_8_0_n69 ) : ( iram_158 ) ;
assign n20589 = wr_addr[7:7] ;
assign n20590 =  ( n20589 ) == ( bv_1_0_n53 )  ;
assign n20591 =  ( wr_addr ) == ( bv_8_158_n385 )  ;
assign n20592 =  ( n20590 ) & (n20591 )  ;
assign n20593 =  ( n20592 ) & (wr )  ;
assign n20594 =  ( n20593 ) ? ( n5071 ) : ( iram_158 ) ;
assign n20595 = wr_addr[7:7] ;
assign n20596 =  ( n20595 ) == ( bv_1_0_n53 )  ;
assign n20597 =  ( wr_addr ) == ( bv_8_158_n385 )  ;
assign n20598 =  ( n20596 ) & (n20597 )  ;
assign n20599 =  ( n20598 ) & (wr )  ;
assign n20600 =  ( n20599 ) ? ( n5096 ) : ( iram_158 ) ;
assign n20601 = wr_addr[7:7] ;
assign n20602 =  ( n20601 ) == ( bv_1_0_n53 )  ;
assign n20603 =  ( wr_addr ) == ( bv_8_158_n385 )  ;
assign n20604 =  ( n20602 ) & (n20603 )  ;
assign n20605 =  ( n20604 ) & (wr )  ;
assign n20606 =  ( n20605 ) ? ( n5123 ) : ( iram_158 ) ;
assign n20607 = wr_addr[7:7] ;
assign n20608 =  ( n20607 ) == ( bv_1_0_n53 )  ;
assign n20609 =  ( wr_addr ) == ( bv_8_158_n385 )  ;
assign n20610 =  ( n20608 ) & (n20609 )  ;
assign n20611 =  ( n20610 ) & (wr )  ;
assign n20612 =  ( n20611 ) ? ( n5165 ) : ( iram_158 ) ;
assign n20613 = wr_addr[7:7] ;
assign n20614 =  ( n20613 ) == ( bv_1_0_n53 )  ;
assign n20615 =  ( wr_addr ) == ( bv_8_158_n385 )  ;
assign n20616 =  ( n20614 ) & (n20615 )  ;
assign n20617 =  ( n20616 ) & (wr )  ;
assign n20618 =  ( n20617 ) ? ( n5204 ) : ( iram_158 ) ;
assign n20619 = wr_addr[7:7] ;
assign n20620 =  ( n20619 ) == ( bv_1_0_n53 )  ;
assign n20621 =  ( wr_addr ) == ( bv_8_158_n385 )  ;
assign n20622 =  ( n20620 ) & (n20621 )  ;
assign n20623 =  ( n20622 ) & (wr )  ;
assign n20624 =  ( n20623 ) ? ( n5262 ) : ( iram_158 ) ;
assign n20625 = wr_addr[7:7] ;
assign n20626 =  ( n20625 ) == ( bv_1_0_n53 )  ;
assign n20627 =  ( wr_addr ) == ( bv_8_158_n385 )  ;
assign n20628 =  ( n20626 ) & (n20627 )  ;
assign n20629 =  ( n20628 ) & (wr )  ;
assign n20630 =  ( n20629 ) ? ( n5298 ) : ( iram_158 ) ;
assign n20631 = wr_addr[7:7] ;
assign n20632 =  ( n20631 ) == ( bv_1_0_n53 )  ;
assign n20633 =  ( wr_addr ) == ( bv_8_158_n385 )  ;
assign n20634 =  ( n20632 ) & (n20633 )  ;
assign n20635 =  ( n20634 ) & (wr )  ;
assign n20636 =  ( n20635 ) ? ( n5325 ) : ( iram_158 ) ;
assign n20637 = wr_addr[7:7] ;
assign n20638 =  ( n20637 ) == ( bv_1_0_n53 )  ;
assign n20639 =  ( wr_addr ) == ( bv_8_159_n387 )  ;
assign n20640 =  ( n20638 ) & (n20639 )  ;
assign n20641 =  ( n20640 ) & (wr )  ;
assign n20642 =  ( n20641 ) ? ( n4782 ) : ( iram_159 ) ;
assign n20643 = wr_addr[7:7] ;
assign n20644 =  ( n20643 ) == ( bv_1_0_n53 )  ;
assign n20645 =  ( wr_addr ) == ( bv_8_159_n387 )  ;
assign n20646 =  ( n20644 ) & (n20645 )  ;
assign n20647 =  ( n20646 ) & (wr )  ;
assign n20648 =  ( n20647 ) ? ( n4841 ) : ( iram_159 ) ;
assign n20649 = wr_addr[7:7] ;
assign n20650 =  ( n20649 ) == ( bv_1_0_n53 )  ;
assign n20651 =  ( wr_addr ) == ( bv_8_159_n387 )  ;
assign n20652 =  ( n20650 ) & (n20651 )  ;
assign n20653 =  ( n20652 ) & (wr )  ;
assign n20654 =  ( n20653 ) ? ( n5449 ) : ( iram_159 ) ;
assign n20655 = wr_addr[7:7] ;
assign n20656 =  ( n20655 ) == ( bv_1_0_n53 )  ;
assign n20657 =  ( wr_addr ) == ( bv_8_159_n387 )  ;
assign n20658 =  ( n20656 ) & (n20657 )  ;
assign n20659 =  ( n20658 ) & (wr )  ;
assign n20660 =  ( n20659 ) ? ( n4906 ) : ( iram_159 ) ;
assign n20661 = wr_addr[7:7] ;
assign n20662 =  ( n20661 ) == ( bv_1_0_n53 )  ;
assign n20663 =  ( wr_addr ) == ( bv_8_159_n387 )  ;
assign n20664 =  ( n20662 ) & (n20663 )  ;
assign n20665 =  ( n20664 ) & (wr )  ;
assign n20666 =  ( n20665 ) ? ( n5485 ) : ( iram_159 ) ;
assign n20667 = wr_addr[7:7] ;
assign n20668 =  ( n20667 ) == ( bv_1_0_n53 )  ;
assign n20669 =  ( wr_addr ) == ( bv_8_159_n387 )  ;
assign n20670 =  ( n20668 ) & (n20669 )  ;
assign n20671 =  ( n20670 ) & (wr )  ;
assign n20672 =  ( n20671 ) ? ( n5512 ) : ( iram_159 ) ;
assign n20673 = wr_addr[7:7] ;
assign n20674 =  ( n20673 ) == ( bv_1_0_n53 )  ;
assign n20675 =  ( wr_addr ) == ( bv_8_159_n387 )  ;
assign n20676 =  ( n20674 ) & (n20675 )  ;
assign n20677 =  ( n20676 ) & (wr )  ;
assign n20678 =  ( n20677 ) ? ( bv_8_0_n69 ) : ( iram_159 ) ;
assign n20679 = wr_addr[7:7] ;
assign n20680 =  ( n20679 ) == ( bv_1_0_n53 )  ;
assign n20681 =  ( wr_addr ) == ( bv_8_159_n387 )  ;
assign n20682 =  ( n20680 ) & (n20681 )  ;
assign n20683 =  ( n20682 ) & (wr )  ;
assign n20684 =  ( n20683 ) ? ( n5071 ) : ( iram_159 ) ;
assign n20685 = wr_addr[7:7] ;
assign n20686 =  ( n20685 ) == ( bv_1_0_n53 )  ;
assign n20687 =  ( wr_addr ) == ( bv_8_159_n387 )  ;
assign n20688 =  ( n20686 ) & (n20687 )  ;
assign n20689 =  ( n20688 ) & (wr )  ;
assign n20690 =  ( n20689 ) ? ( n5096 ) : ( iram_159 ) ;
assign n20691 = wr_addr[7:7] ;
assign n20692 =  ( n20691 ) == ( bv_1_0_n53 )  ;
assign n20693 =  ( wr_addr ) == ( bv_8_159_n387 )  ;
assign n20694 =  ( n20692 ) & (n20693 )  ;
assign n20695 =  ( n20694 ) & (wr )  ;
assign n20696 =  ( n20695 ) ? ( n5123 ) : ( iram_159 ) ;
assign n20697 = wr_addr[7:7] ;
assign n20698 =  ( n20697 ) == ( bv_1_0_n53 )  ;
assign n20699 =  ( wr_addr ) == ( bv_8_159_n387 )  ;
assign n20700 =  ( n20698 ) & (n20699 )  ;
assign n20701 =  ( n20700 ) & (wr )  ;
assign n20702 =  ( n20701 ) ? ( n5165 ) : ( iram_159 ) ;
assign n20703 = wr_addr[7:7] ;
assign n20704 =  ( n20703 ) == ( bv_1_0_n53 )  ;
assign n20705 =  ( wr_addr ) == ( bv_8_159_n387 )  ;
assign n20706 =  ( n20704 ) & (n20705 )  ;
assign n20707 =  ( n20706 ) & (wr )  ;
assign n20708 =  ( n20707 ) ? ( n5204 ) : ( iram_159 ) ;
assign n20709 = wr_addr[7:7] ;
assign n20710 =  ( n20709 ) == ( bv_1_0_n53 )  ;
assign n20711 =  ( wr_addr ) == ( bv_8_159_n387 )  ;
assign n20712 =  ( n20710 ) & (n20711 )  ;
assign n20713 =  ( n20712 ) & (wr )  ;
assign n20714 =  ( n20713 ) ? ( n5262 ) : ( iram_159 ) ;
assign n20715 = wr_addr[7:7] ;
assign n20716 =  ( n20715 ) == ( bv_1_0_n53 )  ;
assign n20717 =  ( wr_addr ) == ( bv_8_159_n387 )  ;
assign n20718 =  ( n20716 ) & (n20717 )  ;
assign n20719 =  ( n20718 ) & (wr )  ;
assign n20720 =  ( n20719 ) ? ( n5298 ) : ( iram_159 ) ;
assign n20721 = wr_addr[7:7] ;
assign n20722 =  ( n20721 ) == ( bv_1_0_n53 )  ;
assign n20723 =  ( wr_addr ) == ( bv_8_159_n387 )  ;
assign n20724 =  ( n20722 ) & (n20723 )  ;
assign n20725 =  ( n20724 ) & (wr )  ;
assign n20726 =  ( n20725 ) ? ( n5325 ) : ( iram_159 ) ;
assign n20727 = wr_addr[7:7] ;
assign n20728 =  ( n20727 ) == ( bv_1_0_n53 )  ;
assign n20729 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n20730 =  ( n20728 ) & (n20729 )  ;
assign n20731 =  ( n20730 ) & (wr )  ;
assign n20732 =  ( n20731 ) ? ( n4782 ) : ( iram_160 ) ;
assign n20733 = wr_addr[7:7] ;
assign n20734 =  ( n20733 ) == ( bv_1_0_n53 )  ;
assign n20735 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n20736 =  ( n20734 ) & (n20735 )  ;
assign n20737 =  ( n20736 ) & (wr )  ;
assign n20738 =  ( n20737 ) ? ( n4841 ) : ( iram_160 ) ;
assign n20739 = wr_addr[7:7] ;
assign n20740 =  ( n20739 ) == ( bv_1_0_n53 )  ;
assign n20741 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n20742 =  ( n20740 ) & (n20741 )  ;
assign n20743 =  ( n20742 ) & (wr )  ;
assign n20744 =  ( n20743 ) ? ( n5449 ) : ( iram_160 ) ;
assign n20745 = wr_addr[7:7] ;
assign n20746 =  ( n20745 ) == ( bv_1_0_n53 )  ;
assign n20747 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n20748 =  ( n20746 ) & (n20747 )  ;
assign n20749 =  ( n20748 ) & (wr )  ;
assign n20750 =  ( n20749 ) ? ( n4906 ) : ( iram_160 ) ;
assign n20751 = wr_addr[7:7] ;
assign n20752 =  ( n20751 ) == ( bv_1_0_n53 )  ;
assign n20753 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n20754 =  ( n20752 ) & (n20753 )  ;
assign n20755 =  ( n20754 ) & (wr )  ;
assign n20756 =  ( n20755 ) ? ( n5485 ) : ( iram_160 ) ;
assign n20757 = wr_addr[7:7] ;
assign n20758 =  ( n20757 ) == ( bv_1_0_n53 )  ;
assign n20759 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n20760 =  ( n20758 ) & (n20759 )  ;
assign n20761 =  ( n20760 ) & (wr )  ;
assign n20762 =  ( n20761 ) ? ( n5512 ) : ( iram_160 ) ;
assign n20763 = wr_addr[7:7] ;
assign n20764 =  ( n20763 ) == ( bv_1_0_n53 )  ;
assign n20765 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n20766 =  ( n20764 ) & (n20765 )  ;
assign n20767 =  ( n20766 ) & (wr )  ;
assign n20768 =  ( n20767 ) ? ( bv_8_0_n69 ) : ( iram_160 ) ;
assign n20769 = wr_addr[7:7] ;
assign n20770 =  ( n20769 ) == ( bv_1_0_n53 )  ;
assign n20771 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n20772 =  ( n20770 ) & (n20771 )  ;
assign n20773 =  ( n20772 ) & (wr )  ;
assign n20774 =  ( n20773 ) ? ( n5071 ) : ( iram_160 ) ;
assign n20775 = wr_addr[7:7] ;
assign n20776 =  ( n20775 ) == ( bv_1_0_n53 )  ;
assign n20777 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n20778 =  ( n20776 ) & (n20777 )  ;
assign n20779 =  ( n20778 ) & (wr )  ;
assign n20780 =  ( n20779 ) ? ( n5096 ) : ( iram_160 ) ;
assign n20781 = wr_addr[7:7] ;
assign n20782 =  ( n20781 ) == ( bv_1_0_n53 )  ;
assign n20783 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n20784 =  ( n20782 ) & (n20783 )  ;
assign n20785 =  ( n20784 ) & (wr )  ;
assign n20786 =  ( n20785 ) ? ( n5123 ) : ( iram_160 ) ;
assign n20787 = wr_addr[7:7] ;
assign n20788 =  ( n20787 ) == ( bv_1_0_n53 )  ;
assign n20789 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n20790 =  ( n20788 ) & (n20789 )  ;
assign n20791 =  ( n20790 ) & (wr )  ;
assign n20792 =  ( n20791 ) ? ( n5165 ) : ( iram_160 ) ;
assign n20793 = wr_addr[7:7] ;
assign n20794 =  ( n20793 ) == ( bv_1_0_n53 )  ;
assign n20795 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n20796 =  ( n20794 ) & (n20795 )  ;
assign n20797 =  ( n20796 ) & (wr )  ;
assign n20798 =  ( n20797 ) ? ( n5204 ) : ( iram_160 ) ;
assign n20799 = wr_addr[7:7] ;
assign n20800 =  ( n20799 ) == ( bv_1_0_n53 )  ;
assign n20801 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n20802 =  ( n20800 ) & (n20801 )  ;
assign n20803 =  ( n20802 ) & (wr )  ;
assign n20804 =  ( n20803 ) ? ( n5262 ) : ( iram_160 ) ;
assign n20805 = wr_addr[7:7] ;
assign n20806 =  ( n20805 ) == ( bv_1_0_n53 )  ;
assign n20807 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n20808 =  ( n20806 ) & (n20807 )  ;
assign n20809 =  ( n20808 ) & (wr )  ;
assign n20810 =  ( n20809 ) ? ( n5298 ) : ( iram_160 ) ;
assign n20811 = wr_addr[7:7] ;
assign n20812 =  ( n20811 ) == ( bv_1_0_n53 )  ;
assign n20813 =  ( wr_addr ) == ( bv_8_160_n389 )  ;
assign n20814 =  ( n20812 ) & (n20813 )  ;
assign n20815 =  ( n20814 ) & (wr )  ;
assign n20816 =  ( n20815 ) ? ( n5325 ) : ( iram_160 ) ;
assign n20817 = wr_addr[7:7] ;
assign n20818 =  ( n20817 ) == ( bv_1_0_n53 )  ;
assign n20819 =  ( wr_addr ) == ( bv_8_161_n391 )  ;
assign n20820 =  ( n20818 ) & (n20819 )  ;
assign n20821 =  ( n20820 ) & (wr )  ;
assign n20822 =  ( n20821 ) ? ( n4782 ) : ( iram_161 ) ;
assign n20823 = wr_addr[7:7] ;
assign n20824 =  ( n20823 ) == ( bv_1_0_n53 )  ;
assign n20825 =  ( wr_addr ) == ( bv_8_161_n391 )  ;
assign n20826 =  ( n20824 ) & (n20825 )  ;
assign n20827 =  ( n20826 ) & (wr )  ;
assign n20828 =  ( n20827 ) ? ( n4841 ) : ( iram_161 ) ;
assign n20829 = wr_addr[7:7] ;
assign n20830 =  ( n20829 ) == ( bv_1_0_n53 )  ;
assign n20831 =  ( wr_addr ) == ( bv_8_161_n391 )  ;
assign n20832 =  ( n20830 ) & (n20831 )  ;
assign n20833 =  ( n20832 ) & (wr )  ;
assign n20834 =  ( n20833 ) ? ( n5449 ) : ( iram_161 ) ;
assign n20835 = wr_addr[7:7] ;
assign n20836 =  ( n20835 ) == ( bv_1_0_n53 )  ;
assign n20837 =  ( wr_addr ) == ( bv_8_161_n391 )  ;
assign n20838 =  ( n20836 ) & (n20837 )  ;
assign n20839 =  ( n20838 ) & (wr )  ;
assign n20840 =  ( n20839 ) ? ( n4906 ) : ( iram_161 ) ;
assign n20841 = wr_addr[7:7] ;
assign n20842 =  ( n20841 ) == ( bv_1_0_n53 )  ;
assign n20843 =  ( wr_addr ) == ( bv_8_161_n391 )  ;
assign n20844 =  ( n20842 ) & (n20843 )  ;
assign n20845 =  ( n20844 ) & (wr )  ;
assign n20846 =  ( n20845 ) ? ( n5485 ) : ( iram_161 ) ;
assign n20847 = wr_addr[7:7] ;
assign n20848 =  ( n20847 ) == ( bv_1_0_n53 )  ;
assign n20849 =  ( wr_addr ) == ( bv_8_161_n391 )  ;
assign n20850 =  ( n20848 ) & (n20849 )  ;
assign n20851 =  ( n20850 ) & (wr )  ;
assign n20852 =  ( n20851 ) ? ( n5512 ) : ( iram_161 ) ;
assign n20853 = wr_addr[7:7] ;
assign n20854 =  ( n20853 ) == ( bv_1_0_n53 )  ;
assign n20855 =  ( wr_addr ) == ( bv_8_161_n391 )  ;
assign n20856 =  ( n20854 ) & (n20855 )  ;
assign n20857 =  ( n20856 ) & (wr )  ;
assign n20858 =  ( n20857 ) ? ( bv_8_0_n69 ) : ( iram_161 ) ;
assign n20859 = wr_addr[7:7] ;
assign n20860 =  ( n20859 ) == ( bv_1_0_n53 )  ;
assign n20861 =  ( wr_addr ) == ( bv_8_161_n391 )  ;
assign n20862 =  ( n20860 ) & (n20861 )  ;
assign n20863 =  ( n20862 ) & (wr )  ;
assign n20864 =  ( n20863 ) ? ( n5071 ) : ( iram_161 ) ;
assign n20865 = wr_addr[7:7] ;
assign n20866 =  ( n20865 ) == ( bv_1_0_n53 )  ;
assign n20867 =  ( wr_addr ) == ( bv_8_161_n391 )  ;
assign n20868 =  ( n20866 ) & (n20867 )  ;
assign n20869 =  ( n20868 ) & (wr )  ;
assign n20870 =  ( n20869 ) ? ( n5096 ) : ( iram_161 ) ;
assign n20871 = wr_addr[7:7] ;
assign n20872 =  ( n20871 ) == ( bv_1_0_n53 )  ;
assign n20873 =  ( wr_addr ) == ( bv_8_161_n391 )  ;
assign n20874 =  ( n20872 ) & (n20873 )  ;
assign n20875 =  ( n20874 ) & (wr )  ;
assign n20876 =  ( n20875 ) ? ( n5123 ) : ( iram_161 ) ;
assign n20877 = wr_addr[7:7] ;
assign n20878 =  ( n20877 ) == ( bv_1_0_n53 )  ;
assign n20879 =  ( wr_addr ) == ( bv_8_161_n391 )  ;
assign n20880 =  ( n20878 ) & (n20879 )  ;
assign n20881 =  ( n20880 ) & (wr )  ;
assign n20882 =  ( n20881 ) ? ( n5165 ) : ( iram_161 ) ;
assign n20883 = wr_addr[7:7] ;
assign n20884 =  ( n20883 ) == ( bv_1_0_n53 )  ;
assign n20885 =  ( wr_addr ) == ( bv_8_161_n391 )  ;
assign n20886 =  ( n20884 ) & (n20885 )  ;
assign n20887 =  ( n20886 ) & (wr )  ;
assign n20888 =  ( n20887 ) ? ( n5204 ) : ( iram_161 ) ;
assign n20889 = wr_addr[7:7] ;
assign n20890 =  ( n20889 ) == ( bv_1_0_n53 )  ;
assign n20891 =  ( wr_addr ) == ( bv_8_161_n391 )  ;
assign n20892 =  ( n20890 ) & (n20891 )  ;
assign n20893 =  ( n20892 ) & (wr )  ;
assign n20894 =  ( n20893 ) ? ( n5262 ) : ( iram_161 ) ;
assign n20895 = wr_addr[7:7] ;
assign n20896 =  ( n20895 ) == ( bv_1_0_n53 )  ;
assign n20897 =  ( wr_addr ) == ( bv_8_161_n391 )  ;
assign n20898 =  ( n20896 ) & (n20897 )  ;
assign n20899 =  ( n20898 ) & (wr )  ;
assign n20900 =  ( n20899 ) ? ( n5298 ) : ( iram_161 ) ;
assign n20901 = wr_addr[7:7] ;
assign n20902 =  ( n20901 ) == ( bv_1_0_n53 )  ;
assign n20903 =  ( wr_addr ) == ( bv_8_161_n391 )  ;
assign n20904 =  ( n20902 ) & (n20903 )  ;
assign n20905 =  ( n20904 ) & (wr )  ;
assign n20906 =  ( n20905 ) ? ( n5325 ) : ( iram_161 ) ;
assign n20907 = wr_addr[7:7] ;
assign n20908 =  ( n20907 ) == ( bv_1_0_n53 )  ;
assign n20909 =  ( wr_addr ) == ( bv_8_162_n393 )  ;
assign n20910 =  ( n20908 ) & (n20909 )  ;
assign n20911 =  ( n20910 ) & (wr )  ;
assign n20912 =  ( n20911 ) ? ( n4782 ) : ( iram_162 ) ;
assign n20913 = wr_addr[7:7] ;
assign n20914 =  ( n20913 ) == ( bv_1_0_n53 )  ;
assign n20915 =  ( wr_addr ) == ( bv_8_162_n393 )  ;
assign n20916 =  ( n20914 ) & (n20915 )  ;
assign n20917 =  ( n20916 ) & (wr )  ;
assign n20918 =  ( n20917 ) ? ( n4841 ) : ( iram_162 ) ;
assign n20919 = wr_addr[7:7] ;
assign n20920 =  ( n20919 ) == ( bv_1_0_n53 )  ;
assign n20921 =  ( wr_addr ) == ( bv_8_162_n393 )  ;
assign n20922 =  ( n20920 ) & (n20921 )  ;
assign n20923 =  ( n20922 ) & (wr )  ;
assign n20924 =  ( n20923 ) ? ( n5449 ) : ( iram_162 ) ;
assign n20925 = wr_addr[7:7] ;
assign n20926 =  ( n20925 ) == ( bv_1_0_n53 )  ;
assign n20927 =  ( wr_addr ) == ( bv_8_162_n393 )  ;
assign n20928 =  ( n20926 ) & (n20927 )  ;
assign n20929 =  ( n20928 ) & (wr )  ;
assign n20930 =  ( n20929 ) ? ( n4906 ) : ( iram_162 ) ;
assign n20931 = wr_addr[7:7] ;
assign n20932 =  ( n20931 ) == ( bv_1_0_n53 )  ;
assign n20933 =  ( wr_addr ) == ( bv_8_162_n393 )  ;
assign n20934 =  ( n20932 ) & (n20933 )  ;
assign n20935 =  ( n20934 ) & (wr )  ;
assign n20936 =  ( n20935 ) ? ( n5485 ) : ( iram_162 ) ;
assign n20937 = wr_addr[7:7] ;
assign n20938 =  ( n20937 ) == ( bv_1_0_n53 )  ;
assign n20939 =  ( wr_addr ) == ( bv_8_162_n393 )  ;
assign n20940 =  ( n20938 ) & (n20939 )  ;
assign n20941 =  ( n20940 ) & (wr )  ;
assign n20942 =  ( n20941 ) ? ( n5512 ) : ( iram_162 ) ;
assign n20943 = wr_addr[7:7] ;
assign n20944 =  ( n20943 ) == ( bv_1_0_n53 )  ;
assign n20945 =  ( wr_addr ) == ( bv_8_162_n393 )  ;
assign n20946 =  ( n20944 ) & (n20945 )  ;
assign n20947 =  ( n20946 ) & (wr )  ;
assign n20948 =  ( n20947 ) ? ( bv_8_0_n69 ) : ( iram_162 ) ;
assign n20949 = wr_addr[7:7] ;
assign n20950 =  ( n20949 ) == ( bv_1_0_n53 )  ;
assign n20951 =  ( wr_addr ) == ( bv_8_162_n393 )  ;
assign n20952 =  ( n20950 ) & (n20951 )  ;
assign n20953 =  ( n20952 ) & (wr )  ;
assign n20954 =  ( n20953 ) ? ( n5071 ) : ( iram_162 ) ;
assign n20955 = wr_addr[7:7] ;
assign n20956 =  ( n20955 ) == ( bv_1_0_n53 )  ;
assign n20957 =  ( wr_addr ) == ( bv_8_162_n393 )  ;
assign n20958 =  ( n20956 ) & (n20957 )  ;
assign n20959 =  ( n20958 ) & (wr )  ;
assign n20960 =  ( n20959 ) ? ( n5096 ) : ( iram_162 ) ;
assign n20961 = wr_addr[7:7] ;
assign n20962 =  ( n20961 ) == ( bv_1_0_n53 )  ;
assign n20963 =  ( wr_addr ) == ( bv_8_162_n393 )  ;
assign n20964 =  ( n20962 ) & (n20963 )  ;
assign n20965 =  ( n20964 ) & (wr )  ;
assign n20966 =  ( n20965 ) ? ( n5123 ) : ( iram_162 ) ;
assign n20967 = wr_addr[7:7] ;
assign n20968 =  ( n20967 ) == ( bv_1_0_n53 )  ;
assign n20969 =  ( wr_addr ) == ( bv_8_162_n393 )  ;
assign n20970 =  ( n20968 ) & (n20969 )  ;
assign n20971 =  ( n20970 ) & (wr )  ;
assign n20972 =  ( n20971 ) ? ( n5165 ) : ( iram_162 ) ;
assign n20973 = wr_addr[7:7] ;
assign n20974 =  ( n20973 ) == ( bv_1_0_n53 )  ;
assign n20975 =  ( wr_addr ) == ( bv_8_162_n393 )  ;
assign n20976 =  ( n20974 ) & (n20975 )  ;
assign n20977 =  ( n20976 ) & (wr )  ;
assign n20978 =  ( n20977 ) ? ( n5204 ) : ( iram_162 ) ;
assign n20979 = wr_addr[7:7] ;
assign n20980 =  ( n20979 ) == ( bv_1_0_n53 )  ;
assign n20981 =  ( wr_addr ) == ( bv_8_162_n393 )  ;
assign n20982 =  ( n20980 ) & (n20981 )  ;
assign n20983 =  ( n20982 ) & (wr )  ;
assign n20984 =  ( n20983 ) ? ( n5262 ) : ( iram_162 ) ;
assign n20985 = wr_addr[7:7] ;
assign n20986 =  ( n20985 ) == ( bv_1_0_n53 )  ;
assign n20987 =  ( wr_addr ) == ( bv_8_162_n393 )  ;
assign n20988 =  ( n20986 ) & (n20987 )  ;
assign n20989 =  ( n20988 ) & (wr )  ;
assign n20990 =  ( n20989 ) ? ( n5298 ) : ( iram_162 ) ;
assign n20991 = wr_addr[7:7] ;
assign n20992 =  ( n20991 ) == ( bv_1_0_n53 )  ;
assign n20993 =  ( wr_addr ) == ( bv_8_162_n393 )  ;
assign n20994 =  ( n20992 ) & (n20993 )  ;
assign n20995 =  ( n20994 ) & (wr )  ;
assign n20996 =  ( n20995 ) ? ( n5325 ) : ( iram_162 ) ;
assign n20997 = wr_addr[7:7] ;
assign n20998 =  ( n20997 ) == ( bv_1_0_n53 )  ;
assign n20999 =  ( wr_addr ) == ( bv_8_163_n395 )  ;
assign n21000 =  ( n20998 ) & (n20999 )  ;
assign n21001 =  ( n21000 ) & (wr )  ;
assign n21002 =  ( n21001 ) ? ( n4782 ) : ( iram_163 ) ;
assign n21003 = wr_addr[7:7] ;
assign n21004 =  ( n21003 ) == ( bv_1_0_n53 )  ;
assign n21005 =  ( wr_addr ) == ( bv_8_163_n395 )  ;
assign n21006 =  ( n21004 ) & (n21005 )  ;
assign n21007 =  ( n21006 ) & (wr )  ;
assign n21008 =  ( n21007 ) ? ( n4841 ) : ( iram_163 ) ;
assign n21009 = wr_addr[7:7] ;
assign n21010 =  ( n21009 ) == ( bv_1_0_n53 )  ;
assign n21011 =  ( wr_addr ) == ( bv_8_163_n395 )  ;
assign n21012 =  ( n21010 ) & (n21011 )  ;
assign n21013 =  ( n21012 ) & (wr )  ;
assign n21014 =  ( n21013 ) ? ( n5449 ) : ( iram_163 ) ;
assign n21015 = wr_addr[7:7] ;
assign n21016 =  ( n21015 ) == ( bv_1_0_n53 )  ;
assign n21017 =  ( wr_addr ) == ( bv_8_163_n395 )  ;
assign n21018 =  ( n21016 ) & (n21017 )  ;
assign n21019 =  ( n21018 ) & (wr )  ;
assign n21020 =  ( n21019 ) ? ( n4906 ) : ( iram_163 ) ;
assign n21021 = wr_addr[7:7] ;
assign n21022 =  ( n21021 ) == ( bv_1_0_n53 )  ;
assign n21023 =  ( wr_addr ) == ( bv_8_163_n395 )  ;
assign n21024 =  ( n21022 ) & (n21023 )  ;
assign n21025 =  ( n21024 ) & (wr )  ;
assign n21026 =  ( n21025 ) ? ( n5485 ) : ( iram_163 ) ;
assign n21027 = wr_addr[7:7] ;
assign n21028 =  ( n21027 ) == ( bv_1_0_n53 )  ;
assign n21029 =  ( wr_addr ) == ( bv_8_163_n395 )  ;
assign n21030 =  ( n21028 ) & (n21029 )  ;
assign n21031 =  ( n21030 ) & (wr )  ;
assign n21032 =  ( n21031 ) ? ( n5512 ) : ( iram_163 ) ;
assign n21033 = wr_addr[7:7] ;
assign n21034 =  ( n21033 ) == ( bv_1_0_n53 )  ;
assign n21035 =  ( wr_addr ) == ( bv_8_163_n395 )  ;
assign n21036 =  ( n21034 ) & (n21035 )  ;
assign n21037 =  ( n21036 ) & (wr )  ;
assign n21038 =  ( n21037 ) ? ( bv_8_0_n69 ) : ( iram_163 ) ;
assign n21039 = wr_addr[7:7] ;
assign n21040 =  ( n21039 ) == ( bv_1_0_n53 )  ;
assign n21041 =  ( wr_addr ) == ( bv_8_163_n395 )  ;
assign n21042 =  ( n21040 ) & (n21041 )  ;
assign n21043 =  ( n21042 ) & (wr )  ;
assign n21044 =  ( n21043 ) ? ( n5071 ) : ( iram_163 ) ;
assign n21045 = wr_addr[7:7] ;
assign n21046 =  ( n21045 ) == ( bv_1_0_n53 )  ;
assign n21047 =  ( wr_addr ) == ( bv_8_163_n395 )  ;
assign n21048 =  ( n21046 ) & (n21047 )  ;
assign n21049 =  ( n21048 ) & (wr )  ;
assign n21050 =  ( n21049 ) ? ( n5096 ) : ( iram_163 ) ;
assign n21051 = wr_addr[7:7] ;
assign n21052 =  ( n21051 ) == ( bv_1_0_n53 )  ;
assign n21053 =  ( wr_addr ) == ( bv_8_163_n395 )  ;
assign n21054 =  ( n21052 ) & (n21053 )  ;
assign n21055 =  ( n21054 ) & (wr )  ;
assign n21056 =  ( n21055 ) ? ( n5123 ) : ( iram_163 ) ;
assign n21057 = wr_addr[7:7] ;
assign n21058 =  ( n21057 ) == ( bv_1_0_n53 )  ;
assign n21059 =  ( wr_addr ) == ( bv_8_163_n395 )  ;
assign n21060 =  ( n21058 ) & (n21059 )  ;
assign n21061 =  ( n21060 ) & (wr )  ;
assign n21062 =  ( n21061 ) ? ( n5165 ) : ( iram_163 ) ;
assign n21063 = wr_addr[7:7] ;
assign n21064 =  ( n21063 ) == ( bv_1_0_n53 )  ;
assign n21065 =  ( wr_addr ) == ( bv_8_163_n395 )  ;
assign n21066 =  ( n21064 ) & (n21065 )  ;
assign n21067 =  ( n21066 ) & (wr )  ;
assign n21068 =  ( n21067 ) ? ( n5204 ) : ( iram_163 ) ;
assign n21069 = wr_addr[7:7] ;
assign n21070 =  ( n21069 ) == ( bv_1_0_n53 )  ;
assign n21071 =  ( wr_addr ) == ( bv_8_163_n395 )  ;
assign n21072 =  ( n21070 ) & (n21071 )  ;
assign n21073 =  ( n21072 ) & (wr )  ;
assign n21074 =  ( n21073 ) ? ( n5262 ) : ( iram_163 ) ;
assign n21075 = wr_addr[7:7] ;
assign n21076 =  ( n21075 ) == ( bv_1_0_n53 )  ;
assign n21077 =  ( wr_addr ) == ( bv_8_163_n395 )  ;
assign n21078 =  ( n21076 ) & (n21077 )  ;
assign n21079 =  ( n21078 ) & (wr )  ;
assign n21080 =  ( n21079 ) ? ( n5298 ) : ( iram_163 ) ;
assign n21081 = wr_addr[7:7] ;
assign n21082 =  ( n21081 ) == ( bv_1_0_n53 )  ;
assign n21083 =  ( wr_addr ) == ( bv_8_163_n395 )  ;
assign n21084 =  ( n21082 ) & (n21083 )  ;
assign n21085 =  ( n21084 ) & (wr )  ;
assign n21086 =  ( n21085 ) ? ( n5325 ) : ( iram_163 ) ;
assign n21087 = wr_addr[7:7] ;
assign n21088 =  ( n21087 ) == ( bv_1_0_n53 )  ;
assign n21089 =  ( wr_addr ) == ( bv_8_164_n397 )  ;
assign n21090 =  ( n21088 ) & (n21089 )  ;
assign n21091 =  ( n21090 ) & (wr )  ;
assign n21092 =  ( n21091 ) ? ( n4782 ) : ( iram_164 ) ;
assign n21093 = wr_addr[7:7] ;
assign n21094 =  ( n21093 ) == ( bv_1_0_n53 )  ;
assign n21095 =  ( wr_addr ) == ( bv_8_164_n397 )  ;
assign n21096 =  ( n21094 ) & (n21095 )  ;
assign n21097 =  ( n21096 ) & (wr )  ;
assign n21098 =  ( n21097 ) ? ( n4841 ) : ( iram_164 ) ;
assign n21099 = wr_addr[7:7] ;
assign n21100 =  ( n21099 ) == ( bv_1_0_n53 )  ;
assign n21101 =  ( wr_addr ) == ( bv_8_164_n397 )  ;
assign n21102 =  ( n21100 ) & (n21101 )  ;
assign n21103 =  ( n21102 ) & (wr )  ;
assign n21104 =  ( n21103 ) ? ( n5449 ) : ( iram_164 ) ;
assign n21105 = wr_addr[7:7] ;
assign n21106 =  ( n21105 ) == ( bv_1_0_n53 )  ;
assign n21107 =  ( wr_addr ) == ( bv_8_164_n397 )  ;
assign n21108 =  ( n21106 ) & (n21107 )  ;
assign n21109 =  ( n21108 ) & (wr )  ;
assign n21110 =  ( n21109 ) ? ( n4906 ) : ( iram_164 ) ;
assign n21111 = wr_addr[7:7] ;
assign n21112 =  ( n21111 ) == ( bv_1_0_n53 )  ;
assign n21113 =  ( wr_addr ) == ( bv_8_164_n397 )  ;
assign n21114 =  ( n21112 ) & (n21113 )  ;
assign n21115 =  ( n21114 ) & (wr )  ;
assign n21116 =  ( n21115 ) ? ( n5485 ) : ( iram_164 ) ;
assign n21117 = wr_addr[7:7] ;
assign n21118 =  ( n21117 ) == ( bv_1_0_n53 )  ;
assign n21119 =  ( wr_addr ) == ( bv_8_164_n397 )  ;
assign n21120 =  ( n21118 ) & (n21119 )  ;
assign n21121 =  ( n21120 ) & (wr )  ;
assign n21122 =  ( n21121 ) ? ( n5512 ) : ( iram_164 ) ;
assign n21123 = wr_addr[7:7] ;
assign n21124 =  ( n21123 ) == ( bv_1_0_n53 )  ;
assign n21125 =  ( wr_addr ) == ( bv_8_164_n397 )  ;
assign n21126 =  ( n21124 ) & (n21125 )  ;
assign n21127 =  ( n21126 ) & (wr )  ;
assign n21128 =  ( n21127 ) ? ( bv_8_0_n69 ) : ( iram_164 ) ;
assign n21129 = wr_addr[7:7] ;
assign n21130 =  ( n21129 ) == ( bv_1_0_n53 )  ;
assign n21131 =  ( wr_addr ) == ( bv_8_164_n397 )  ;
assign n21132 =  ( n21130 ) & (n21131 )  ;
assign n21133 =  ( n21132 ) & (wr )  ;
assign n21134 =  ( n21133 ) ? ( n5071 ) : ( iram_164 ) ;
assign n21135 = wr_addr[7:7] ;
assign n21136 =  ( n21135 ) == ( bv_1_0_n53 )  ;
assign n21137 =  ( wr_addr ) == ( bv_8_164_n397 )  ;
assign n21138 =  ( n21136 ) & (n21137 )  ;
assign n21139 =  ( n21138 ) & (wr )  ;
assign n21140 =  ( n21139 ) ? ( n5096 ) : ( iram_164 ) ;
assign n21141 = wr_addr[7:7] ;
assign n21142 =  ( n21141 ) == ( bv_1_0_n53 )  ;
assign n21143 =  ( wr_addr ) == ( bv_8_164_n397 )  ;
assign n21144 =  ( n21142 ) & (n21143 )  ;
assign n21145 =  ( n21144 ) & (wr )  ;
assign n21146 =  ( n21145 ) ? ( n5123 ) : ( iram_164 ) ;
assign n21147 = wr_addr[7:7] ;
assign n21148 =  ( n21147 ) == ( bv_1_0_n53 )  ;
assign n21149 =  ( wr_addr ) == ( bv_8_164_n397 )  ;
assign n21150 =  ( n21148 ) & (n21149 )  ;
assign n21151 =  ( n21150 ) & (wr )  ;
assign n21152 =  ( n21151 ) ? ( n5165 ) : ( iram_164 ) ;
assign n21153 = wr_addr[7:7] ;
assign n21154 =  ( n21153 ) == ( bv_1_0_n53 )  ;
assign n21155 =  ( wr_addr ) == ( bv_8_164_n397 )  ;
assign n21156 =  ( n21154 ) & (n21155 )  ;
assign n21157 =  ( n21156 ) & (wr )  ;
assign n21158 =  ( n21157 ) ? ( n5204 ) : ( iram_164 ) ;
assign n21159 = wr_addr[7:7] ;
assign n21160 =  ( n21159 ) == ( bv_1_0_n53 )  ;
assign n21161 =  ( wr_addr ) == ( bv_8_164_n397 )  ;
assign n21162 =  ( n21160 ) & (n21161 )  ;
assign n21163 =  ( n21162 ) & (wr )  ;
assign n21164 =  ( n21163 ) ? ( n5262 ) : ( iram_164 ) ;
assign n21165 = wr_addr[7:7] ;
assign n21166 =  ( n21165 ) == ( bv_1_0_n53 )  ;
assign n21167 =  ( wr_addr ) == ( bv_8_164_n397 )  ;
assign n21168 =  ( n21166 ) & (n21167 )  ;
assign n21169 =  ( n21168 ) & (wr )  ;
assign n21170 =  ( n21169 ) ? ( n5298 ) : ( iram_164 ) ;
assign n21171 = wr_addr[7:7] ;
assign n21172 =  ( n21171 ) == ( bv_1_0_n53 )  ;
assign n21173 =  ( wr_addr ) == ( bv_8_164_n397 )  ;
assign n21174 =  ( n21172 ) & (n21173 )  ;
assign n21175 =  ( n21174 ) & (wr )  ;
assign n21176 =  ( n21175 ) ? ( n5325 ) : ( iram_164 ) ;
assign n21177 = wr_addr[7:7] ;
assign n21178 =  ( n21177 ) == ( bv_1_0_n53 )  ;
assign n21179 =  ( wr_addr ) == ( bv_8_165_n399 )  ;
assign n21180 =  ( n21178 ) & (n21179 )  ;
assign n21181 =  ( n21180 ) & (wr )  ;
assign n21182 =  ( n21181 ) ? ( n4782 ) : ( iram_165 ) ;
assign n21183 = wr_addr[7:7] ;
assign n21184 =  ( n21183 ) == ( bv_1_0_n53 )  ;
assign n21185 =  ( wr_addr ) == ( bv_8_165_n399 )  ;
assign n21186 =  ( n21184 ) & (n21185 )  ;
assign n21187 =  ( n21186 ) & (wr )  ;
assign n21188 =  ( n21187 ) ? ( n4841 ) : ( iram_165 ) ;
assign n21189 = wr_addr[7:7] ;
assign n21190 =  ( n21189 ) == ( bv_1_0_n53 )  ;
assign n21191 =  ( wr_addr ) == ( bv_8_165_n399 )  ;
assign n21192 =  ( n21190 ) & (n21191 )  ;
assign n21193 =  ( n21192 ) & (wr )  ;
assign n21194 =  ( n21193 ) ? ( n5449 ) : ( iram_165 ) ;
assign n21195 = wr_addr[7:7] ;
assign n21196 =  ( n21195 ) == ( bv_1_0_n53 )  ;
assign n21197 =  ( wr_addr ) == ( bv_8_165_n399 )  ;
assign n21198 =  ( n21196 ) & (n21197 )  ;
assign n21199 =  ( n21198 ) & (wr )  ;
assign n21200 =  ( n21199 ) ? ( n4906 ) : ( iram_165 ) ;
assign n21201 = wr_addr[7:7] ;
assign n21202 =  ( n21201 ) == ( bv_1_0_n53 )  ;
assign n21203 =  ( wr_addr ) == ( bv_8_165_n399 )  ;
assign n21204 =  ( n21202 ) & (n21203 )  ;
assign n21205 =  ( n21204 ) & (wr )  ;
assign n21206 =  ( n21205 ) ? ( n5485 ) : ( iram_165 ) ;
assign n21207 = wr_addr[7:7] ;
assign n21208 =  ( n21207 ) == ( bv_1_0_n53 )  ;
assign n21209 =  ( wr_addr ) == ( bv_8_165_n399 )  ;
assign n21210 =  ( n21208 ) & (n21209 )  ;
assign n21211 =  ( n21210 ) & (wr )  ;
assign n21212 =  ( n21211 ) ? ( n5512 ) : ( iram_165 ) ;
assign n21213 = wr_addr[7:7] ;
assign n21214 =  ( n21213 ) == ( bv_1_0_n53 )  ;
assign n21215 =  ( wr_addr ) == ( bv_8_165_n399 )  ;
assign n21216 =  ( n21214 ) & (n21215 )  ;
assign n21217 =  ( n21216 ) & (wr )  ;
assign n21218 =  ( n21217 ) ? ( bv_8_0_n69 ) : ( iram_165 ) ;
assign n21219 = wr_addr[7:7] ;
assign n21220 =  ( n21219 ) == ( bv_1_0_n53 )  ;
assign n21221 =  ( wr_addr ) == ( bv_8_165_n399 )  ;
assign n21222 =  ( n21220 ) & (n21221 )  ;
assign n21223 =  ( n21222 ) & (wr )  ;
assign n21224 =  ( n21223 ) ? ( n5071 ) : ( iram_165 ) ;
assign n21225 = wr_addr[7:7] ;
assign n21226 =  ( n21225 ) == ( bv_1_0_n53 )  ;
assign n21227 =  ( wr_addr ) == ( bv_8_165_n399 )  ;
assign n21228 =  ( n21226 ) & (n21227 )  ;
assign n21229 =  ( n21228 ) & (wr )  ;
assign n21230 =  ( n21229 ) ? ( n5096 ) : ( iram_165 ) ;
assign n21231 = wr_addr[7:7] ;
assign n21232 =  ( n21231 ) == ( bv_1_0_n53 )  ;
assign n21233 =  ( wr_addr ) == ( bv_8_165_n399 )  ;
assign n21234 =  ( n21232 ) & (n21233 )  ;
assign n21235 =  ( n21234 ) & (wr )  ;
assign n21236 =  ( n21235 ) ? ( n5123 ) : ( iram_165 ) ;
assign n21237 = wr_addr[7:7] ;
assign n21238 =  ( n21237 ) == ( bv_1_0_n53 )  ;
assign n21239 =  ( wr_addr ) == ( bv_8_165_n399 )  ;
assign n21240 =  ( n21238 ) & (n21239 )  ;
assign n21241 =  ( n21240 ) & (wr )  ;
assign n21242 =  ( n21241 ) ? ( n5165 ) : ( iram_165 ) ;
assign n21243 = wr_addr[7:7] ;
assign n21244 =  ( n21243 ) == ( bv_1_0_n53 )  ;
assign n21245 =  ( wr_addr ) == ( bv_8_165_n399 )  ;
assign n21246 =  ( n21244 ) & (n21245 )  ;
assign n21247 =  ( n21246 ) & (wr )  ;
assign n21248 =  ( n21247 ) ? ( n5204 ) : ( iram_165 ) ;
assign n21249 = wr_addr[7:7] ;
assign n21250 =  ( n21249 ) == ( bv_1_0_n53 )  ;
assign n21251 =  ( wr_addr ) == ( bv_8_165_n399 )  ;
assign n21252 =  ( n21250 ) & (n21251 )  ;
assign n21253 =  ( n21252 ) & (wr )  ;
assign n21254 =  ( n21253 ) ? ( n5262 ) : ( iram_165 ) ;
assign n21255 = wr_addr[7:7] ;
assign n21256 =  ( n21255 ) == ( bv_1_0_n53 )  ;
assign n21257 =  ( wr_addr ) == ( bv_8_165_n399 )  ;
assign n21258 =  ( n21256 ) & (n21257 )  ;
assign n21259 =  ( n21258 ) & (wr )  ;
assign n21260 =  ( n21259 ) ? ( n5298 ) : ( iram_165 ) ;
assign n21261 = wr_addr[7:7] ;
assign n21262 =  ( n21261 ) == ( bv_1_0_n53 )  ;
assign n21263 =  ( wr_addr ) == ( bv_8_165_n399 )  ;
assign n21264 =  ( n21262 ) & (n21263 )  ;
assign n21265 =  ( n21264 ) & (wr )  ;
assign n21266 =  ( n21265 ) ? ( n5325 ) : ( iram_165 ) ;
assign n21267 = wr_addr[7:7] ;
assign n21268 =  ( n21267 ) == ( bv_1_0_n53 )  ;
assign n21269 =  ( wr_addr ) == ( bv_8_166_n401 )  ;
assign n21270 =  ( n21268 ) & (n21269 )  ;
assign n21271 =  ( n21270 ) & (wr )  ;
assign n21272 =  ( n21271 ) ? ( n4782 ) : ( iram_166 ) ;
assign n21273 = wr_addr[7:7] ;
assign n21274 =  ( n21273 ) == ( bv_1_0_n53 )  ;
assign n21275 =  ( wr_addr ) == ( bv_8_166_n401 )  ;
assign n21276 =  ( n21274 ) & (n21275 )  ;
assign n21277 =  ( n21276 ) & (wr )  ;
assign n21278 =  ( n21277 ) ? ( n4841 ) : ( iram_166 ) ;
assign n21279 = wr_addr[7:7] ;
assign n21280 =  ( n21279 ) == ( bv_1_0_n53 )  ;
assign n21281 =  ( wr_addr ) == ( bv_8_166_n401 )  ;
assign n21282 =  ( n21280 ) & (n21281 )  ;
assign n21283 =  ( n21282 ) & (wr )  ;
assign n21284 =  ( n21283 ) ? ( n5449 ) : ( iram_166 ) ;
assign n21285 = wr_addr[7:7] ;
assign n21286 =  ( n21285 ) == ( bv_1_0_n53 )  ;
assign n21287 =  ( wr_addr ) == ( bv_8_166_n401 )  ;
assign n21288 =  ( n21286 ) & (n21287 )  ;
assign n21289 =  ( n21288 ) & (wr )  ;
assign n21290 =  ( n21289 ) ? ( n4906 ) : ( iram_166 ) ;
assign n21291 = wr_addr[7:7] ;
assign n21292 =  ( n21291 ) == ( bv_1_0_n53 )  ;
assign n21293 =  ( wr_addr ) == ( bv_8_166_n401 )  ;
assign n21294 =  ( n21292 ) & (n21293 )  ;
assign n21295 =  ( n21294 ) & (wr )  ;
assign n21296 =  ( n21295 ) ? ( n5485 ) : ( iram_166 ) ;
assign n21297 = wr_addr[7:7] ;
assign n21298 =  ( n21297 ) == ( bv_1_0_n53 )  ;
assign n21299 =  ( wr_addr ) == ( bv_8_166_n401 )  ;
assign n21300 =  ( n21298 ) & (n21299 )  ;
assign n21301 =  ( n21300 ) & (wr )  ;
assign n21302 =  ( n21301 ) ? ( n5512 ) : ( iram_166 ) ;
assign n21303 = wr_addr[7:7] ;
assign n21304 =  ( n21303 ) == ( bv_1_0_n53 )  ;
assign n21305 =  ( wr_addr ) == ( bv_8_166_n401 )  ;
assign n21306 =  ( n21304 ) & (n21305 )  ;
assign n21307 =  ( n21306 ) & (wr )  ;
assign n21308 =  ( n21307 ) ? ( bv_8_0_n69 ) : ( iram_166 ) ;
assign n21309 = wr_addr[7:7] ;
assign n21310 =  ( n21309 ) == ( bv_1_0_n53 )  ;
assign n21311 =  ( wr_addr ) == ( bv_8_166_n401 )  ;
assign n21312 =  ( n21310 ) & (n21311 )  ;
assign n21313 =  ( n21312 ) & (wr )  ;
assign n21314 =  ( n21313 ) ? ( n5071 ) : ( iram_166 ) ;
assign n21315 = wr_addr[7:7] ;
assign n21316 =  ( n21315 ) == ( bv_1_0_n53 )  ;
assign n21317 =  ( wr_addr ) == ( bv_8_166_n401 )  ;
assign n21318 =  ( n21316 ) & (n21317 )  ;
assign n21319 =  ( n21318 ) & (wr )  ;
assign n21320 =  ( n21319 ) ? ( n5096 ) : ( iram_166 ) ;
assign n21321 = wr_addr[7:7] ;
assign n21322 =  ( n21321 ) == ( bv_1_0_n53 )  ;
assign n21323 =  ( wr_addr ) == ( bv_8_166_n401 )  ;
assign n21324 =  ( n21322 ) & (n21323 )  ;
assign n21325 =  ( n21324 ) & (wr )  ;
assign n21326 =  ( n21325 ) ? ( n5123 ) : ( iram_166 ) ;
assign n21327 = wr_addr[7:7] ;
assign n21328 =  ( n21327 ) == ( bv_1_0_n53 )  ;
assign n21329 =  ( wr_addr ) == ( bv_8_166_n401 )  ;
assign n21330 =  ( n21328 ) & (n21329 )  ;
assign n21331 =  ( n21330 ) & (wr )  ;
assign n21332 =  ( n21331 ) ? ( n5165 ) : ( iram_166 ) ;
assign n21333 = wr_addr[7:7] ;
assign n21334 =  ( n21333 ) == ( bv_1_0_n53 )  ;
assign n21335 =  ( wr_addr ) == ( bv_8_166_n401 )  ;
assign n21336 =  ( n21334 ) & (n21335 )  ;
assign n21337 =  ( n21336 ) & (wr )  ;
assign n21338 =  ( n21337 ) ? ( n5204 ) : ( iram_166 ) ;
assign n21339 = wr_addr[7:7] ;
assign n21340 =  ( n21339 ) == ( bv_1_0_n53 )  ;
assign n21341 =  ( wr_addr ) == ( bv_8_166_n401 )  ;
assign n21342 =  ( n21340 ) & (n21341 )  ;
assign n21343 =  ( n21342 ) & (wr )  ;
assign n21344 =  ( n21343 ) ? ( n5262 ) : ( iram_166 ) ;
assign n21345 = wr_addr[7:7] ;
assign n21346 =  ( n21345 ) == ( bv_1_0_n53 )  ;
assign n21347 =  ( wr_addr ) == ( bv_8_166_n401 )  ;
assign n21348 =  ( n21346 ) & (n21347 )  ;
assign n21349 =  ( n21348 ) & (wr )  ;
assign n21350 =  ( n21349 ) ? ( n5298 ) : ( iram_166 ) ;
assign n21351 = wr_addr[7:7] ;
assign n21352 =  ( n21351 ) == ( bv_1_0_n53 )  ;
assign n21353 =  ( wr_addr ) == ( bv_8_166_n401 )  ;
assign n21354 =  ( n21352 ) & (n21353 )  ;
assign n21355 =  ( n21354 ) & (wr )  ;
assign n21356 =  ( n21355 ) ? ( n5325 ) : ( iram_166 ) ;
assign n21357 = wr_addr[7:7] ;
assign n21358 =  ( n21357 ) == ( bv_1_0_n53 )  ;
assign n21359 =  ( wr_addr ) == ( bv_8_167_n403 )  ;
assign n21360 =  ( n21358 ) & (n21359 )  ;
assign n21361 =  ( n21360 ) & (wr )  ;
assign n21362 =  ( n21361 ) ? ( n4782 ) : ( iram_167 ) ;
assign n21363 = wr_addr[7:7] ;
assign n21364 =  ( n21363 ) == ( bv_1_0_n53 )  ;
assign n21365 =  ( wr_addr ) == ( bv_8_167_n403 )  ;
assign n21366 =  ( n21364 ) & (n21365 )  ;
assign n21367 =  ( n21366 ) & (wr )  ;
assign n21368 =  ( n21367 ) ? ( n4841 ) : ( iram_167 ) ;
assign n21369 = wr_addr[7:7] ;
assign n21370 =  ( n21369 ) == ( bv_1_0_n53 )  ;
assign n21371 =  ( wr_addr ) == ( bv_8_167_n403 )  ;
assign n21372 =  ( n21370 ) & (n21371 )  ;
assign n21373 =  ( n21372 ) & (wr )  ;
assign n21374 =  ( n21373 ) ? ( n5449 ) : ( iram_167 ) ;
assign n21375 = wr_addr[7:7] ;
assign n21376 =  ( n21375 ) == ( bv_1_0_n53 )  ;
assign n21377 =  ( wr_addr ) == ( bv_8_167_n403 )  ;
assign n21378 =  ( n21376 ) & (n21377 )  ;
assign n21379 =  ( n21378 ) & (wr )  ;
assign n21380 =  ( n21379 ) ? ( n4906 ) : ( iram_167 ) ;
assign n21381 = wr_addr[7:7] ;
assign n21382 =  ( n21381 ) == ( bv_1_0_n53 )  ;
assign n21383 =  ( wr_addr ) == ( bv_8_167_n403 )  ;
assign n21384 =  ( n21382 ) & (n21383 )  ;
assign n21385 =  ( n21384 ) & (wr )  ;
assign n21386 =  ( n21385 ) ? ( n5485 ) : ( iram_167 ) ;
assign n21387 = wr_addr[7:7] ;
assign n21388 =  ( n21387 ) == ( bv_1_0_n53 )  ;
assign n21389 =  ( wr_addr ) == ( bv_8_167_n403 )  ;
assign n21390 =  ( n21388 ) & (n21389 )  ;
assign n21391 =  ( n21390 ) & (wr )  ;
assign n21392 =  ( n21391 ) ? ( n5512 ) : ( iram_167 ) ;
assign n21393 = wr_addr[7:7] ;
assign n21394 =  ( n21393 ) == ( bv_1_0_n53 )  ;
assign n21395 =  ( wr_addr ) == ( bv_8_167_n403 )  ;
assign n21396 =  ( n21394 ) & (n21395 )  ;
assign n21397 =  ( n21396 ) & (wr )  ;
assign n21398 =  ( n21397 ) ? ( bv_8_0_n69 ) : ( iram_167 ) ;
assign n21399 = wr_addr[7:7] ;
assign n21400 =  ( n21399 ) == ( bv_1_0_n53 )  ;
assign n21401 =  ( wr_addr ) == ( bv_8_167_n403 )  ;
assign n21402 =  ( n21400 ) & (n21401 )  ;
assign n21403 =  ( n21402 ) & (wr )  ;
assign n21404 =  ( n21403 ) ? ( n5071 ) : ( iram_167 ) ;
assign n21405 = wr_addr[7:7] ;
assign n21406 =  ( n21405 ) == ( bv_1_0_n53 )  ;
assign n21407 =  ( wr_addr ) == ( bv_8_167_n403 )  ;
assign n21408 =  ( n21406 ) & (n21407 )  ;
assign n21409 =  ( n21408 ) & (wr )  ;
assign n21410 =  ( n21409 ) ? ( n5096 ) : ( iram_167 ) ;
assign n21411 = wr_addr[7:7] ;
assign n21412 =  ( n21411 ) == ( bv_1_0_n53 )  ;
assign n21413 =  ( wr_addr ) == ( bv_8_167_n403 )  ;
assign n21414 =  ( n21412 ) & (n21413 )  ;
assign n21415 =  ( n21414 ) & (wr )  ;
assign n21416 =  ( n21415 ) ? ( n5123 ) : ( iram_167 ) ;
assign n21417 = wr_addr[7:7] ;
assign n21418 =  ( n21417 ) == ( bv_1_0_n53 )  ;
assign n21419 =  ( wr_addr ) == ( bv_8_167_n403 )  ;
assign n21420 =  ( n21418 ) & (n21419 )  ;
assign n21421 =  ( n21420 ) & (wr )  ;
assign n21422 =  ( n21421 ) ? ( n5165 ) : ( iram_167 ) ;
assign n21423 = wr_addr[7:7] ;
assign n21424 =  ( n21423 ) == ( bv_1_0_n53 )  ;
assign n21425 =  ( wr_addr ) == ( bv_8_167_n403 )  ;
assign n21426 =  ( n21424 ) & (n21425 )  ;
assign n21427 =  ( n21426 ) & (wr )  ;
assign n21428 =  ( n21427 ) ? ( n5204 ) : ( iram_167 ) ;
assign n21429 = wr_addr[7:7] ;
assign n21430 =  ( n21429 ) == ( bv_1_0_n53 )  ;
assign n21431 =  ( wr_addr ) == ( bv_8_167_n403 )  ;
assign n21432 =  ( n21430 ) & (n21431 )  ;
assign n21433 =  ( n21432 ) & (wr )  ;
assign n21434 =  ( n21433 ) ? ( n5262 ) : ( iram_167 ) ;
assign n21435 = wr_addr[7:7] ;
assign n21436 =  ( n21435 ) == ( bv_1_0_n53 )  ;
assign n21437 =  ( wr_addr ) == ( bv_8_167_n403 )  ;
assign n21438 =  ( n21436 ) & (n21437 )  ;
assign n21439 =  ( n21438 ) & (wr )  ;
assign n21440 =  ( n21439 ) ? ( n5298 ) : ( iram_167 ) ;
assign n21441 = wr_addr[7:7] ;
assign n21442 =  ( n21441 ) == ( bv_1_0_n53 )  ;
assign n21443 =  ( wr_addr ) == ( bv_8_167_n403 )  ;
assign n21444 =  ( n21442 ) & (n21443 )  ;
assign n21445 =  ( n21444 ) & (wr )  ;
assign n21446 =  ( n21445 ) ? ( n5325 ) : ( iram_167 ) ;
assign n21447 = wr_addr[7:7] ;
assign n21448 =  ( n21447 ) == ( bv_1_0_n53 )  ;
assign n21449 =  ( wr_addr ) == ( bv_8_168_n405 )  ;
assign n21450 =  ( n21448 ) & (n21449 )  ;
assign n21451 =  ( n21450 ) & (wr )  ;
assign n21452 =  ( n21451 ) ? ( n4782 ) : ( iram_168 ) ;
assign n21453 = wr_addr[7:7] ;
assign n21454 =  ( n21453 ) == ( bv_1_0_n53 )  ;
assign n21455 =  ( wr_addr ) == ( bv_8_168_n405 )  ;
assign n21456 =  ( n21454 ) & (n21455 )  ;
assign n21457 =  ( n21456 ) & (wr )  ;
assign n21458 =  ( n21457 ) ? ( n4841 ) : ( iram_168 ) ;
assign n21459 = wr_addr[7:7] ;
assign n21460 =  ( n21459 ) == ( bv_1_0_n53 )  ;
assign n21461 =  ( wr_addr ) == ( bv_8_168_n405 )  ;
assign n21462 =  ( n21460 ) & (n21461 )  ;
assign n21463 =  ( n21462 ) & (wr )  ;
assign n21464 =  ( n21463 ) ? ( n5449 ) : ( iram_168 ) ;
assign n21465 = wr_addr[7:7] ;
assign n21466 =  ( n21465 ) == ( bv_1_0_n53 )  ;
assign n21467 =  ( wr_addr ) == ( bv_8_168_n405 )  ;
assign n21468 =  ( n21466 ) & (n21467 )  ;
assign n21469 =  ( n21468 ) & (wr )  ;
assign n21470 =  ( n21469 ) ? ( n4906 ) : ( iram_168 ) ;
assign n21471 = wr_addr[7:7] ;
assign n21472 =  ( n21471 ) == ( bv_1_0_n53 )  ;
assign n21473 =  ( wr_addr ) == ( bv_8_168_n405 )  ;
assign n21474 =  ( n21472 ) & (n21473 )  ;
assign n21475 =  ( n21474 ) & (wr )  ;
assign n21476 =  ( n21475 ) ? ( n5485 ) : ( iram_168 ) ;
assign n21477 = wr_addr[7:7] ;
assign n21478 =  ( n21477 ) == ( bv_1_0_n53 )  ;
assign n21479 =  ( wr_addr ) == ( bv_8_168_n405 )  ;
assign n21480 =  ( n21478 ) & (n21479 )  ;
assign n21481 =  ( n21480 ) & (wr )  ;
assign n21482 =  ( n21481 ) ? ( n5512 ) : ( iram_168 ) ;
assign n21483 = wr_addr[7:7] ;
assign n21484 =  ( n21483 ) == ( bv_1_0_n53 )  ;
assign n21485 =  ( wr_addr ) == ( bv_8_168_n405 )  ;
assign n21486 =  ( n21484 ) & (n21485 )  ;
assign n21487 =  ( n21486 ) & (wr )  ;
assign n21488 =  ( n21487 ) ? ( bv_8_0_n69 ) : ( iram_168 ) ;
assign n21489 = wr_addr[7:7] ;
assign n21490 =  ( n21489 ) == ( bv_1_0_n53 )  ;
assign n21491 =  ( wr_addr ) == ( bv_8_168_n405 )  ;
assign n21492 =  ( n21490 ) & (n21491 )  ;
assign n21493 =  ( n21492 ) & (wr )  ;
assign n21494 =  ( n21493 ) ? ( n5071 ) : ( iram_168 ) ;
assign n21495 = wr_addr[7:7] ;
assign n21496 =  ( n21495 ) == ( bv_1_0_n53 )  ;
assign n21497 =  ( wr_addr ) == ( bv_8_168_n405 )  ;
assign n21498 =  ( n21496 ) & (n21497 )  ;
assign n21499 =  ( n21498 ) & (wr )  ;
assign n21500 =  ( n21499 ) ? ( n5096 ) : ( iram_168 ) ;
assign n21501 = wr_addr[7:7] ;
assign n21502 =  ( n21501 ) == ( bv_1_0_n53 )  ;
assign n21503 =  ( wr_addr ) == ( bv_8_168_n405 )  ;
assign n21504 =  ( n21502 ) & (n21503 )  ;
assign n21505 =  ( n21504 ) & (wr )  ;
assign n21506 =  ( n21505 ) ? ( n5123 ) : ( iram_168 ) ;
assign n21507 = wr_addr[7:7] ;
assign n21508 =  ( n21507 ) == ( bv_1_0_n53 )  ;
assign n21509 =  ( wr_addr ) == ( bv_8_168_n405 )  ;
assign n21510 =  ( n21508 ) & (n21509 )  ;
assign n21511 =  ( n21510 ) & (wr )  ;
assign n21512 =  ( n21511 ) ? ( n5165 ) : ( iram_168 ) ;
assign n21513 = wr_addr[7:7] ;
assign n21514 =  ( n21513 ) == ( bv_1_0_n53 )  ;
assign n21515 =  ( wr_addr ) == ( bv_8_168_n405 )  ;
assign n21516 =  ( n21514 ) & (n21515 )  ;
assign n21517 =  ( n21516 ) & (wr )  ;
assign n21518 =  ( n21517 ) ? ( n5204 ) : ( iram_168 ) ;
assign n21519 = wr_addr[7:7] ;
assign n21520 =  ( n21519 ) == ( bv_1_0_n53 )  ;
assign n21521 =  ( wr_addr ) == ( bv_8_168_n405 )  ;
assign n21522 =  ( n21520 ) & (n21521 )  ;
assign n21523 =  ( n21522 ) & (wr )  ;
assign n21524 =  ( n21523 ) ? ( n5262 ) : ( iram_168 ) ;
assign n21525 = wr_addr[7:7] ;
assign n21526 =  ( n21525 ) == ( bv_1_0_n53 )  ;
assign n21527 =  ( wr_addr ) == ( bv_8_168_n405 )  ;
assign n21528 =  ( n21526 ) & (n21527 )  ;
assign n21529 =  ( n21528 ) & (wr )  ;
assign n21530 =  ( n21529 ) ? ( n5298 ) : ( iram_168 ) ;
assign n21531 = wr_addr[7:7] ;
assign n21532 =  ( n21531 ) == ( bv_1_0_n53 )  ;
assign n21533 =  ( wr_addr ) == ( bv_8_168_n405 )  ;
assign n21534 =  ( n21532 ) & (n21533 )  ;
assign n21535 =  ( n21534 ) & (wr )  ;
assign n21536 =  ( n21535 ) ? ( n5325 ) : ( iram_168 ) ;
assign n21537 = wr_addr[7:7] ;
assign n21538 =  ( n21537 ) == ( bv_1_0_n53 )  ;
assign n21539 =  ( wr_addr ) == ( bv_8_169_n407 )  ;
assign n21540 =  ( n21538 ) & (n21539 )  ;
assign n21541 =  ( n21540 ) & (wr )  ;
assign n21542 =  ( n21541 ) ? ( n4782 ) : ( iram_169 ) ;
assign n21543 = wr_addr[7:7] ;
assign n21544 =  ( n21543 ) == ( bv_1_0_n53 )  ;
assign n21545 =  ( wr_addr ) == ( bv_8_169_n407 )  ;
assign n21546 =  ( n21544 ) & (n21545 )  ;
assign n21547 =  ( n21546 ) & (wr )  ;
assign n21548 =  ( n21547 ) ? ( n4841 ) : ( iram_169 ) ;
assign n21549 = wr_addr[7:7] ;
assign n21550 =  ( n21549 ) == ( bv_1_0_n53 )  ;
assign n21551 =  ( wr_addr ) == ( bv_8_169_n407 )  ;
assign n21552 =  ( n21550 ) & (n21551 )  ;
assign n21553 =  ( n21552 ) & (wr )  ;
assign n21554 =  ( n21553 ) ? ( n5449 ) : ( iram_169 ) ;
assign n21555 = wr_addr[7:7] ;
assign n21556 =  ( n21555 ) == ( bv_1_0_n53 )  ;
assign n21557 =  ( wr_addr ) == ( bv_8_169_n407 )  ;
assign n21558 =  ( n21556 ) & (n21557 )  ;
assign n21559 =  ( n21558 ) & (wr )  ;
assign n21560 =  ( n21559 ) ? ( n4906 ) : ( iram_169 ) ;
assign n21561 = wr_addr[7:7] ;
assign n21562 =  ( n21561 ) == ( bv_1_0_n53 )  ;
assign n21563 =  ( wr_addr ) == ( bv_8_169_n407 )  ;
assign n21564 =  ( n21562 ) & (n21563 )  ;
assign n21565 =  ( n21564 ) & (wr )  ;
assign n21566 =  ( n21565 ) ? ( n5485 ) : ( iram_169 ) ;
assign n21567 = wr_addr[7:7] ;
assign n21568 =  ( n21567 ) == ( bv_1_0_n53 )  ;
assign n21569 =  ( wr_addr ) == ( bv_8_169_n407 )  ;
assign n21570 =  ( n21568 ) & (n21569 )  ;
assign n21571 =  ( n21570 ) & (wr )  ;
assign n21572 =  ( n21571 ) ? ( n5512 ) : ( iram_169 ) ;
assign n21573 = wr_addr[7:7] ;
assign n21574 =  ( n21573 ) == ( bv_1_0_n53 )  ;
assign n21575 =  ( wr_addr ) == ( bv_8_169_n407 )  ;
assign n21576 =  ( n21574 ) & (n21575 )  ;
assign n21577 =  ( n21576 ) & (wr )  ;
assign n21578 =  ( n21577 ) ? ( bv_8_0_n69 ) : ( iram_169 ) ;
assign n21579 = wr_addr[7:7] ;
assign n21580 =  ( n21579 ) == ( bv_1_0_n53 )  ;
assign n21581 =  ( wr_addr ) == ( bv_8_169_n407 )  ;
assign n21582 =  ( n21580 ) & (n21581 )  ;
assign n21583 =  ( n21582 ) & (wr )  ;
assign n21584 =  ( n21583 ) ? ( n5071 ) : ( iram_169 ) ;
assign n21585 = wr_addr[7:7] ;
assign n21586 =  ( n21585 ) == ( bv_1_0_n53 )  ;
assign n21587 =  ( wr_addr ) == ( bv_8_169_n407 )  ;
assign n21588 =  ( n21586 ) & (n21587 )  ;
assign n21589 =  ( n21588 ) & (wr )  ;
assign n21590 =  ( n21589 ) ? ( n5096 ) : ( iram_169 ) ;
assign n21591 = wr_addr[7:7] ;
assign n21592 =  ( n21591 ) == ( bv_1_0_n53 )  ;
assign n21593 =  ( wr_addr ) == ( bv_8_169_n407 )  ;
assign n21594 =  ( n21592 ) & (n21593 )  ;
assign n21595 =  ( n21594 ) & (wr )  ;
assign n21596 =  ( n21595 ) ? ( n5123 ) : ( iram_169 ) ;
assign n21597 = wr_addr[7:7] ;
assign n21598 =  ( n21597 ) == ( bv_1_0_n53 )  ;
assign n21599 =  ( wr_addr ) == ( bv_8_169_n407 )  ;
assign n21600 =  ( n21598 ) & (n21599 )  ;
assign n21601 =  ( n21600 ) & (wr )  ;
assign n21602 =  ( n21601 ) ? ( n5165 ) : ( iram_169 ) ;
assign n21603 = wr_addr[7:7] ;
assign n21604 =  ( n21603 ) == ( bv_1_0_n53 )  ;
assign n21605 =  ( wr_addr ) == ( bv_8_169_n407 )  ;
assign n21606 =  ( n21604 ) & (n21605 )  ;
assign n21607 =  ( n21606 ) & (wr )  ;
assign n21608 =  ( n21607 ) ? ( n5204 ) : ( iram_169 ) ;
assign n21609 = wr_addr[7:7] ;
assign n21610 =  ( n21609 ) == ( bv_1_0_n53 )  ;
assign n21611 =  ( wr_addr ) == ( bv_8_169_n407 )  ;
assign n21612 =  ( n21610 ) & (n21611 )  ;
assign n21613 =  ( n21612 ) & (wr )  ;
assign n21614 =  ( n21613 ) ? ( n5262 ) : ( iram_169 ) ;
assign n21615 = wr_addr[7:7] ;
assign n21616 =  ( n21615 ) == ( bv_1_0_n53 )  ;
assign n21617 =  ( wr_addr ) == ( bv_8_169_n407 )  ;
assign n21618 =  ( n21616 ) & (n21617 )  ;
assign n21619 =  ( n21618 ) & (wr )  ;
assign n21620 =  ( n21619 ) ? ( n5298 ) : ( iram_169 ) ;
assign n21621 = wr_addr[7:7] ;
assign n21622 =  ( n21621 ) == ( bv_1_0_n53 )  ;
assign n21623 =  ( wr_addr ) == ( bv_8_169_n407 )  ;
assign n21624 =  ( n21622 ) & (n21623 )  ;
assign n21625 =  ( n21624 ) & (wr )  ;
assign n21626 =  ( n21625 ) ? ( n5325 ) : ( iram_169 ) ;
assign n21627 = wr_addr[7:7] ;
assign n21628 =  ( n21627 ) == ( bv_1_0_n53 )  ;
assign n21629 =  ( wr_addr ) == ( bv_8_170_n409 )  ;
assign n21630 =  ( n21628 ) & (n21629 )  ;
assign n21631 =  ( n21630 ) & (wr )  ;
assign n21632 =  ( n21631 ) ? ( n4782 ) : ( iram_170 ) ;
assign n21633 = wr_addr[7:7] ;
assign n21634 =  ( n21633 ) == ( bv_1_0_n53 )  ;
assign n21635 =  ( wr_addr ) == ( bv_8_170_n409 )  ;
assign n21636 =  ( n21634 ) & (n21635 )  ;
assign n21637 =  ( n21636 ) & (wr )  ;
assign n21638 =  ( n21637 ) ? ( n4841 ) : ( iram_170 ) ;
assign n21639 = wr_addr[7:7] ;
assign n21640 =  ( n21639 ) == ( bv_1_0_n53 )  ;
assign n21641 =  ( wr_addr ) == ( bv_8_170_n409 )  ;
assign n21642 =  ( n21640 ) & (n21641 )  ;
assign n21643 =  ( n21642 ) & (wr )  ;
assign n21644 =  ( n21643 ) ? ( n5449 ) : ( iram_170 ) ;
assign n21645 = wr_addr[7:7] ;
assign n21646 =  ( n21645 ) == ( bv_1_0_n53 )  ;
assign n21647 =  ( wr_addr ) == ( bv_8_170_n409 )  ;
assign n21648 =  ( n21646 ) & (n21647 )  ;
assign n21649 =  ( n21648 ) & (wr )  ;
assign n21650 =  ( n21649 ) ? ( n4906 ) : ( iram_170 ) ;
assign n21651 = wr_addr[7:7] ;
assign n21652 =  ( n21651 ) == ( bv_1_0_n53 )  ;
assign n21653 =  ( wr_addr ) == ( bv_8_170_n409 )  ;
assign n21654 =  ( n21652 ) & (n21653 )  ;
assign n21655 =  ( n21654 ) & (wr )  ;
assign n21656 =  ( n21655 ) ? ( n5485 ) : ( iram_170 ) ;
assign n21657 = wr_addr[7:7] ;
assign n21658 =  ( n21657 ) == ( bv_1_0_n53 )  ;
assign n21659 =  ( wr_addr ) == ( bv_8_170_n409 )  ;
assign n21660 =  ( n21658 ) & (n21659 )  ;
assign n21661 =  ( n21660 ) & (wr )  ;
assign n21662 =  ( n21661 ) ? ( n5512 ) : ( iram_170 ) ;
assign n21663 = wr_addr[7:7] ;
assign n21664 =  ( n21663 ) == ( bv_1_0_n53 )  ;
assign n21665 =  ( wr_addr ) == ( bv_8_170_n409 )  ;
assign n21666 =  ( n21664 ) & (n21665 )  ;
assign n21667 =  ( n21666 ) & (wr )  ;
assign n21668 =  ( n21667 ) ? ( bv_8_0_n69 ) : ( iram_170 ) ;
assign n21669 = wr_addr[7:7] ;
assign n21670 =  ( n21669 ) == ( bv_1_0_n53 )  ;
assign n21671 =  ( wr_addr ) == ( bv_8_170_n409 )  ;
assign n21672 =  ( n21670 ) & (n21671 )  ;
assign n21673 =  ( n21672 ) & (wr )  ;
assign n21674 =  ( n21673 ) ? ( n5071 ) : ( iram_170 ) ;
assign n21675 = wr_addr[7:7] ;
assign n21676 =  ( n21675 ) == ( bv_1_0_n53 )  ;
assign n21677 =  ( wr_addr ) == ( bv_8_170_n409 )  ;
assign n21678 =  ( n21676 ) & (n21677 )  ;
assign n21679 =  ( n21678 ) & (wr )  ;
assign n21680 =  ( n21679 ) ? ( n5096 ) : ( iram_170 ) ;
assign n21681 = wr_addr[7:7] ;
assign n21682 =  ( n21681 ) == ( bv_1_0_n53 )  ;
assign n21683 =  ( wr_addr ) == ( bv_8_170_n409 )  ;
assign n21684 =  ( n21682 ) & (n21683 )  ;
assign n21685 =  ( n21684 ) & (wr )  ;
assign n21686 =  ( n21685 ) ? ( n5123 ) : ( iram_170 ) ;
assign n21687 = wr_addr[7:7] ;
assign n21688 =  ( n21687 ) == ( bv_1_0_n53 )  ;
assign n21689 =  ( wr_addr ) == ( bv_8_170_n409 )  ;
assign n21690 =  ( n21688 ) & (n21689 )  ;
assign n21691 =  ( n21690 ) & (wr )  ;
assign n21692 =  ( n21691 ) ? ( n5165 ) : ( iram_170 ) ;
assign n21693 = wr_addr[7:7] ;
assign n21694 =  ( n21693 ) == ( bv_1_0_n53 )  ;
assign n21695 =  ( wr_addr ) == ( bv_8_170_n409 )  ;
assign n21696 =  ( n21694 ) & (n21695 )  ;
assign n21697 =  ( n21696 ) & (wr )  ;
assign n21698 =  ( n21697 ) ? ( n5204 ) : ( iram_170 ) ;
assign n21699 = wr_addr[7:7] ;
assign n21700 =  ( n21699 ) == ( bv_1_0_n53 )  ;
assign n21701 =  ( wr_addr ) == ( bv_8_170_n409 )  ;
assign n21702 =  ( n21700 ) & (n21701 )  ;
assign n21703 =  ( n21702 ) & (wr )  ;
assign n21704 =  ( n21703 ) ? ( n5262 ) : ( iram_170 ) ;
assign n21705 = wr_addr[7:7] ;
assign n21706 =  ( n21705 ) == ( bv_1_0_n53 )  ;
assign n21707 =  ( wr_addr ) == ( bv_8_170_n409 )  ;
assign n21708 =  ( n21706 ) & (n21707 )  ;
assign n21709 =  ( n21708 ) & (wr )  ;
assign n21710 =  ( n21709 ) ? ( n5298 ) : ( iram_170 ) ;
assign n21711 = wr_addr[7:7] ;
assign n21712 =  ( n21711 ) == ( bv_1_0_n53 )  ;
assign n21713 =  ( wr_addr ) == ( bv_8_170_n409 )  ;
assign n21714 =  ( n21712 ) & (n21713 )  ;
assign n21715 =  ( n21714 ) & (wr )  ;
assign n21716 =  ( n21715 ) ? ( n5325 ) : ( iram_170 ) ;
assign n21717 = wr_addr[7:7] ;
assign n21718 =  ( n21717 ) == ( bv_1_0_n53 )  ;
assign n21719 =  ( wr_addr ) == ( bv_8_171_n411 )  ;
assign n21720 =  ( n21718 ) & (n21719 )  ;
assign n21721 =  ( n21720 ) & (wr )  ;
assign n21722 =  ( n21721 ) ? ( n4782 ) : ( iram_171 ) ;
assign n21723 = wr_addr[7:7] ;
assign n21724 =  ( n21723 ) == ( bv_1_0_n53 )  ;
assign n21725 =  ( wr_addr ) == ( bv_8_171_n411 )  ;
assign n21726 =  ( n21724 ) & (n21725 )  ;
assign n21727 =  ( n21726 ) & (wr )  ;
assign n21728 =  ( n21727 ) ? ( n4841 ) : ( iram_171 ) ;
assign n21729 = wr_addr[7:7] ;
assign n21730 =  ( n21729 ) == ( bv_1_0_n53 )  ;
assign n21731 =  ( wr_addr ) == ( bv_8_171_n411 )  ;
assign n21732 =  ( n21730 ) & (n21731 )  ;
assign n21733 =  ( n21732 ) & (wr )  ;
assign n21734 =  ( n21733 ) ? ( n5449 ) : ( iram_171 ) ;
assign n21735 = wr_addr[7:7] ;
assign n21736 =  ( n21735 ) == ( bv_1_0_n53 )  ;
assign n21737 =  ( wr_addr ) == ( bv_8_171_n411 )  ;
assign n21738 =  ( n21736 ) & (n21737 )  ;
assign n21739 =  ( n21738 ) & (wr )  ;
assign n21740 =  ( n21739 ) ? ( n4906 ) : ( iram_171 ) ;
assign n21741 = wr_addr[7:7] ;
assign n21742 =  ( n21741 ) == ( bv_1_0_n53 )  ;
assign n21743 =  ( wr_addr ) == ( bv_8_171_n411 )  ;
assign n21744 =  ( n21742 ) & (n21743 )  ;
assign n21745 =  ( n21744 ) & (wr )  ;
assign n21746 =  ( n21745 ) ? ( n5485 ) : ( iram_171 ) ;
assign n21747 = wr_addr[7:7] ;
assign n21748 =  ( n21747 ) == ( bv_1_0_n53 )  ;
assign n21749 =  ( wr_addr ) == ( bv_8_171_n411 )  ;
assign n21750 =  ( n21748 ) & (n21749 )  ;
assign n21751 =  ( n21750 ) & (wr )  ;
assign n21752 =  ( n21751 ) ? ( n5512 ) : ( iram_171 ) ;
assign n21753 = wr_addr[7:7] ;
assign n21754 =  ( n21753 ) == ( bv_1_0_n53 )  ;
assign n21755 =  ( wr_addr ) == ( bv_8_171_n411 )  ;
assign n21756 =  ( n21754 ) & (n21755 )  ;
assign n21757 =  ( n21756 ) & (wr )  ;
assign n21758 =  ( n21757 ) ? ( bv_8_0_n69 ) : ( iram_171 ) ;
assign n21759 = wr_addr[7:7] ;
assign n21760 =  ( n21759 ) == ( bv_1_0_n53 )  ;
assign n21761 =  ( wr_addr ) == ( bv_8_171_n411 )  ;
assign n21762 =  ( n21760 ) & (n21761 )  ;
assign n21763 =  ( n21762 ) & (wr )  ;
assign n21764 =  ( n21763 ) ? ( n5071 ) : ( iram_171 ) ;
assign n21765 = wr_addr[7:7] ;
assign n21766 =  ( n21765 ) == ( bv_1_0_n53 )  ;
assign n21767 =  ( wr_addr ) == ( bv_8_171_n411 )  ;
assign n21768 =  ( n21766 ) & (n21767 )  ;
assign n21769 =  ( n21768 ) & (wr )  ;
assign n21770 =  ( n21769 ) ? ( n5096 ) : ( iram_171 ) ;
assign n21771 = wr_addr[7:7] ;
assign n21772 =  ( n21771 ) == ( bv_1_0_n53 )  ;
assign n21773 =  ( wr_addr ) == ( bv_8_171_n411 )  ;
assign n21774 =  ( n21772 ) & (n21773 )  ;
assign n21775 =  ( n21774 ) & (wr )  ;
assign n21776 =  ( n21775 ) ? ( n5123 ) : ( iram_171 ) ;
assign n21777 = wr_addr[7:7] ;
assign n21778 =  ( n21777 ) == ( bv_1_0_n53 )  ;
assign n21779 =  ( wr_addr ) == ( bv_8_171_n411 )  ;
assign n21780 =  ( n21778 ) & (n21779 )  ;
assign n21781 =  ( n21780 ) & (wr )  ;
assign n21782 =  ( n21781 ) ? ( n5165 ) : ( iram_171 ) ;
assign n21783 = wr_addr[7:7] ;
assign n21784 =  ( n21783 ) == ( bv_1_0_n53 )  ;
assign n21785 =  ( wr_addr ) == ( bv_8_171_n411 )  ;
assign n21786 =  ( n21784 ) & (n21785 )  ;
assign n21787 =  ( n21786 ) & (wr )  ;
assign n21788 =  ( n21787 ) ? ( n5204 ) : ( iram_171 ) ;
assign n21789 = wr_addr[7:7] ;
assign n21790 =  ( n21789 ) == ( bv_1_0_n53 )  ;
assign n21791 =  ( wr_addr ) == ( bv_8_171_n411 )  ;
assign n21792 =  ( n21790 ) & (n21791 )  ;
assign n21793 =  ( n21792 ) & (wr )  ;
assign n21794 =  ( n21793 ) ? ( n5262 ) : ( iram_171 ) ;
assign n21795 = wr_addr[7:7] ;
assign n21796 =  ( n21795 ) == ( bv_1_0_n53 )  ;
assign n21797 =  ( wr_addr ) == ( bv_8_171_n411 )  ;
assign n21798 =  ( n21796 ) & (n21797 )  ;
assign n21799 =  ( n21798 ) & (wr )  ;
assign n21800 =  ( n21799 ) ? ( n5298 ) : ( iram_171 ) ;
assign n21801 = wr_addr[7:7] ;
assign n21802 =  ( n21801 ) == ( bv_1_0_n53 )  ;
assign n21803 =  ( wr_addr ) == ( bv_8_171_n411 )  ;
assign n21804 =  ( n21802 ) & (n21803 )  ;
assign n21805 =  ( n21804 ) & (wr )  ;
assign n21806 =  ( n21805 ) ? ( n5325 ) : ( iram_171 ) ;
assign n21807 = wr_addr[7:7] ;
assign n21808 =  ( n21807 ) == ( bv_1_0_n53 )  ;
assign n21809 =  ( wr_addr ) == ( bv_8_172_n413 )  ;
assign n21810 =  ( n21808 ) & (n21809 )  ;
assign n21811 =  ( n21810 ) & (wr )  ;
assign n21812 =  ( n21811 ) ? ( n4782 ) : ( iram_172 ) ;
assign n21813 = wr_addr[7:7] ;
assign n21814 =  ( n21813 ) == ( bv_1_0_n53 )  ;
assign n21815 =  ( wr_addr ) == ( bv_8_172_n413 )  ;
assign n21816 =  ( n21814 ) & (n21815 )  ;
assign n21817 =  ( n21816 ) & (wr )  ;
assign n21818 =  ( n21817 ) ? ( n4841 ) : ( iram_172 ) ;
assign n21819 = wr_addr[7:7] ;
assign n21820 =  ( n21819 ) == ( bv_1_0_n53 )  ;
assign n21821 =  ( wr_addr ) == ( bv_8_172_n413 )  ;
assign n21822 =  ( n21820 ) & (n21821 )  ;
assign n21823 =  ( n21822 ) & (wr )  ;
assign n21824 =  ( n21823 ) ? ( n5449 ) : ( iram_172 ) ;
assign n21825 = wr_addr[7:7] ;
assign n21826 =  ( n21825 ) == ( bv_1_0_n53 )  ;
assign n21827 =  ( wr_addr ) == ( bv_8_172_n413 )  ;
assign n21828 =  ( n21826 ) & (n21827 )  ;
assign n21829 =  ( n21828 ) & (wr )  ;
assign n21830 =  ( n21829 ) ? ( n4906 ) : ( iram_172 ) ;
assign n21831 = wr_addr[7:7] ;
assign n21832 =  ( n21831 ) == ( bv_1_0_n53 )  ;
assign n21833 =  ( wr_addr ) == ( bv_8_172_n413 )  ;
assign n21834 =  ( n21832 ) & (n21833 )  ;
assign n21835 =  ( n21834 ) & (wr )  ;
assign n21836 =  ( n21835 ) ? ( n5485 ) : ( iram_172 ) ;
assign n21837 = wr_addr[7:7] ;
assign n21838 =  ( n21837 ) == ( bv_1_0_n53 )  ;
assign n21839 =  ( wr_addr ) == ( bv_8_172_n413 )  ;
assign n21840 =  ( n21838 ) & (n21839 )  ;
assign n21841 =  ( n21840 ) & (wr )  ;
assign n21842 =  ( n21841 ) ? ( n5512 ) : ( iram_172 ) ;
assign n21843 = wr_addr[7:7] ;
assign n21844 =  ( n21843 ) == ( bv_1_0_n53 )  ;
assign n21845 =  ( wr_addr ) == ( bv_8_172_n413 )  ;
assign n21846 =  ( n21844 ) & (n21845 )  ;
assign n21847 =  ( n21846 ) & (wr )  ;
assign n21848 =  ( n21847 ) ? ( bv_8_0_n69 ) : ( iram_172 ) ;
assign n21849 = wr_addr[7:7] ;
assign n21850 =  ( n21849 ) == ( bv_1_0_n53 )  ;
assign n21851 =  ( wr_addr ) == ( bv_8_172_n413 )  ;
assign n21852 =  ( n21850 ) & (n21851 )  ;
assign n21853 =  ( n21852 ) & (wr )  ;
assign n21854 =  ( n21853 ) ? ( n5071 ) : ( iram_172 ) ;
assign n21855 = wr_addr[7:7] ;
assign n21856 =  ( n21855 ) == ( bv_1_0_n53 )  ;
assign n21857 =  ( wr_addr ) == ( bv_8_172_n413 )  ;
assign n21858 =  ( n21856 ) & (n21857 )  ;
assign n21859 =  ( n21858 ) & (wr )  ;
assign n21860 =  ( n21859 ) ? ( n5096 ) : ( iram_172 ) ;
assign n21861 = wr_addr[7:7] ;
assign n21862 =  ( n21861 ) == ( bv_1_0_n53 )  ;
assign n21863 =  ( wr_addr ) == ( bv_8_172_n413 )  ;
assign n21864 =  ( n21862 ) & (n21863 )  ;
assign n21865 =  ( n21864 ) & (wr )  ;
assign n21866 =  ( n21865 ) ? ( n5123 ) : ( iram_172 ) ;
assign n21867 = wr_addr[7:7] ;
assign n21868 =  ( n21867 ) == ( bv_1_0_n53 )  ;
assign n21869 =  ( wr_addr ) == ( bv_8_172_n413 )  ;
assign n21870 =  ( n21868 ) & (n21869 )  ;
assign n21871 =  ( n21870 ) & (wr )  ;
assign n21872 =  ( n21871 ) ? ( n5165 ) : ( iram_172 ) ;
assign n21873 = wr_addr[7:7] ;
assign n21874 =  ( n21873 ) == ( bv_1_0_n53 )  ;
assign n21875 =  ( wr_addr ) == ( bv_8_172_n413 )  ;
assign n21876 =  ( n21874 ) & (n21875 )  ;
assign n21877 =  ( n21876 ) & (wr )  ;
assign n21878 =  ( n21877 ) ? ( n5204 ) : ( iram_172 ) ;
assign n21879 = wr_addr[7:7] ;
assign n21880 =  ( n21879 ) == ( bv_1_0_n53 )  ;
assign n21881 =  ( wr_addr ) == ( bv_8_172_n413 )  ;
assign n21882 =  ( n21880 ) & (n21881 )  ;
assign n21883 =  ( n21882 ) & (wr )  ;
assign n21884 =  ( n21883 ) ? ( n5262 ) : ( iram_172 ) ;
assign n21885 = wr_addr[7:7] ;
assign n21886 =  ( n21885 ) == ( bv_1_0_n53 )  ;
assign n21887 =  ( wr_addr ) == ( bv_8_172_n413 )  ;
assign n21888 =  ( n21886 ) & (n21887 )  ;
assign n21889 =  ( n21888 ) & (wr )  ;
assign n21890 =  ( n21889 ) ? ( n5298 ) : ( iram_172 ) ;
assign n21891 = wr_addr[7:7] ;
assign n21892 =  ( n21891 ) == ( bv_1_0_n53 )  ;
assign n21893 =  ( wr_addr ) == ( bv_8_172_n413 )  ;
assign n21894 =  ( n21892 ) & (n21893 )  ;
assign n21895 =  ( n21894 ) & (wr )  ;
assign n21896 =  ( n21895 ) ? ( n5325 ) : ( iram_172 ) ;
assign n21897 = wr_addr[7:7] ;
assign n21898 =  ( n21897 ) == ( bv_1_0_n53 )  ;
assign n21899 =  ( wr_addr ) == ( bv_8_173_n415 )  ;
assign n21900 =  ( n21898 ) & (n21899 )  ;
assign n21901 =  ( n21900 ) & (wr )  ;
assign n21902 =  ( n21901 ) ? ( n4782 ) : ( iram_173 ) ;
assign n21903 = wr_addr[7:7] ;
assign n21904 =  ( n21903 ) == ( bv_1_0_n53 )  ;
assign n21905 =  ( wr_addr ) == ( bv_8_173_n415 )  ;
assign n21906 =  ( n21904 ) & (n21905 )  ;
assign n21907 =  ( n21906 ) & (wr )  ;
assign n21908 =  ( n21907 ) ? ( n4841 ) : ( iram_173 ) ;
assign n21909 = wr_addr[7:7] ;
assign n21910 =  ( n21909 ) == ( bv_1_0_n53 )  ;
assign n21911 =  ( wr_addr ) == ( bv_8_173_n415 )  ;
assign n21912 =  ( n21910 ) & (n21911 )  ;
assign n21913 =  ( n21912 ) & (wr )  ;
assign n21914 =  ( n21913 ) ? ( n5449 ) : ( iram_173 ) ;
assign n21915 = wr_addr[7:7] ;
assign n21916 =  ( n21915 ) == ( bv_1_0_n53 )  ;
assign n21917 =  ( wr_addr ) == ( bv_8_173_n415 )  ;
assign n21918 =  ( n21916 ) & (n21917 )  ;
assign n21919 =  ( n21918 ) & (wr )  ;
assign n21920 =  ( n21919 ) ? ( n4906 ) : ( iram_173 ) ;
assign n21921 = wr_addr[7:7] ;
assign n21922 =  ( n21921 ) == ( bv_1_0_n53 )  ;
assign n21923 =  ( wr_addr ) == ( bv_8_173_n415 )  ;
assign n21924 =  ( n21922 ) & (n21923 )  ;
assign n21925 =  ( n21924 ) & (wr )  ;
assign n21926 =  ( n21925 ) ? ( n5485 ) : ( iram_173 ) ;
assign n21927 = wr_addr[7:7] ;
assign n21928 =  ( n21927 ) == ( bv_1_0_n53 )  ;
assign n21929 =  ( wr_addr ) == ( bv_8_173_n415 )  ;
assign n21930 =  ( n21928 ) & (n21929 )  ;
assign n21931 =  ( n21930 ) & (wr )  ;
assign n21932 =  ( n21931 ) ? ( n5512 ) : ( iram_173 ) ;
assign n21933 = wr_addr[7:7] ;
assign n21934 =  ( n21933 ) == ( bv_1_0_n53 )  ;
assign n21935 =  ( wr_addr ) == ( bv_8_173_n415 )  ;
assign n21936 =  ( n21934 ) & (n21935 )  ;
assign n21937 =  ( n21936 ) & (wr )  ;
assign n21938 =  ( n21937 ) ? ( bv_8_0_n69 ) : ( iram_173 ) ;
assign n21939 = wr_addr[7:7] ;
assign n21940 =  ( n21939 ) == ( bv_1_0_n53 )  ;
assign n21941 =  ( wr_addr ) == ( bv_8_173_n415 )  ;
assign n21942 =  ( n21940 ) & (n21941 )  ;
assign n21943 =  ( n21942 ) & (wr )  ;
assign n21944 =  ( n21943 ) ? ( n5071 ) : ( iram_173 ) ;
assign n21945 = wr_addr[7:7] ;
assign n21946 =  ( n21945 ) == ( bv_1_0_n53 )  ;
assign n21947 =  ( wr_addr ) == ( bv_8_173_n415 )  ;
assign n21948 =  ( n21946 ) & (n21947 )  ;
assign n21949 =  ( n21948 ) & (wr )  ;
assign n21950 =  ( n21949 ) ? ( n5096 ) : ( iram_173 ) ;
assign n21951 = wr_addr[7:7] ;
assign n21952 =  ( n21951 ) == ( bv_1_0_n53 )  ;
assign n21953 =  ( wr_addr ) == ( bv_8_173_n415 )  ;
assign n21954 =  ( n21952 ) & (n21953 )  ;
assign n21955 =  ( n21954 ) & (wr )  ;
assign n21956 =  ( n21955 ) ? ( n5123 ) : ( iram_173 ) ;
assign n21957 = wr_addr[7:7] ;
assign n21958 =  ( n21957 ) == ( bv_1_0_n53 )  ;
assign n21959 =  ( wr_addr ) == ( bv_8_173_n415 )  ;
assign n21960 =  ( n21958 ) & (n21959 )  ;
assign n21961 =  ( n21960 ) & (wr )  ;
assign n21962 =  ( n21961 ) ? ( n5165 ) : ( iram_173 ) ;
assign n21963 = wr_addr[7:7] ;
assign n21964 =  ( n21963 ) == ( bv_1_0_n53 )  ;
assign n21965 =  ( wr_addr ) == ( bv_8_173_n415 )  ;
assign n21966 =  ( n21964 ) & (n21965 )  ;
assign n21967 =  ( n21966 ) & (wr )  ;
assign n21968 =  ( n21967 ) ? ( n5204 ) : ( iram_173 ) ;
assign n21969 = wr_addr[7:7] ;
assign n21970 =  ( n21969 ) == ( bv_1_0_n53 )  ;
assign n21971 =  ( wr_addr ) == ( bv_8_173_n415 )  ;
assign n21972 =  ( n21970 ) & (n21971 )  ;
assign n21973 =  ( n21972 ) & (wr )  ;
assign n21974 =  ( n21973 ) ? ( n5262 ) : ( iram_173 ) ;
assign n21975 = wr_addr[7:7] ;
assign n21976 =  ( n21975 ) == ( bv_1_0_n53 )  ;
assign n21977 =  ( wr_addr ) == ( bv_8_173_n415 )  ;
assign n21978 =  ( n21976 ) & (n21977 )  ;
assign n21979 =  ( n21978 ) & (wr )  ;
assign n21980 =  ( n21979 ) ? ( n5298 ) : ( iram_173 ) ;
assign n21981 = wr_addr[7:7] ;
assign n21982 =  ( n21981 ) == ( bv_1_0_n53 )  ;
assign n21983 =  ( wr_addr ) == ( bv_8_173_n415 )  ;
assign n21984 =  ( n21982 ) & (n21983 )  ;
assign n21985 =  ( n21984 ) & (wr )  ;
assign n21986 =  ( n21985 ) ? ( n5325 ) : ( iram_173 ) ;
assign n21987 = wr_addr[7:7] ;
assign n21988 =  ( n21987 ) == ( bv_1_0_n53 )  ;
assign n21989 =  ( wr_addr ) == ( bv_8_174_n417 )  ;
assign n21990 =  ( n21988 ) & (n21989 )  ;
assign n21991 =  ( n21990 ) & (wr )  ;
assign n21992 =  ( n21991 ) ? ( n4782 ) : ( iram_174 ) ;
assign n21993 = wr_addr[7:7] ;
assign n21994 =  ( n21993 ) == ( bv_1_0_n53 )  ;
assign n21995 =  ( wr_addr ) == ( bv_8_174_n417 )  ;
assign n21996 =  ( n21994 ) & (n21995 )  ;
assign n21997 =  ( n21996 ) & (wr )  ;
assign n21998 =  ( n21997 ) ? ( n4841 ) : ( iram_174 ) ;
assign n21999 = wr_addr[7:7] ;
assign n22000 =  ( n21999 ) == ( bv_1_0_n53 )  ;
assign n22001 =  ( wr_addr ) == ( bv_8_174_n417 )  ;
assign n22002 =  ( n22000 ) & (n22001 )  ;
assign n22003 =  ( n22002 ) & (wr )  ;
assign n22004 =  ( n22003 ) ? ( n5449 ) : ( iram_174 ) ;
assign n22005 = wr_addr[7:7] ;
assign n22006 =  ( n22005 ) == ( bv_1_0_n53 )  ;
assign n22007 =  ( wr_addr ) == ( bv_8_174_n417 )  ;
assign n22008 =  ( n22006 ) & (n22007 )  ;
assign n22009 =  ( n22008 ) & (wr )  ;
assign n22010 =  ( n22009 ) ? ( n4906 ) : ( iram_174 ) ;
assign n22011 = wr_addr[7:7] ;
assign n22012 =  ( n22011 ) == ( bv_1_0_n53 )  ;
assign n22013 =  ( wr_addr ) == ( bv_8_174_n417 )  ;
assign n22014 =  ( n22012 ) & (n22013 )  ;
assign n22015 =  ( n22014 ) & (wr )  ;
assign n22016 =  ( n22015 ) ? ( n5485 ) : ( iram_174 ) ;
assign n22017 = wr_addr[7:7] ;
assign n22018 =  ( n22017 ) == ( bv_1_0_n53 )  ;
assign n22019 =  ( wr_addr ) == ( bv_8_174_n417 )  ;
assign n22020 =  ( n22018 ) & (n22019 )  ;
assign n22021 =  ( n22020 ) & (wr )  ;
assign n22022 =  ( n22021 ) ? ( n5512 ) : ( iram_174 ) ;
assign n22023 = wr_addr[7:7] ;
assign n22024 =  ( n22023 ) == ( bv_1_0_n53 )  ;
assign n22025 =  ( wr_addr ) == ( bv_8_174_n417 )  ;
assign n22026 =  ( n22024 ) & (n22025 )  ;
assign n22027 =  ( n22026 ) & (wr )  ;
assign n22028 =  ( n22027 ) ? ( bv_8_0_n69 ) : ( iram_174 ) ;
assign n22029 = wr_addr[7:7] ;
assign n22030 =  ( n22029 ) == ( bv_1_0_n53 )  ;
assign n22031 =  ( wr_addr ) == ( bv_8_174_n417 )  ;
assign n22032 =  ( n22030 ) & (n22031 )  ;
assign n22033 =  ( n22032 ) & (wr )  ;
assign n22034 =  ( n22033 ) ? ( n5071 ) : ( iram_174 ) ;
assign n22035 = wr_addr[7:7] ;
assign n22036 =  ( n22035 ) == ( bv_1_0_n53 )  ;
assign n22037 =  ( wr_addr ) == ( bv_8_174_n417 )  ;
assign n22038 =  ( n22036 ) & (n22037 )  ;
assign n22039 =  ( n22038 ) & (wr )  ;
assign n22040 =  ( n22039 ) ? ( n5096 ) : ( iram_174 ) ;
assign n22041 = wr_addr[7:7] ;
assign n22042 =  ( n22041 ) == ( bv_1_0_n53 )  ;
assign n22043 =  ( wr_addr ) == ( bv_8_174_n417 )  ;
assign n22044 =  ( n22042 ) & (n22043 )  ;
assign n22045 =  ( n22044 ) & (wr )  ;
assign n22046 =  ( n22045 ) ? ( n5123 ) : ( iram_174 ) ;
assign n22047 = wr_addr[7:7] ;
assign n22048 =  ( n22047 ) == ( bv_1_0_n53 )  ;
assign n22049 =  ( wr_addr ) == ( bv_8_174_n417 )  ;
assign n22050 =  ( n22048 ) & (n22049 )  ;
assign n22051 =  ( n22050 ) & (wr )  ;
assign n22052 =  ( n22051 ) ? ( n5165 ) : ( iram_174 ) ;
assign n22053 = wr_addr[7:7] ;
assign n22054 =  ( n22053 ) == ( bv_1_0_n53 )  ;
assign n22055 =  ( wr_addr ) == ( bv_8_174_n417 )  ;
assign n22056 =  ( n22054 ) & (n22055 )  ;
assign n22057 =  ( n22056 ) & (wr )  ;
assign n22058 =  ( n22057 ) ? ( n5204 ) : ( iram_174 ) ;
assign n22059 = wr_addr[7:7] ;
assign n22060 =  ( n22059 ) == ( bv_1_0_n53 )  ;
assign n22061 =  ( wr_addr ) == ( bv_8_174_n417 )  ;
assign n22062 =  ( n22060 ) & (n22061 )  ;
assign n22063 =  ( n22062 ) & (wr )  ;
assign n22064 =  ( n22063 ) ? ( n5262 ) : ( iram_174 ) ;
assign n22065 = wr_addr[7:7] ;
assign n22066 =  ( n22065 ) == ( bv_1_0_n53 )  ;
assign n22067 =  ( wr_addr ) == ( bv_8_174_n417 )  ;
assign n22068 =  ( n22066 ) & (n22067 )  ;
assign n22069 =  ( n22068 ) & (wr )  ;
assign n22070 =  ( n22069 ) ? ( n5298 ) : ( iram_174 ) ;
assign n22071 = wr_addr[7:7] ;
assign n22072 =  ( n22071 ) == ( bv_1_0_n53 )  ;
assign n22073 =  ( wr_addr ) == ( bv_8_174_n417 )  ;
assign n22074 =  ( n22072 ) & (n22073 )  ;
assign n22075 =  ( n22074 ) & (wr )  ;
assign n22076 =  ( n22075 ) ? ( n5325 ) : ( iram_174 ) ;
assign n22077 = wr_addr[7:7] ;
assign n22078 =  ( n22077 ) == ( bv_1_0_n53 )  ;
assign n22079 =  ( wr_addr ) == ( bv_8_175_n419 )  ;
assign n22080 =  ( n22078 ) & (n22079 )  ;
assign n22081 =  ( n22080 ) & (wr )  ;
assign n22082 =  ( n22081 ) ? ( n4782 ) : ( iram_175 ) ;
assign n22083 = wr_addr[7:7] ;
assign n22084 =  ( n22083 ) == ( bv_1_0_n53 )  ;
assign n22085 =  ( wr_addr ) == ( bv_8_175_n419 )  ;
assign n22086 =  ( n22084 ) & (n22085 )  ;
assign n22087 =  ( n22086 ) & (wr )  ;
assign n22088 =  ( n22087 ) ? ( n4841 ) : ( iram_175 ) ;
assign n22089 = wr_addr[7:7] ;
assign n22090 =  ( n22089 ) == ( bv_1_0_n53 )  ;
assign n22091 =  ( wr_addr ) == ( bv_8_175_n419 )  ;
assign n22092 =  ( n22090 ) & (n22091 )  ;
assign n22093 =  ( n22092 ) & (wr )  ;
assign n22094 =  ( n22093 ) ? ( n5449 ) : ( iram_175 ) ;
assign n22095 = wr_addr[7:7] ;
assign n22096 =  ( n22095 ) == ( bv_1_0_n53 )  ;
assign n22097 =  ( wr_addr ) == ( bv_8_175_n419 )  ;
assign n22098 =  ( n22096 ) & (n22097 )  ;
assign n22099 =  ( n22098 ) & (wr )  ;
assign n22100 =  ( n22099 ) ? ( n4906 ) : ( iram_175 ) ;
assign n22101 = wr_addr[7:7] ;
assign n22102 =  ( n22101 ) == ( bv_1_0_n53 )  ;
assign n22103 =  ( wr_addr ) == ( bv_8_175_n419 )  ;
assign n22104 =  ( n22102 ) & (n22103 )  ;
assign n22105 =  ( n22104 ) & (wr )  ;
assign n22106 =  ( n22105 ) ? ( n5485 ) : ( iram_175 ) ;
assign n22107 = wr_addr[7:7] ;
assign n22108 =  ( n22107 ) == ( bv_1_0_n53 )  ;
assign n22109 =  ( wr_addr ) == ( bv_8_175_n419 )  ;
assign n22110 =  ( n22108 ) & (n22109 )  ;
assign n22111 =  ( n22110 ) & (wr )  ;
assign n22112 =  ( n22111 ) ? ( n5512 ) : ( iram_175 ) ;
assign n22113 = wr_addr[7:7] ;
assign n22114 =  ( n22113 ) == ( bv_1_0_n53 )  ;
assign n22115 =  ( wr_addr ) == ( bv_8_175_n419 )  ;
assign n22116 =  ( n22114 ) & (n22115 )  ;
assign n22117 =  ( n22116 ) & (wr )  ;
assign n22118 =  ( n22117 ) ? ( bv_8_0_n69 ) : ( iram_175 ) ;
assign n22119 = wr_addr[7:7] ;
assign n22120 =  ( n22119 ) == ( bv_1_0_n53 )  ;
assign n22121 =  ( wr_addr ) == ( bv_8_175_n419 )  ;
assign n22122 =  ( n22120 ) & (n22121 )  ;
assign n22123 =  ( n22122 ) & (wr )  ;
assign n22124 =  ( n22123 ) ? ( n5071 ) : ( iram_175 ) ;
assign n22125 = wr_addr[7:7] ;
assign n22126 =  ( n22125 ) == ( bv_1_0_n53 )  ;
assign n22127 =  ( wr_addr ) == ( bv_8_175_n419 )  ;
assign n22128 =  ( n22126 ) & (n22127 )  ;
assign n22129 =  ( n22128 ) & (wr )  ;
assign n22130 =  ( n22129 ) ? ( n5096 ) : ( iram_175 ) ;
assign n22131 = wr_addr[7:7] ;
assign n22132 =  ( n22131 ) == ( bv_1_0_n53 )  ;
assign n22133 =  ( wr_addr ) == ( bv_8_175_n419 )  ;
assign n22134 =  ( n22132 ) & (n22133 )  ;
assign n22135 =  ( n22134 ) & (wr )  ;
assign n22136 =  ( n22135 ) ? ( n5123 ) : ( iram_175 ) ;
assign n22137 = wr_addr[7:7] ;
assign n22138 =  ( n22137 ) == ( bv_1_0_n53 )  ;
assign n22139 =  ( wr_addr ) == ( bv_8_175_n419 )  ;
assign n22140 =  ( n22138 ) & (n22139 )  ;
assign n22141 =  ( n22140 ) & (wr )  ;
assign n22142 =  ( n22141 ) ? ( n5165 ) : ( iram_175 ) ;
assign n22143 = wr_addr[7:7] ;
assign n22144 =  ( n22143 ) == ( bv_1_0_n53 )  ;
assign n22145 =  ( wr_addr ) == ( bv_8_175_n419 )  ;
assign n22146 =  ( n22144 ) & (n22145 )  ;
assign n22147 =  ( n22146 ) & (wr )  ;
assign n22148 =  ( n22147 ) ? ( n5204 ) : ( iram_175 ) ;
assign n22149 = wr_addr[7:7] ;
assign n22150 =  ( n22149 ) == ( bv_1_0_n53 )  ;
assign n22151 =  ( wr_addr ) == ( bv_8_175_n419 )  ;
assign n22152 =  ( n22150 ) & (n22151 )  ;
assign n22153 =  ( n22152 ) & (wr )  ;
assign n22154 =  ( n22153 ) ? ( n5262 ) : ( iram_175 ) ;
assign n22155 = wr_addr[7:7] ;
assign n22156 =  ( n22155 ) == ( bv_1_0_n53 )  ;
assign n22157 =  ( wr_addr ) == ( bv_8_175_n419 )  ;
assign n22158 =  ( n22156 ) & (n22157 )  ;
assign n22159 =  ( n22158 ) & (wr )  ;
assign n22160 =  ( n22159 ) ? ( n5298 ) : ( iram_175 ) ;
assign n22161 = wr_addr[7:7] ;
assign n22162 =  ( n22161 ) == ( bv_1_0_n53 )  ;
assign n22163 =  ( wr_addr ) == ( bv_8_175_n419 )  ;
assign n22164 =  ( n22162 ) & (n22163 )  ;
assign n22165 =  ( n22164 ) & (wr )  ;
assign n22166 =  ( n22165 ) ? ( n5325 ) : ( iram_175 ) ;
assign n22167 = wr_addr[7:7] ;
assign n22168 =  ( n22167 ) == ( bv_1_0_n53 )  ;
assign n22169 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n22170 =  ( n22168 ) & (n22169 )  ;
assign n22171 =  ( n22170 ) & (wr )  ;
assign n22172 =  ( n22171 ) ? ( n4782 ) : ( iram_176 ) ;
assign n22173 = wr_addr[7:7] ;
assign n22174 =  ( n22173 ) == ( bv_1_0_n53 )  ;
assign n22175 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n22176 =  ( n22174 ) & (n22175 )  ;
assign n22177 =  ( n22176 ) & (wr )  ;
assign n22178 =  ( n22177 ) ? ( n4841 ) : ( iram_176 ) ;
assign n22179 = wr_addr[7:7] ;
assign n22180 =  ( n22179 ) == ( bv_1_0_n53 )  ;
assign n22181 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n22182 =  ( n22180 ) & (n22181 )  ;
assign n22183 =  ( n22182 ) & (wr )  ;
assign n22184 =  ( n22183 ) ? ( n5449 ) : ( iram_176 ) ;
assign n22185 = wr_addr[7:7] ;
assign n22186 =  ( n22185 ) == ( bv_1_0_n53 )  ;
assign n22187 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n22188 =  ( n22186 ) & (n22187 )  ;
assign n22189 =  ( n22188 ) & (wr )  ;
assign n22190 =  ( n22189 ) ? ( n4906 ) : ( iram_176 ) ;
assign n22191 = wr_addr[7:7] ;
assign n22192 =  ( n22191 ) == ( bv_1_0_n53 )  ;
assign n22193 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n22194 =  ( n22192 ) & (n22193 )  ;
assign n22195 =  ( n22194 ) & (wr )  ;
assign n22196 =  ( n22195 ) ? ( n5485 ) : ( iram_176 ) ;
assign n22197 = wr_addr[7:7] ;
assign n22198 =  ( n22197 ) == ( bv_1_0_n53 )  ;
assign n22199 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n22200 =  ( n22198 ) & (n22199 )  ;
assign n22201 =  ( n22200 ) & (wr )  ;
assign n22202 =  ( n22201 ) ? ( n5512 ) : ( iram_176 ) ;
assign n22203 = wr_addr[7:7] ;
assign n22204 =  ( n22203 ) == ( bv_1_0_n53 )  ;
assign n22205 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n22206 =  ( n22204 ) & (n22205 )  ;
assign n22207 =  ( n22206 ) & (wr )  ;
assign n22208 =  ( n22207 ) ? ( bv_8_0_n69 ) : ( iram_176 ) ;
assign n22209 = wr_addr[7:7] ;
assign n22210 =  ( n22209 ) == ( bv_1_0_n53 )  ;
assign n22211 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n22212 =  ( n22210 ) & (n22211 )  ;
assign n22213 =  ( n22212 ) & (wr )  ;
assign n22214 =  ( n22213 ) ? ( n5071 ) : ( iram_176 ) ;
assign n22215 = wr_addr[7:7] ;
assign n22216 =  ( n22215 ) == ( bv_1_0_n53 )  ;
assign n22217 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n22218 =  ( n22216 ) & (n22217 )  ;
assign n22219 =  ( n22218 ) & (wr )  ;
assign n22220 =  ( n22219 ) ? ( n5096 ) : ( iram_176 ) ;
assign n22221 = wr_addr[7:7] ;
assign n22222 =  ( n22221 ) == ( bv_1_0_n53 )  ;
assign n22223 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n22224 =  ( n22222 ) & (n22223 )  ;
assign n22225 =  ( n22224 ) & (wr )  ;
assign n22226 =  ( n22225 ) ? ( n5123 ) : ( iram_176 ) ;
assign n22227 = wr_addr[7:7] ;
assign n22228 =  ( n22227 ) == ( bv_1_0_n53 )  ;
assign n22229 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n22230 =  ( n22228 ) & (n22229 )  ;
assign n22231 =  ( n22230 ) & (wr )  ;
assign n22232 =  ( n22231 ) ? ( n5165 ) : ( iram_176 ) ;
assign n22233 = wr_addr[7:7] ;
assign n22234 =  ( n22233 ) == ( bv_1_0_n53 )  ;
assign n22235 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n22236 =  ( n22234 ) & (n22235 )  ;
assign n22237 =  ( n22236 ) & (wr )  ;
assign n22238 =  ( n22237 ) ? ( n5204 ) : ( iram_176 ) ;
assign n22239 = wr_addr[7:7] ;
assign n22240 =  ( n22239 ) == ( bv_1_0_n53 )  ;
assign n22241 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n22242 =  ( n22240 ) & (n22241 )  ;
assign n22243 =  ( n22242 ) & (wr )  ;
assign n22244 =  ( n22243 ) ? ( n5262 ) : ( iram_176 ) ;
assign n22245 = wr_addr[7:7] ;
assign n22246 =  ( n22245 ) == ( bv_1_0_n53 )  ;
assign n22247 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n22248 =  ( n22246 ) & (n22247 )  ;
assign n22249 =  ( n22248 ) & (wr )  ;
assign n22250 =  ( n22249 ) ? ( n5298 ) : ( iram_176 ) ;
assign n22251 = wr_addr[7:7] ;
assign n22252 =  ( n22251 ) == ( bv_1_0_n53 )  ;
assign n22253 =  ( wr_addr ) == ( bv_8_176_n421 )  ;
assign n22254 =  ( n22252 ) & (n22253 )  ;
assign n22255 =  ( n22254 ) & (wr )  ;
assign n22256 =  ( n22255 ) ? ( n5325 ) : ( iram_176 ) ;
assign n22257 = wr_addr[7:7] ;
assign n22258 =  ( n22257 ) == ( bv_1_0_n53 )  ;
assign n22259 =  ( wr_addr ) == ( bv_8_177_n423 )  ;
assign n22260 =  ( n22258 ) & (n22259 )  ;
assign n22261 =  ( n22260 ) & (wr )  ;
assign n22262 =  ( n22261 ) ? ( n4782 ) : ( iram_177 ) ;
assign n22263 = wr_addr[7:7] ;
assign n22264 =  ( n22263 ) == ( bv_1_0_n53 )  ;
assign n22265 =  ( wr_addr ) == ( bv_8_177_n423 )  ;
assign n22266 =  ( n22264 ) & (n22265 )  ;
assign n22267 =  ( n22266 ) & (wr )  ;
assign n22268 =  ( n22267 ) ? ( n4841 ) : ( iram_177 ) ;
assign n22269 = wr_addr[7:7] ;
assign n22270 =  ( n22269 ) == ( bv_1_0_n53 )  ;
assign n22271 =  ( wr_addr ) == ( bv_8_177_n423 )  ;
assign n22272 =  ( n22270 ) & (n22271 )  ;
assign n22273 =  ( n22272 ) & (wr )  ;
assign n22274 =  ( n22273 ) ? ( n5449 ) : ( iram_177 ) ;
assign n22275 = wr_addr[7:7] ;
assign n22276 =  ( n22275 ) == ( bv_1_0_n53 )  ;
assign n22277 =  ( wr_addr ) == ( bv_8_177_n423 )  ;
assign n22278 =  ( n22276 ) & (n22277 )  ;
assign n22279 =  ( n22278 ) & (wr )  ;
assign n22280 =  ( n22279 ) ? ( n4906 ) : ( iram_177 ) ;
assign n22281 = wr_addr[7:7] ;
assign n22282 =  ( n22281 ) == ( bv_1_0_n53 )  ;
assign n22283 =  ( wr_addr ) == ( bv_8_177_n423 )  ;
assign n22284 =  ( n22282 ) & (n22283 )  ;
assign n22285 =  ( n22284 ) & (wr )  ;
assign n22286 =  ( n22285 ) ? ( n5485 ) : ( iram_177 ) ;
assign n22287 = wr_addr[7:7] ;
assign n22288 =  ( n22287 ) == ( bv_1_0_n53 )  ;
assign n22289 =  ( wr_addr ) == ( bv_8_177_n423 )  ;
assign n22290 =  ( n22288 ) & (n22289 )  ;
assign n22291 =  ( n22290 ) & (wr )  ;
assign n22292 =  ( n22291 ) ? ( n5512 ) : ( iram_177 ) ;
assign n22293 = wr_addr[7:7] ;
assign n22294 =  ( n22293 ) == ( bv_1_0_n53 )  ;
assign n22295 =  ( wr_addr ) == ( bv_8_177_n423 )  ;
assign n22296 =  ( n22294 ) & (n22295 )  ;
assign n22297 =  ( n22296 ) & (wr )  ;
assign n22298 =  ( n22297 ) ? ( bv_8_0_n69 ) : ( iram_177 ) ;
assign n22299 = wr_addr[7:7] ;
assign n22300 =  ( n22299 ) == ( bv_1_0_n53 )  ;
assign n22301 =  ( wr_addr ) == ( bv_8_177_n423 )  ;
assign n22302 =  ( n22300 ) & (n22301 )  ;
assign n22303 =  ( n22302 ) & (wr )  ;
assign n22304 =  ( n22303 ) ? ( n5071 ) : ( iram_177 ) ;
assign n22305 = wr_addr[7:7] ;
assign n22306 =  ( n22305 ) == ( bv_1_0_n53 )  ;
assign n22307 =  ( wr_addr ) == ( bv_8_177_n423 )  ;
assign n22308 =  ( n22306 ) & (n22307 )  ;
assign n22309 =  ( n22308 ) & (wr )  ;
assign n22310 =  ( n22309 ) ? ( n5096 ) : ( iram_177 ) ;
assign n22311 = wr_addr[7:7] ;
assign n22312 =  ( n22311 ) == ( bv_1_0_n53 )  ;
assign n22313 =  ( wr_addr ) == ( bv_8_177_n423 )  ;
assign n22314 =  ( n22312 ) & (n22313 )  ;
assign n22315 =  ( n22314 ) & (wr )  ;
assign n22316 =  ( n22315 ) ? ( n5123 ) : ( iram_177 ) ;
assign n22317 = wr_addr[7:7] ;
assign n22318 =  ( n22317 ) == ( bv_1_0_n53 )  ;
assign n22319 =  ( wr_addr ) == ( bv_8_177_n423 )  ;
assign n22320 =  ( n22318 ) & (n22319 )  ;
assign n22321 =  ( n22320 ) & (wr )  ;
assign n22322 =  ( n22321 ) ? ( n5165 ) : ( iram_177 ) ;
assign n22323 = wr_addr[7:7] ;
assign n22324 =  ( n22323 ) == ( bv_1_0_n53 )  ;
assign n22325 =  ( wr_addr ) == ( bv_8_177_n423 )  ;
assign n22326 =  ( n22324 ) & (n22325 )  ;
assign n22327 =  ( n22326 ) & (wr )  ;
assign n22328 =  ( n22327 ) ? ( n5204 ) : ( iram_177 ) ;
assign n22329 = wr_addr[7:7] ;
assign n22330 =  ( n22329 ) == ( bv_1_0_n53 )  ;
assign n22331 =  ( wr_addr ) == ( bv_8_177_n423 )  ;
assign n22332 =  ( n22330 ) & (n22331 )  ;
assign n22333 =  ( n22332 ) & (wr )  ;
assign n22334 =  ( n22333 ) ? ( n5262 ) : ( iram_177 ) ;
assign n22335 = wr_addr[7:7] ;
assign n22336 =  ( n22335 ) == ( bv_1_0_n53 )  ;
assign n22337 =  ( wr_addr ) == ( bv_8_177_n423 )  ;
assign n22338 =  ( n22336 ) & (n22337 )  ;
assign n22339 =  ( n22338 ) & (wr )  ;
assign n22340 =  ( n22339 ) ? ( n5298 ) : ( iram_177 ) ;
assign n22341 = wr_addr[7:7] ;
assign n22342 =  ( n22341 ) == ( bv_1_0_n53 )  ;
assign n22343 =  ( wr_addr ) == ( bv_8_177_n423 )  ;
assign n22344 =  ( n22342 ) & (n22343 )  ;
assign n22345 =  ( n22344 ) & (wr )  ;
assign n22346 =  ( n22345 ) ? ( n5325 ) : ( iram_177 ) ;
assign n22347 = wr_addr[7:7] ;
assign n22348 =  ( n22347 ) == ( bv_1_0_n53 )  ;
assign n22349 =  ( wr_addr ) == ( bv_8_178_n425 )  ;
assign n22350 =  ( n22348 ) & (n22349 )  ;
assign n22351 =  ( n22350 ) & (wr )  ;
assign n22352 =  ( n22351 ) ? ( n4782 ) : ( iram_178 ) ;
assign n22353 = wr_addr[7:7] ;
assign n22354 =  ( n22353 ) == ( bv_1_0_n53 )  ;
assign n22355 =  ( wr_addr ) == ( bv_8_178_n425 )  ;
assign n22356 =  ( n22354 ) & (n22355 )  ;
assign n22357 =  ( n22356 ) & (wr )  ;
assign n22358 =  ( n22357 ) ? ( n4841 ) : ( iram_178 ) ;
assign n22359 = wr_addr[7:7] ;
assign n22360 =  ( n22359 ) == ( bv_1_0_n53 )  ;
assign n22361 =  ( wr_addr ) == ( bv_8_178_n425 )  ;
assign n22362 =  ( n22360 ) & (n22361 )  ;
assign n22363 =  ( n22362 ) & (wr )  ;
assign n22364 =  ( n22363 ) ? ( n5449 ) : ( iram_178 ) ;
assign n22365 = wr_addr[7:7] ;
assign n22366 =  ( n22365 ) == ( bv_1_0_n53 )  ;
assign n22367 =  ( wr_addr ) == ( bv_8_178_n425 )  ;
assign n22368 =  ( n22366 ) & (n22367 )  ;
assign n22369 =  ( n22368 ) & (wr )  ;
assign n22370 =  ( n22369 ) ? ( n4906 ) : ( iram_178 ) ;
assign n22371 = wr_addr[7:7] ;
assign n22372 =  ( n22371 ) == ( bv_1_0_n53 )  ;
assign n22373 =  ( wr_addr ) == ( bv_8_178_n425 )  ;
assign n22374 =  ( n22372 ) & (n22373 )  ;
assign n22375 =  ( n22374 ) & (wr )  ;
assign n22376 =  ( n22375 ) ? ( n5485 ) : ( iram_178 ) ;
assign n22377 = wr_addr[7:7] ;
assign n22378 =  ( n22377 ) == ( bv_1_0_n53 )  ;
assign n22379 =  ( wr_addr ) == ( bv_8_178_n425 )  ;
assign n22380 =  ( n22378 ) & (n22379 )  ;
assign n22381 =  ( n22380 ) & (wr )  ;
assign n22382 =  ( n22381 ) ? ( n5512 ) : ( iram_178 ) ;
assign n22383 = wr_addr[7:7] ;
assign n22384 =  ( n22383 ) == ( bv_1_0_n53 )  ;
assign n22385 =  ( wr_addr ) == ( bv_8_178_n425 )  ;
assign n22386 =  ( n22384 ) & (n22385 )  ;
assign n22387 =  ( n22386 ) & (wr )  ;
assign n22388 =  ( n22387 ) ? ( bv_8_0_n69 ) : ( iram_178 ) ;
assign n22389 = wr_addr[7:7] ;
assign n22390 =  ( n22389 ) == ( bv_1_0_n53 )  ;
assign n22391 =  ( wr_addr ) == ( bv_8_178_n425 )  ;
assign n22392 =  ( n22390 ) & (n22391 )  ;
assign n22393 =  ( n22392 ) & (wr )  ;
assign n22394 =  ( n22393 ) ? ( n5071 ) : ( iram_178 ) ;
assign n22395 = wr_addr[7:7] ;
assign n22396 =  ( n22395 ) == ( bv_1_0_n53 )  ;
assign n22397 =  ( wr_addr ) == ( bv_8_178_n425 )  ;
assign n22398 =  ( n22396 ) & (n22397 )  ;
assign n22399 =  ( n22398 ) & (wr )  ;
assign n22400 =  ( n22399 ) ? ( n5096 ) : ( iram_178 ) ;
assign n22401 = wr_addr[7:7] ;
assign n22402 =  ( n22401 ) == ( bv_1_0_n53 )  ;
assign n22403 =  ( wr_addr ) == ( bv_8_178_n425 )  ;
assign n22404 =  ( n22402 ) & (n22403 )  ;
assign n22405 =  ( n22404 ) & (wr )  ;
assign n22406 =  ( n22405 ) ? ( n5123 ) : ( iram_178 ) ;
assign n22407 = wr_addr[7:7] ;
assign n22408 =  ( n22407 ) == ( bv_1_0_n53 )  ;
assign n22409 =  ( wr_addr ) == ( bv_8_178_n425 )  ;
assign n22410 =  ( n22408 ) & (n22409 )  ;
assign n22411 =  ( n22410 ) & (wr )  ;
assign n22412 =  ( n22411 ) ? ( n5165 ) : ( iram_178 ) ;
assign n22413 = wr_addr[7:7] ;
assign n22414 =  ( n22413 ) == ( bv_1_0_n53 )  ;
assign n22415 =  ( wr_addr ) == ( bv_8_178_n425 )  ;
assign n22416 =  ( n22414 ) & (n22415 )  ;
assign n22417 =  ( n22416 ) & (wr )  ;
assign n22418 =  ( n22417 ) ? ( n5204 ) : ( iram_178 ) ;
assign n22419 = wr_addr[7:7] ;
assign n22420 =  ( n22419 ) == ( bv_1_0_n53 )  ;
assign n22421 =  ( wr_addr ) == ( bv_8_178_n425 )  ;
assign n22422 =  ( n22420 ) & (n22421 )  ;
assign n22423 =  ( n22422 ) & (wr )  ;
assign n22424 =  ( n22423 ) ? ( n5262 ) : ( iram_178 ) ;
assign n22425 = wr_addr[7:7] ;
assign n22426 =  ( n22425 ) == ( bv_1_0_n53 )  ;
assign n22427 =  ( wr_addr ) == ( bv_8_178_n425 )  ;
assign n22428 =  ( n22426 ) & (n22427 )  ;
assign n22429 =  ( n22428 ) & (wr )  ;
assign n22430 =  ( n22429 ) ? ( n5298 ) : ( iram_178 ) ;
assign n22431 = wr_addr[7:7] ;
assign n22432 =  ( n22431 ) == ( bv_1_0_n53 )  ;
assign n22433 =  ( wr_addr ) == ( bv_8_178_n425 )  ;
assign n22434 =  ( n22432 ) & (n22433 )  ;
assign n22435 =  ( n22434 ) & (wr )  ;
assign n22436 =  ( n22435 ) ? ( n5325 ) : ( iram_178 ) ;
assign n22437 = wr_addr[7:7] ;
assign n22438 =  ( n22437 ) == ( bv_1_0_n53 )  ;
assign n22439 =  ( wr_addr ) == ( bv_8_179_n427 )  ;
assign n22440 =  ( n22438 ) & (n22439 )  ;
assign n22441 =  ( n22440 ) & (wr )  ;
assign n22442 =  ( n22441 ) ? ( n4782 ) : ( iram_179 ) ;
assign n22443 = wr_addr[7:7] ;
assign n22444 =  ( n22443 ) == ( bv_1_0_n53 )  ;
assign n22445 =  ( wr_addr ) == ( bv_8_179_n427 )  ;
assign n22446 =  ( n22444 ) & (n22445 )  ;
assign n22447 =  ( n22446 ) & (wr )  ;
assign n22448 =  ( n22447 ) ? ( n4841 ) : ( iram_179 ) ;
assign n22449 = wr_addr[7:7] ;
assign n22450 =  ( n22449 ) == ( bv_1_0_n53 )  ;
assign n22451 =  ( wr_addr ) == ( bv_8_179_n427 )  ;
assign n22452 =  ( n22450 ) & (n22451 )  ;
assign n22453 =  ( n22452 ) & (wr )  ;
assign n22454 =  ( n22453 ) ? ( n5449 ) : ( iram_179 ) ;
assign n22455 = wr_addr[7:7] ;
assign n22456 =  ( n22455 ) == ( bv_1_0_n53 )  ;
assign n22457 =  ( wr_addr ) == ( bv_8_179_n427 )  ;
assign n22458 =  ( n22456 ) & (n22457 )  ;
assign n22459 =  ( n22458 ) & (wr )  ;
assign n22460 =  ( n22459 ) ? ( n4906 ) : ( iram_179 ) ;
assign n22461 = wr_addr[7:7] ;
assign n22462 =  ( n22461 ) == ( bv_1_0_n53 )  ;
assign n22463 =  ( wr_addr ) == ( bv_8_179_n427 )  ;
assign n22464 =  ( n22462 ) & (n22463 )  ;
assign n22465 =  ( n22464 ) & (wr )  ;
assign n22466 =  ( n22465 ) ? ( n5485 ) : ( iram_179 ) ;
assign n22467 = wr_addr[7:7] ;
assign n22468 =  ( n22467 ) == ( bv_1_0_n53 )  ;
assign n22469 =  ( wr_addr ) == ( bv_8_179_n427 )  ;
assign n22470 =  ( n22468 ) & (n22469 )  ;
assign n22471 =  ( n22470 ) & (wr )  ;
assign n22472 =  ( n22471 ) ? ( n5512 ) : ( iram_179 ) ;
assign n22473 = wr_addr[7:7] ;
assign n22474 =  ( n22473 ) == ( bv_1_0_n53 )  ;
assign n22475 =  ( wr_addr ) == ( bv_8_179_n427 )  ;
assign n22476 =  ( n22474 ) & (n22475 )  ;
assign n22477 =  ( n22476 ) & (wr )  ;
assign n22478 =  ( n22477 ) ? ( bv_8_0_n69 ) : ( iram_179 ) ;
assign n22479 = wr_addr[7:7] ;
assign n22480 =  ( n22479 ) == ( bv_1_0_n53 )  ;
assign n22481 =  ( wr_addr ) == ( bv_8_179_n427 )  ;
assign n22482 =  ( n22480 ) & (n22481 )  ;
assign n22483 =  ( n22482 ) & (wr )  ;
assign n22484 =  ( n22483 ) ? ( n5071 ) : ( iram_179 ) ;
assign n22485 = wr_addr[7:7] ;
assign n22486 =  ( n22485 ) == ( bv_1_0_n53 )  ;
assign n22487 =  ( wr_addr ) == ( bv_8_179_n427 )  ;
assign n22488 =  ( n22486 ) & (n22487 )  ;
assign n22489 =  ( n22488 ) & (wr )  ;
assign n22490 =  ( n22489 ) ? ( n5096 ) : ( iram_179 ) ;
assign n22491 = wr_addr[7:7] ;
assign n22492 =  ( n22491 ) == ( bv_1_0_n53 )  ;
assign n22493 =  ( wr_addr ) == ( bv_8_179_n427 )  ;
assign n22494 =  ( n22492 ) & (n22493 )  ;
assign n22495 =  ( n22494 ) & (wr )  ;
assign n22496 =  ( n22495 ) ? ( n5123 ) : ( iram_179 ) ;
assign n22497 = wr_addr[7:7] ;
assign n22498 =  ( n22497 ) == ( bv_1_0_n53 )  ;
assign n22499 =  ( wr_addr ) == ( bv_8_179_n427 )  ;
assign n22500 =  ( n22498 ) & (n22499 )  ;
assign n22501 =  ( n22500 ) & (wr )  ;
assign n22502 =  ( n22501 ) ? ( n5165 ) : ( iram_179 ) ;
assign n22503 = wr_addr[7:7] ;
assign n22504 =  ( n22503 ) == ( bv_1_0_n53 )  ;
assign n22505 =  ( wr_addr ) == ( bv_8_179_n427 )  ;
assign n22506 =  ( n22504 ) & (n22505 )  ;
assign n22507 =  ( n22506 ) & (wr )  ;
assign n22508 =  ( n22507 ) ? ( n5204 ) : ( iram_179 ) ;
assign n22509 = wr_addr[7:7] ;
assign n22510 =  ( n22509 ) == ( bv_1_0_n53 )  ;
assign n22511 =  ( wr_addr ) == ( bv_8_179_n427 )  ;
assign n22512 =  ( n22510 ) & (n22511 )  ;
assign n22513 =  ( n22512 ) & (wr )  ;
assign n22514 =  ( n22513 ) ? ( n5262 ) : ( iram_179 ) ;
assign n22515 = wr_addr[7:7] ;
assign n22516 =  ( n22515 ) == ( bv_1_0_n53 )  ;
assign n22517 =  ( wr_addr ) == ( bv_8_179_n427 )  ;
assign n22518 =  ( n22516 ) & (n22517 )  ;
assign n22519 =  ( n22518 ) & (wr )  ;
assign n22520 =  ( n22519 ) ? ( n5298 ) : ( iram_179 ) ;
assign n22521 = wr_addr[7:7] ;
assign n22522 =  ( n22521 ) == ( bv_1_0_n53 )  ;
assign n22523 =  ( wr_addr ) == ( bv_8_179_n427 )  ;
assign n22524 =  ( n22522 ) & (n22523 )  ;
assign n22525 =  ( n22524 ) & (wr )  ;
assign n22526 =  ( n22525 ) ? ( n5325 ) : ( iram_179 ) ;
assign n22527 = wr_addr[7:7] ;
assign n22528 =  ( n22527 ) == ( bv_1_0_n53 )  ;
assign n22529 =  ( wr_addr ) == ( bv_8_180_n429 )  ;
assign n22530 =  ( n22528 ) & (n22529 )  ;
assign n22531 =  ( n22530 ) & (wr )  ;
assign n22532 =  ( n22531 ) ? ( n4782 ) : ( iram_180 ) ;
assign n22533 = wr_addr[7:7] ;
assign n22534 =  ( n22533 ) == ( bv_1_0_n53 )  ;
assign n22535 =  ( wr_addr ) == ( bv_8_180_n429 )  ;
assign n22536 =  ( n22534 ) & (n22535 )  ;
assign n22537 =  ( n22536 ) & (wr )  ;
assign n22538 =  ( n22537 ) ? ( n4841 ) : ( iram_180 ) ;
assign n22539 = wr_addr[7:7] ;
assign n22540 =  ( n22539 ) == ( bv_1_0_n53 )  ;
assign n22541 =  ( wr_addr ) == ( bv_8_180_n429 )  ;
assign n22542 =  ( n22540 ) & (n22541 )  ;
assign n22543 =  ( n22542 ) & (wr )  ;
assign n22544 =  ( n22543 ) ? ( n5449 ) : ( iram_180 ) ;
assign n22545 = wr_addr[7:7] ;
assign n22546 =  ( n22545 ) == ( bv_1_0_n53 )  ;
assign n22547 =  ( wr_addr ) == ( bv_8_180_n429 )  ;
assign n22548 =  ( n22546 ) & (n22547 )  ;
assign n22549 =  ( n22548 ) & (wr )  ;
assign n22550 =  ( n22549 ) ? ( n4906 ) : ( iram_180 ) ;
assign n22551 = wr_addr[7:7] ;
assign n22552 =  ( n22551 ) == ( bv_1_0_n53 )  ;
assign n22553 =  ( wr_addr ) == ( bv_8_180_n429 )  ;
assign n22554 =  ( n22552 ) & (n22553 )  ;
assign n22555 =  ( n22554 ) & (wr )  ;
assign n22556 =  ( n22555 ) ? ( n5485 ) : ( iram_180 ) ;
assign n22557 = wr_addr[7:7] ;
assign n22558 =  ( n22557 ) == ( bv_1_0_n53 )  ;
assign n22559 =  ( wr_addr ) == ( bv_8_180_n429 )  ;
assign n22560 =  ( n22558 ) & (n22559 )  ;
assign n22561 =  ( n22560 ) & (wr )  ;
assign n22562 =  ( n22561 ) ? ( n5512 ) : ( iram_180 ) ;
assign n22563 = wr_addr[7:7] ;
assign n22564 =  ( n22563 ) == ( bv_1_0_n53 )  ;
assign n22565 =  ( wr_addr ) == ( bv_8_180_n429 )  ;
assign n22566 =  ( n22564 ) & (n22565 )  ;
assign n22567 =  ( n22566 ) & (wr )  ;
assign n22568 =  ( n22567 ) ? ( bv_8_0_n69 ) : ( iram_180 ) ;
assign n22569 = wr_addr[7:7] ;
assign n22570 =  ( n22569 ) == ( bv_1_0_n53 )  ;
assign n22571 =  ( wr_addr ) == ( bv_8_180_n429 )  ;
assign n22572 =  ( n22570 ) & (n22571 )  ;
assign n22573 =  ( n22572 ) & (wr )  ;
assign n22574 =  ( n22573 ) ? ( n5071 ) : ( iram_180 ) ;
assign n22575 = wr_addr[7:7] ;
assign n22576 =  ( n22575 ) == ( bv_1_0_n53 )  ;
assign n22577 =  ( wr_addr ) == ( bv_8_180_n429 )  ;
assign n22578 =  ( n22576 ) & (n22577 )  ;
assign n22579 =  ( n22578 ) & (wr )  ;
assign n22580 =  ( n22579 ) ? ( n5096 ) : ( iram_180 ) ;
assign n22581 = wr_addr[7:7] ;
assign n22582 =  ( n22581 ) == ( bv_1_0_n53 )  ;
assign n22583 =  ( wr_addr ) == ( bv_8_180_n429 )  ;
assign n22584 =  ( n22582 ) & (n22583 )  ;
assign n22585 =  ( n22584 ) & (wr )  ;
assign n22586 =  ( n22585 ) ? ( n5123 ) : ( iram_180 ) ;
assign n22587 = wr_addr[7:7] ;
assign n22588 =  ( n22587 ) == ( bv_1_0_n53 )  ;
assign n22589 =  ( wr_addr ) == ( bv_8_180_n429 )  ;
assign n22590 =  ( n22588 ) & (n22589 )  ;
assign n22591 =  ( n22590 ) & (wr )  ;
assign n22592 =  ( n22591 ) ? ( n5165 ) : ( iram_180 ) ;
assign n22593 = wr_addr[7:7] ;
assign n22594 =  ( n22593 ) == ( bv_1_0_n53 )  ;
assign n22595 =  ( wr_addr ) == ( bv_8_180_n429 )  ;
assign n22596 =  ( n22594 ) & (n22595 )  ;
assign n22597 =  ( n22596 ) & (wr )  ;
assign n22598 =  ( n22597 ) ? ( n5204 ) : ( iram_180 ) ;
assign n22599 = wr_addr[7:7] ;
assign n22600 =  ( n22599 ) == ( bv_1_0_n53 )  ;
assign n22601 =  ( wr_addr ) == ( bv_8_180_n429 )  ;
assign n22602 =  ( n22600 ) & (n22601 )  ;
assign n22603 =  ( n22602 ) & (wr )  ;
assign n22604 =  ( n22603 ) ? ( n5262 ) : ( iram_180 ) ;
assign n22605 = wr_addr[7:7] ;
assign n22606 =  ( n22605 ) == ( bv_1_0_n53 )  ;
assign n22607 =  ( wr_addr ) == ( bv_8_180_n429 )  ;
assign n22608 =  ( n22606 ) & (n22607 )  ;
assign n22609 =  ( n22608 ) & (wr )  ;
assign n22610 =  ( n22609 ) ? ( n5298 ) : ( iram_180 ) ;
assign n22611 = wr_addr[7:7] ;
assign n22612 =  ( n22611 ) == ( bv_1_0_n53 )  ;
assign n22613 =  ( wr_addr ) == ( bv_8_180_n429 )  ;
assign n22614 =  ( n22612 ) & (n22613 )  ;
assign n22615 =  ( n22614 ) & (wr )  ;
assign n22616 =  ( n22615 ) ? ( n5325 ) : ( iram_180 ) ;
assign n22617 = wr_addr[7:7] ;
assign n22618 =  ( n22617 ) == ( bv_1_0_n53 )  ;
assign n22619 =  ( wr_addr ) == ( bv_8_181_n431 )  ;
assign n22620 =  ( n22618 ) & (n22619 )  ;
assign n22621 =  ( n22620 ) & (wr )  ;
assign n22622 =  ( n22621 ) ? ( n4782 ) : ( iram_181 ) ;
assign n22623 = wr_addr[7:7] ;
assign n22624 =  ( n22623 ) == ( bv_1_0_n53 )  ;
assign n22625 =  ( wr_addr ) == ( bv_8_181_n431 )  ;
assign n22626 =  ( n22624 ) & (n22625 )  ;
assign n22627 =  ( n22626 ) & (wr )  ;
assign n22628 =  ( n22627 ) ? ( n4841 ) : ( iram_181 ) ;
assign n22629 = wr_addr[7:7] ;
assign n22630 =  ( n22629 ) == ( bv_1_0_n53 )  ;
assign n22631 =  ( wr_addr ) == ( bv_8_181_n431 )  ;
assign n22632 =  ( n22630 ) & (n22631 )  ;
assign n22633 =  ( n22632 ) & (wr )  ;
assign n22634 =  ( n22633 ) ? ( n5449 ) : ( iram_181 ) ;
assign n22635 = wr_addr[7:7] ;
assign n22636 =  ( n22635 ) == ( bv_1_0_n53 )  ;
assign n22637 =  ( wr_addr ) == ( bv_8_181_n431 )  ;
assign n22638 =  ( n22636 ) & (n22637 )  ;
assign n22639 =  ( n22638 ) & (wr )  ;
assign n22640 =  ( n22639 ) ? ( n4906 ) : ( iram_181 ) ;
assign n22641 = wr_addr[7:7] ;
assign n22642 =  ( n22641 ) == ( bv_1_0_n53 )  ;
assign n22643 =  ( wr_addr ) == ( bv_8_181_n431 )  ;
assign n22644 =  ( n22642 ) & (n22643 )  ;
assign n22645 =  ( n22644 ) & (wr )  ;
assign n22646 =  ( n22645 ) ? ( n5485 ) : ( iram_181 ) ;
assign n22647 = wr_addr[7:7] ;
assign n22648 =  ( n22647 ) == ( bv_1_0_n53 )  ;
assign n22649 =  ( wr_addr ) == ( bv_8_181_n431 )  ;
assign n22650 =  ( n22648 ) & (n22649 )  ;
assign n22651 =  ( n22650 ) & (wr )  ;
assign n22652 =  ( n22651 ) ? ( n5512 ) : ( iram_181 ) ;
assign n22653 = wr_addr[7:7] ;
assign n22654 =  ( n22653 ) == ( bv_1_0_n53 )  ;
assign n22655 =  ( wr_addr ) == ( bv_8_181_n431 )  ;
assign n22656 =  ( n22654 ) & (n22655 )  ;
assign n22657 =  ( n22656 ) & (wr )  ;
assign n22658 =  ( n22657 ) ? ( bv_8_0_n69 ) : ( iram_181 ) ;
assign n22659 = wr_addr[7:7] ;
assign n22660 =  ( n22659 ) == ( bv_1_0_n53 )  ;
assign n22661 =  ( wr_addr ) == ( bv_8_181_n431 )  ;
assign n22662 =  ( n22660 ) & (n22661 )  ;
assign n22663 =  ( n22662 ) & (wr )  ;
assign n22664 =  ( n22663 ) ? ( n5071 ) : ( iram_181 ) ;
assign n22665 = wr_addr[7:7] ;
assign n22666 =  ( n22665 ) == ( bv_1_0_n53 )  ;
assign n22667 =  ( wr_addr ) == ( bv_8_181_n431 )  ;
assign n22668 =  ( n22666 ) & (n22667 )  ;
assign n22669 =  ( n22668 ) & (wr )  ;
assign n22670 =  ( n22669 ) ? ( n5096 ) : ( iram_181 ) ;
assign n22671 = wr_addr[7:7] ;
assign n22672 =  ( n22671 ) == ( bv_1_0_n53 )  ;
assign n22673 =  ( wr_addr ) == ( bv_8_181_n431 )  ;
assign n22674 =  ( n22672 ) & (n22673 )  ;
assign n22675 =  ( n22674 ) & (wr )  ;
assign n22676 =  ( n22675 ) ? ( n5123 ) : ( iram_181 ) ;
assign n22677 = wr_addr[7:7] ;
assign n22678 =  ( n22677 ) == ( bv_1_0_n53 )  ;
assign n22679 =  ( wr_addr ) == ( bv_8_181_n431 )  ;
assign n22680 =  ( n22678 ) & (n22679 )  ;
assign n22681 =  ( n22680 ) & (wr )  ;
assign n22682 =  ( n22681 ) ? ( n5165 ) : ( iram_181 ) ;
assign n22683 = wr_addr[7:7] ;
assign n22684 =  ( n22683 ) == ( bv_1_0_n53 )  ;
assign n22685 =  ( wr_addr ) == ( bv_8_181_n431 )  ;
assign n22686 =  ( n22684 ) & (n22685 )  ;
assign n22687 =  ( n22686 ) & (wr )  ;
assign n22688 =  ( n22687 ) ? ( n5204 ) : ( iram_181 ) ;
assign n22689 = wr_addr[7:7] ;
assign n22690 =  ( n22689 ) == ( bv_1_0_n53 )  ;
assign n22691 =  ( wr_addr ) == ( bv_8_181_n431 )  ;
assign n22692 =  ( n22690 ) & (n22691 )  ;
assign n22693 =  ( n22692 ) & (wr )  ;
assign n22694 =  ( n22693 ) ? ( n5262 ) : ( iram_181 ) ;
assign n22695 = wr_addr[7:7] ;
assign n22696 =  ( n22695 ) == ( bv_1_0_n53 )  ;
assign n22697 =  ( wr_addr ) == ( bv_8_181_n431 )  ;
assign n22698 =  ( n22696 ) & (n22697 )  ;
assign n22699 =  ( n22698 ) & (wr )  ;
assign n22700 =  ( n22699 ) ? ( n5298 ) : ( iram_181 ) ;
assign n22701 = wr_addr[7:7] ;
assign n22702 =  ( n22701 ) == ( bv_1_0_n53 )  ;
assign n22703 =  ( wr_addr ) == ( bv_8_181_n431 )  ;
assign n22704 =  ( n22702 ) & (n22703 )  ;
assign n22705 =  ( n22704 ) & (wr )  ;
assign n22706 =  ( n22705 ) ? ( n5325 ) : ( iram_181 ) ;
assign n22707 = wr_addr[7:7] ;
assign n22708 =  ( n22707 ) == ( bv_1_0_n53 )  ;
assign n22709 =  ( wr_addr ) == ( bv_8_182_n433 )  ;
assign n22710 =  ( n22708 ) & (n22709 )  ;
assign n22711 =  ( n22710 ) & (wr )  ;
assign n22712 =  ( n22711 ) ? ( n4782 ) : ( iram_182 ) ;
assign n22713 = wr_addr[7:7] ;
assign n22714 =  ( n22713 ) == ( bv_1_0_n53 )  ;
assign n22715 =  ( wr_addr ) == ( bv_8_182_n433 )  ;
assign n22716 =  ( n22714 ) & (n22715 )  ;
assign n22717 =  ( n22716 ) & (wr )  ;
assign n22718 =  ( n22717 ) ? ( n4841 ) : ( iram_182 ) ;
assign n22719 = wr_addr[7:7] ;
assign n22720 =  ( n22719 ) == ( bv_1_0_n53 )  ;
assign n22721 =  ( wr_addr ) == ( bv_8_182_n433 )  ;
assign n22722 =  ( n22720 ) & (n22721 )  ;
assign n22723 =  ( n22722 ) & (wr )  ;
assign n22724 =  ( n22723 ) ? ( n5449 ) : ( iram_182 ) ;
assign n22725 = wr_addr[7:7] ;
assign n22726 =  ( n22725 ) == ( bv_1_0_n53 )  ;
assign n22727 =  ( wr_addr ) == ( bv_8_182_n433 )  ;
assign n22728 =  ( n22726 ) & (n22727 )  ;
assign n22729 =  ( n22728 ) & (wr )  ;
assign n22730 =  ( n22729 ) ? ( n4906 ) : ( iram_182 ) ;
assign n22731 = wr_addr[7:7] ;
assign n22732 =  ( n22731 ) == ( bv_1_0_n53 )  ;
assign n22733 =  ( wr_addr ) == ( bv_8_182_n433 )  ;
assign n22734 =  ( n22732 ) & (n22733 )  ;
assign n22735 =  ( n22734 ) & (wr )  ;
assign n22736 =  ( n22735 ) ? ( n5485 ) : ( iram_182 ) ;
assign n22737 = wr_addr[7:7] ;
assign n22738 =  ( n22737 ) == ( bv_1_0_n53 )  ;
assign n22739 =  ( wr_addr ) == ( bv_8_182_n433 )  ;
assign n22740 =  ( n22738 ) & (n22739 )  ;
assign n22741 =  ( n22740 ) & (wr )  ;
assign n22742 =  ( n22741 ) ? ( n5512 ) : ( iram_182 ) ;
assign n22743 = wr_addr[7:7] ;
assign n22744 =  ( n22743 ) == ( bv_1_0_n53 )  ;
assign n22745 =  ( wr_addr ) == ( bv_8_182_n433 )  ;
assign n22746 =  ( n22744 ) & (n22745 )  ;
assign n22747 =  ( n22746 ) & (wr )  ;
assign n22748 =  ( n22747 ) ? ( bv_8_0_n69 ) : ( iram_182 ) ;
assign n22749 = wr_addr[7:7] ;
assign n22750 =  ( n22749 ) == ( bv_1_0_n53 )  ;
assign n22751 =  ( wr_addr ) == ( bv_8_182_n433 )  ;
assign n22752 =  ( n22750 ) & (n22751 )  ;
assign n22753 =  ( n22752 ) & (wr )  ;
assign n22754 =  ( n22753 ) ? ( n5071 ) : ( iram_182 ) ;
assign n22755 = wr_addr[7:7] ;
assign n22756 =  ( n22755 ) == ( bv_1_0_n53 )  ;
assign n22757 =  ( wr_addr ) == ( bv_8_182_n433 )  ;
assign n22758 =  ( n22756 ) & (n22757 )  ;
assign n22759 =  ( n22758 ) & (wr )  ;
assign n22760 =  ( n22759 ) ? ( n5096 ) : ( iram_182 ) ;
assign n22761 = wr_addr[7:7] ;
assign n22762 =  ( n22761 ) == ( bv_1_0_n53 )  ;
assign n22763 =  ( wr_addr ) == ( bv_8_182_n433 )  ;
assign n22764 =  ( n22762 ) & (n22763 )  ;
assign n22765 =  ( n22764 ) & (wr )  ;
assign n22766 =  ( n22765 ) ? ( n5123 ) : ( iram_182 ) ;
assign n22767 = wr_addr[7:7] ;
assign n22768 =  ( n22767 ) == ( bv_1_0_n53 )  ;
assign n22769 =  ( wr_addr ) == ( bv_8_182_n433 )  ;
assign n22770 =  ( n22768 ) & (n22769 )  ;
assign n22771 =  ( n22770 ) & (wr )  ;
assign n22772 =  ( n22771 ) ? ( n5165 ) : ( iram_182 ) ;
assign n22773 = wr_addr[7:7] ;
assign n22774 =  ( n22773 ) == ( bv_1_0_n53 )  ;
assign n22775 =  ( wr_addr ) == ( bv_8_182_n433 )  ;
assign n22776 =  ( n22774 ) & (n22775 )  ;
assign n22777 =  ( n22776 ) & (wr )  ;
assign n22778 =  ( n22777 ) ? ( n5204 ) : ( iram_182 ) ;
assign n22779 = wr_addr[7:7] ;
assign n22780 =  ( n22779 ) == ( bv_1_0_n53 )  ;
assign n22781 =  ( wr_addr ) == ( bv_8_182_n433 )  ;
assign n22782 =  ( n22780 ) & (n22781 )  ;
assign n22783 =  ( n22782 ) & (wr )  ;
assign n22784 =  ( n22783 ) ? ( n5262 ) : ( iram_182 ) ;
assign n22785 = wr_addr[7:7] ;
assign n22786 =  ( n22785 ) == ( bv_1_0_n53 )  ;
assign n22787 =  ( wr_addr ) == ( bv_8_182_n433 )  ;
assign n22788 =  ( n22786 ) & (n22787 )  ;
assign n22789 =  ( n22788 ) & (wr )  ;
assign n22790 =  ( n22789 ) ? ( n5298 ) : ( iram_182 ) ;
assign n22791 = wr_addr[7:7] ;
assign n22792 =  ( n22791 ) == ( bv_1_0_n53 )  ;
assign n22793 =  ( wr_addr ) == ( bv_8_182_n433 )  ;
assign n22794 =  ( n22792 ) & (n22793 )  ;
assign n22795 =  ( n22794 ) & (wr )  ;
assign n22796 =  ( n22795 ) ? ( n5325 ) : ( iram_182 ) ;
assign n22797 = wr_addr[7:7] ;
assign n22798 =  ( n22797 ) == ( bv_1_0_n53 )  ;
assign n22799 =  ( wr_addr ) == ( bv_8_183_n435 )  ;
assign n22800 =  ( n22798 ) & (n22799 )  ;
assign n22801 =  ( n22800 ) & (wr )  ;
assign n22802 =  ( n22801 ) ? ( n4782 ) : ( iram_183 ) ;
assign n22803 = wr_addr[7:7] ;
assign n22804 =  ( n22803 ) == ( bv_1_0_n53 )  ;
assign n22805 =  ( wr_addr ) == ( bv_8_183_n435 )  ;
assign n22806 =  ( n22804 ) & (n22805 )  ;
assign n22807 =  ( n22806 ) & (wr )  ;
assign n22808 =  ( n22807 ) ? ( n4841 ) : ( iram_183 ) ;
assign n22809 = wr_addr[7:7] ;
assign n22810 =  ( n22809 ) == ( bv_1_0_n53 )  ;
assign n22811 =  ( wr_addr ) == ( bv_8_183_n435 )  ;
assign n22812 =  ( n22810 ) & (n22811 )  ;
assign n22813 =  ( n22812 ) & (wr )  ;
assign n22814 =  ( n22813 ) ? ( n5449 ) : ( iram_183 ) ;
assign n22815 = wr_addr[7:7] ;
assign n22816 =  ( n22815 ) == ( bv_1_0_n53 )  ;
assign n22817 =  ( wr_addr ) == ( bv_8_183_n435 )  ;
assign n22818 =  ( n22816 ) & (n22817 )  ;
assign n22819 =  ( n22818 ) & (wr )  ;
assign n22820 =  ( n22819 ) ? ( n4906 ) : ( iram_183 ) ;
assign n22821 = wr_addr[7:7] ;
assign n22822 =  ( n22821 ) == ( bv_1_0_n53 )  ;
assign n22823 =  ( wr_addr ) == ( bv_8_183_n435 )  ;
assign n22824 =  ( n22822 ) & (n22823 )  ;
assign n22825 =  ( n22824 ) & (wr )  ;
assign n22826 =  ( n22825 ) ? ( n5485 ) : ( iram_183 ) ;
assign n22827 = wr_addr[7:7] ;
assign n22828 =  ( n22827 ) == ( bv_1_0_n53 )  ;
assign n22829 =  ( wr_addr ) == ( bv_8_183_n435 )  ;
assign n22830 =  ( n22828 ) & (n22829 )  ;
assign n22831 =  ( n22830 ) & (wr )  ;
assign n22832 =  ( n22831 ) ? ( n5512 ) : ( iram_183 ) ;
assign n22833 = wr_addr[7:7] ;
assign n22834 =  ( n22833 ) == ( bv_1_0_n53 )  ;
assign n22835 =  ( wr_addr ) == ( bv_8_183_n435 )  ;
assign n22836 =  ( n22834 ) & (n22835 )  ;
assign n22837 =  ( n22836 ) & (wr )  ;
assign n22838 =  ( n22837 ) ? ( bv_8_0_n69 ) : ( iram_183 ) ;
assign n22839 = wr_addr[7:7] ;
assign n22840 =  ( n22839 ) == ( bv_1_0_n53 )  ;
assign n22841 =  ( wr_addr ) == ( bv_8_183_n435 )  ;
assign n22842 =  ( n22840 ) & (n22841 )  ;
assign n22843 =  ( n22842 ) & (wr )  ;
assign n22844 =  ( n22843 ) ? ( n5071 ) : ( iram_183 ) ;
assign n22845 = wr_addr[7:7] ;
assign n22846 =  ( n22845 ) == ( bv_1_0_n53 )  ;
assign n22847 =  ( wr_addr ) == ( bv_8_183_n435 )  ;
assign n22848 =  ( n22846 ) & (n22847 )  ;
assign n22849 =  ( n22848 ) & (wr )  ;
assign n22850 =  ( n22849 ) ? ( n5096 ) : ( iram_183 ) ;
assign n22851 = wr_addr[7:7] ;
assign n22852 =  ( n22851 ) == ( bv_1_0_n53 )  ;
assign n22853 =  ( wr_addr ) == ( bv_8_183_n435 )  ;
assign n22854 =  ( n22852 ) & (n22853 )  ;
assign n22855 =  ( n22854 ) & (wr )  ;
assign n22856 =  ( n22855 ) ? ( n5123 ) : ( iram_183 ) ;
assign n22857 = wr_addr[7:7] ;
assign n22858 =  ( n22857 ) == ( bv_1_0_n53 )  ;
assign n22859 =  ( wr_addr ) == ( bv_8_183_n435 )  ;
assign n22860 =  ( n22858 ) & (n22859 )  ;
assign n22861 =  ( n22860 ) & (wr )  ;
assign n22862 =  ( n22861 ) ? ( n5165 ) : ( iram_183 ) ;
assign n22863 = wr_addr[7:7] ;
assign n22864 =  ( n22863 ) == ( bv_1_0_n53 )  ;
assign n22865 =  ( wr_addr ) == ( bv_8_183_n435 )  ;
assign n22866 =  ( n22864 ) & (n22865 )  ;
assign n22867 =  ( n22866 ) & (wr )  ;
assign n22868 =  ( n22867 ) ? ( n5204 ) : ( iram_183 ) ;
assign n22869 = wr_addr[7:7] ;
assign n22870 =  ( n22869 ) == ( bv_1_0_n53 )  ;
assign n22871 =  ( wr_addr ) == ( bv_8_183_n435 )  ;
assign n22872 =  ( n22870 ) & (n22871 )  ;
assign n22873 =  ( n22872 ) & (wr )  ;
assign n22874 =  ( n22873 ) ? ( n5262 ) : ( iram_183 ) ;
assign n22875 = wr_addr[7:7] ;
assign n22876 =  ( n22875 ) == ( bv_1_0_n53 )  ;
assign n22877 =  ( wr_addr ) == ( bv_8_183_n435 )  ;
assign n22878 =  ( n22876 ) & (n22877 )  ;
assign n22879 =  ( n22878 ) & (wr )  ;
assign n22880 =  ( n22879 ) ? ( n5298 ) : ( iram_183 ) ;
assign n22881 = wr_addr[7:7] ;
assign n22882 =  ( n22881 ) == ( bv_1_0_n53 )  ;
assign n22883 =  ( wr_addr ) == ( bv_8_183_n435 )  ;
assign n22884 =  ( n22882 ) & (n22883 )  ;
assign n22885 =  ( n22884 ) & (wr )  ;
assign n22886 =  ( n22885 ) ? ( n5325 ) : ( iram_183 ) ;
assign n22887 = wr_addr[7:7] ;
assign n22888 =  ( n22887 ) == ( bv_1_0_n53 )  ;
assign n22889 =  ( wr_addr ) == ( bv_8_184_n437 )  ;
assign n22890 =  ( n22888 ) & (n22889 )  ;
assign n22891 =  ( n22890 ) & (wr )  ;
assign n22892 =  ( n22891 ) ? ( n4782 ) : ( iram_184 ) ;
assign n22893 = wr_addr[7:7] ;
assign n22894 =  ( n22893 ) == ( bv_1_0_n53 )  ;
assign n22895 =  ( wr_addr ) == ( bv_8_184_n437 )  ;
assign n22896 =  ( n22894 ) & (n22895 )  ;
assign n22897 =  ( n22896 ) & (wr )  ;
assign n22898 =  ( n22897 ) ? ( n4841 ) : ( iram_184 ) ;
assign n22899 = wr_addr[7:7] ;
assign n22900 =  ( n22899 ) == ( bv_1_0_n53 )  ;
assign n22901 =  ( wr_addr ) == ( bv_8_184_n437 )  ;
assign n22902 =  ( n22900 ) & (n22901 )  ;
assign n22903 =  ( n22902 ) & (wr )  ;
assign n22904 =  ( n22903 ) ? ( n5449 ) : ( iram_184 ) ;
assign n22905 = wr_addr[7:7] ;
assign n22906 =  ( n22905 ) == ( bv_1_0_n53 )  ;
assign n22907 =  ( wr_addr ) == ( bv_8_184_n437 )  ;
assign n22908 =  ( n22906 ) & (n22907 )  ;
assign n22909 =  ( n22908 ) & (wr )  ;
assign n22910 =  ( n22909 ) ? ( n4906 ) : ( iram_184 ) ;
assign n22911 = wr_addr[7:7] ;
assign n22912 =  ( n22911 ) == ( bv_1_0_n53 )  ;
assign n22913 =  ( wr_addr ) == ( bv_8_184_n437 )  ;
assign n22914 =  ( n22912 ) & (n22913 )  ;
assign n22915 =  ( n22914 ) & (wr )  ;
assign n22916 =  ( n22915 ) ? ( n5485 ) : ( iram_184 ) ;
assign n22917 = wr_addr[7:7] ;
assign n22918 =  ( n22917 ) == ( bv_1_0_n53 )  ;
assign n22919 =  ( wr_addr ) == ( bv_8_184_n437 )  ;
assign n22920 =  ( n22918 ) & (n22919 )  ;
assign n22921 =  ( n22920 ) & (wr )  ;
assign n22922 =  ( n22921 ) ? ( n5512 ) : ( iram_184 ) ;
assign n22923 = wr_addr[7:7] ;
assign n22924 =  ( n22923 ) == ( bv_1_0_n53 )  ;
assign n22925 =  ( wr_addr ) == ( bv_8_184_n437 )  ;
assign n22926 =  ( n22924 ) & (n22925 )  ;
assign n22927 =  ( n22926 ) & (wr )  ;
assign n22928 =  ( n22927 ) ? ( bv_8_0_n69 ) : ( iram_184 ) ;
assign n22929 = wr_addr[7:7] ;
assign n22930 =  ( n22929 ) == ( bv_1_0_n53 )  ;
assign n22931 =  ( wr_addr ) == ( bv_8_184_n437 )  ;
assign n22932 =  ( n22930 ) & (n22931 )  ;
assign n22933 =  ( n22932 ) & (wr )  ;
assign n22934 =  ( n22933 ) ? ( n5071 ) : ( iram_184 ) ;
assign n22935 = wr_addr[7:7] ;
assign n22936 =  ( n22935 ) == ( bv_1_0_n53 )  ;
assign n22937 =  ( wr_addr ) == ( bv_8_184_n437 )  ;
assign n22938 =  ( n22936 ) & (n22937 )  ;
assign n22939 =  ( n22938 ) & (wr )  ;
assign n22940 =  ( n22939 ) ? ( n5096 ) : ( iram_184 ) ;
assign n22941 = wr_addr[7:7] ;
assign n22942 =  ( n22941 ) == ( bv_1_0_n53 )  ;
assign n22943 =  ( wr_addr ) == ( bv_8_184_n437 )  ;
assign n22944 =  ( n22942 ) & (n22943 )  ;
assign n22945 =  ( n22944 ) & (wr )  ;
assign n22946 =  ( n22945 ) ? ( n5123 ) : ( iram_184 ) ;
assign n22947 = wr_addr[7:7] ;
assign n22948 =  ( n22947 ) == ( bv_1_0_n53 )  ;
assign n22949 =  ( wr_addr ) == ( bv_8_184_n437 )  ;
assign n22950 =  ( n22948 ) & (n22949 )  ;
assign n22951 =  ( n22950 ) & (wr )  ;
assign n22952 =  ( n22951 ) ? ( n5165 ) : ( iram_184 ) ;
assign n22953 = wr_addr[7:7] ;
assign n22954 =  ( n22953 ) == ( bv_1_0_n53 )  ;
assign n22955 =  ( wr_addr ) == ( bv_8_184_n437 )  ;
assign n22956 =  ( n22954 ) & (n22955 )  ;
assign n22957 =  ( n22956 ) & (wr )  ;
assign n22958 =  ( n22957 ) ? ( n5204 ) : ( iram_184 ) ;
assign n22959 = wr_addr[7:7] ;
assign n22960 =  ( n22959 ) == ( bv_1_0_n53 )  ;
assign n22961 =  ( wr_addr ) == ( bv_8_184_n437 )  ;
assign n22962 =  ( n22960 ) & (n22961 )  ;
assign n22963 =  ( n22962 ) & (wr )  ;
assign n22964 =  ( n22963 ) ? ( n5262 ) : ( iram_184 ) ;
assign n22965 = wr_addr[7:7] ;
assign n22966 =  ( n22965 ) == ( bv_1_0_n53 )  ;
assign n22967 =  ( wr_addr ) == ( bv_8_184_n437 )  ;
assign n22968 =  ( n22966 ) & (n22967 )  ;
assign n22969 =  ( n22968 ) & (wr )  ;
assign n22970 =  ( n22969 ) ? ( n5298 ) : ( iram_184 ) ;
assign n22971 = wr_addr[7:7] ;
assign n22972 =  ( n22971 ) == ( bv_1_0_n53 )  ;
assign n22973 =  ( wr_addr ) == ( bv_8_184_n437 )  ;
assign n22974 =  ( n22972 ) & (n22973 )  ;
assign n22975 =  ( n22974 ) & (wr )  ;
assign n22976 =  ( n22975 ) ? ( n5325 ) : ( iram_184 ) ;
assign n22977 = wr_addr[7:7] ;
assign n22978 =  ( n22977 ) == ( bv_1_0_n53 )  ;
assign n22979 =  ( wr_addr ) == ( bv_8_185_n439 )  ;
assign n22980 =  ( n22978 ) & (n22979 )  ;
assign n22981 =  ( n22980 ) & (wr )  ;
assign n22982 =  ( n22981 ) ? ( n4782 ) : ( iram_185 ) ;
assign n22983 = wr_addr[7:7] ;
assign n22984 =  ( n22983 ) == ( bv_1_0_n53 )  ;
assign n22985 =  ( wr_addr ) == ( bv_8_185_n439 )  ;
assign n22986 =  ( n22984 ) & (n22985 )  ;
assign n22987 =  ( n22986 ) & (wr )  ;
assign n22988 =  ( n22987 ) ? ( n4841 ) : ( iram_185 ) ;
assign n22989 = wr_addr[7:7] ;
assign n22990 =  ( n22989 ) == ( bv_1_0_n53 )  ;
assign n22991 =  ( wr_addr ) == ( bv_8_185_n439 )  ;
assign n22992 =  ( n22990 ) & (n22991 )  ;
assign n22993 =  ( n22992 ) & (wr )  ;
assign n22994 =  ( n22993 ) ? ( n5449 ) : ( iram_185 ) ;
assign n22995 = wr_addr[7:7] ;
assign n22996 =  ( n22995 ) == ( bv_1_0_n53 )  ;
assign n22997 =  ( wr_addr ) == ( bv_8_185_n439 )  ;
assign n22998 =  ( n22996 ) & (n22997 )  ;
assign n22999 =  ( n22998 ) & (wr )  ;
assign n23000 =  ( n22999 ) ? ( n4906 ) : ( iram_185 ) ;
assign n23001 = wr_addr[7:7] ;
assign n23002 =  ( n23001 ) == ( bv_1_0_n53 )  ;
assign n23003 =  ( wr_addr ) == ( bv_8_185_n439 )  ;
assign n23004 =  ( n23002 ) & (n23003 )  ;
assign n23005 =  ( n23004 ) & (wr )  ;
assign n23006 =  ( n23005 ) ? ( n5485 ) : ( iram_185 ) ;
assign n23007 = wr_addr[7:7] ;
assign n23008 =  ( n23007 ) == ( bv_1_0_n53 )  ;
assign n23009 =  ( wr_addr ) == ( bv_8_185_n439 )  ;
assign n23010 =  ( n23008 ) & (n23009 )  ;
assign n23011 =  ( n23010 ) & (wr )  ;
assign n23012 =  ( n23011 ) ? ( n5512 ) : ( iram_185 ) ;
assign n23013 = wr_addr[7:7] ;
assign n23014 =  ( n23013 ) == ( bv_1_0_n53 )  ;
assign n23015 =  ( wr_addr ) == ( bv_8_185_n439 )  ;
assign n23016 =  ( n23014 ) & (n23015 )  ;
assign n23017 =  ( n23016 ) & (wr )  ;
assign n23018 =  ( n23017 ) ? ( bv_8_0_n69 ) : ( iram_185 ) ;
assign n23019 = wr_addr[7:7] ;
assign n23020 =  ( n23019 ) == ( bv_1_0_n53 )  ;
assign n23021 =  ( wr_addr ) == ( bv_8_185_n439 )  ;
assign n23022 =  ( n23020 ) & (n23021 )  ;
assign n23023 =  ( n23022 ) & (wr )  ;
assign n23024 =  ( n23023 ) ? ( n5071 ) : ( iram_185 ) ;
assign n23025 = wr_addr[7:7] ;
assign n23026 =  ( n23025 ) == ( bv_1_0_n53 )  ;
assign n23027 =  ( wr_addr ) == ( bv_8_185_n439 )  ;
assign n23028 =  ( n23026 ) & (n23027 )  ;
assign n23029 =  ( n23028 ) & (wr )  ;
assign n23030 =  ( n23029 ) ? ( n5096 ) : ( iram_185 ) ;
assign n23031 = wr_addr[7:7] ;
assign n23032 =  ( n23031 ) == ( bv_1_0_n53 )  ;
assign n23033 =  ( wr_addr ) == ( bv_8_185_n439 )  ;
assign n23034 =  ( n23032 ) & (n23033 )  ;
assign n23035 =  ( n23034 ) & (wr )  ;
assign n23036 =  ( n23035 ) ? ( n5123 ) : ( iram_185 ) ;
assign n23037 = wr_addr[7:7] ;
assign n23038 =  ( n23037 ) == ( bv_1_0_n53 )  ;
assign n23039 =  ( wr_addr ) == ( bv_8_185_n439 )  ;
assign n23040 =  ( n23038 ) & (n23039 )  ;
assign n23041 =  ( n23040 ) & (wr )  ;
assign n23042 =  ( n23041 ) ? ( n5165 ) : ( iram_185 ) ;
assign n23043 = wr_addr[7:7] ;
assign n23044 =  ( n23043 ) == ( bv_1_0_n53 )  ;
assign n23045 =  ( wr_addr ) == ( bv_8_185_n439 )  ;
assign n23046 =  ( n23044 ) & (n23045 )  ;
assign n23047 =  ( n23046 ) & (wr )  ;
assign n23048 =  ( n23047 ) ? ( n5204 ) : ( iram_185 ) ;
assign n23049 = wr_addr[7:7] ;
assign n23050 =  ( n23049 ) == ( bv_1_0_n53 )  ;
assign n23051 =  ( wr_addr ) == ( bv_8_185_n439 )  ;
assign n23052 =  ( n23050 ) & (n23051 )  ;
assign n23053 =  ( n23052 ) & (wr )  ;
assign n23054 =  ( n23053 ) ? ( n5262 ) : ( iram_185 ) ;
assign n23055 = wr_addr[7:7] ;
assign n23056 =  ( n23055 ) == ( bv_1_0_n53 )  ;
assign n23057 =  ( wr_addr ) == ( bv_8_185_n439 )  ;
assign n23058 =  ( n23056 ) & (n23057 )  ;
assign n23059 =  ( n23058 ) & (wr )  ;
assign n23060 =  ( n23059 ) ? ( n5298 ) : ( iram_185 ) ;
assign n23061 = wr_addr[7:7] ;
assign n23062 =  ( n23061 ) == ( bv_1_0_n53 )  ;
assign n23063 =  ( wr_addr ) == ( bv_8_185_n439 )  ;
assign n23064 =  ( n23062 ) & (n23063 )  ;
assign n23065 =  ( n23064 ) & (wr )  ;
assign n23066 =  ( n23065 ) ? ( n5325 ) : ( iram_185 ) ;
assign n23067 = wr_addr[7:7] ;
assign n23068 =  ( n23067 ) == ( bv_1_0_n53 )  ;
assign n23069 =  ( wr_addr ) == ( bv_8_186_n441 )  ;
assign n23070 =  ( n23068 ) & (n23069 )  ;
assign n23071 =  ( n23070 ) & (wr )  ;
assign n23072 =  ( n23071 ) ? ( n4782 ) : ( iram_186 ) ;
assign n23073 = wr_addr[7:7] ;
assign n23074 =  ( n23073 ) == ( bv_1_0_n53 )  ;
assign n23075 =  ( wr_addr ) == ( bv_8_186_n441 )  ;
assign n23076 =  ( n23074 ) & (n23075 )  ;
assign n23077 =  ( n23076 ) & (wr )  ;
assign n23078 =  ( n23077 ) ? ( n4841 ) : ( iram_186 ) ;
assign n23079 = wr_addr[7:7] ;
assign n23080 =  ( n23079 ) == ( bv_1_0_n53 )  ;
assign n23081 =  ( wr_addr ) == ( bv_8_186_n441 )  ;
assign n23082 =  ( n23080 ) & (n23081 )  ;
assign n23083 =  ( n23082 ) & (wr )  ;
assign n23084 =  ( n23083 ) ? ( n5449 ) : ( iram_186 ) ;
assign n23085 = wr_addr[7:7] ;
assign n23086 =  ( n23085 ) == ( bv_1_0_n53 )  ;
assign n23087 =  ( wr_addr ) == ( bv_8_186_n441 )  ;
assign n23088 =  ( n23086 ) & (n23087 )  ;
assign n23089 =  ( n23088 ) & (wr )  ;
assign n23090 =  ( n23089 ) ? ( n4906 ) : ( iram_186 ) ;
assign n23091 = wr_addr[7:7] ;
assign n23092 =  ( n23091 ) == ( bv_1_0_n53 )  ;
assign n23093 =  ( wr_addr ) == ( bv_8_186_n441 )  ;
assign n23094 =  ( n23092 ) & (n23093 )  ;
assign n23095 =  ( n23094 ) & (wr )  ;
assign n23096 =  ( n23095 ) ? ( n5485 ) : ( iram_186 ) ;
assign n23097 = wr_addr[7:7] ;
assign n23098 =  ( n23097 ) == ( bv_1_0_n53 )  ;
assign n23099 =  ( wr_addr ) == ( bv_8_186_n441 )  ;
assign n23100 =  ( n23098 ) & (n23099 )  ;
assign n23101 =  ( n23100 ) & (wr )  ;
assign n23102 =  ( n23101 ) ? ( n5512 ) : ( iram_186 ) ;
assign n23103 = wr_addr[7:7] ;
assign n23104 =  ( n23103 ) == ( bv_1_0_n53 )  ;
assign n23105 =  ( wr_addr ) == ( bv_8_186_n441 )  ;
assign n23106 =  ( n23104 ) & (n23105 )  ;
assign n23107 =  ( n23106 ) & (wr )  ;
assign n23108 =  ( n23107 ) ? ( bv_8_0_n69 ) : ( iram_186 ) ;
assign n23109 = wr_addr[7:7] ;
assign n23110 =  ( n23109 ) == ( bv_1_0_n53 )  ;
assign n23111 =  ( wr_addr ) == ( bv_8_186_n441 )  ;
assign n23112 =  ( n23110 ) & (n23111 )  ;
assign n23113 =  ( n23112 ) & (wr )  ;
assign n23114 =  ( n23113 ) ? ( n5071 ) : ( iram_186 ) ;
assign n23115 = wr_addr[7:7] ;
assign n23116 =  ( n23115 ) == ( bv_1_0_n53 )  ;
assign n23117 =  ( wr_addr ) == ( bv_8_186_n441 )  ;
assign n23118 =  ( n23116 ) & (n23117 )  ;
assign n23119 =  ( n23118 ) & (wr )  ;
assign n23120 =  ( n23119 ) ? ( n5096 ) : ( iram_186 ) ;
assign n23121 = wr_addr[7:7] ;
assign n23122 =  ( n23121 ) == ( bv_1_0_n53 )  ;
assign n23123 =  ( wr_addr ) == ( bv_8_186_n441 )  ;
assign n23124 =  ( n23122 ) & (n23123 )  ;
assign n23125 =  ( n23124 ) & (wr )  ;
assign n23126 =  ( n23125 ) ? ( n5123 ) : ( iram_186 ) ;
assign n23127 = wr_addr[7:7] ;
assign n23128 =  ( n23127 ) == ( bv_1_0_n53 )  ;
assign n23129 =  ( wr_addr ) == ( bv_8_186_n441 )  ;
assign n23130 =  ( n23128 ) & (n23129 )  ;
assign n23131 =  ( n23130 ) & (wr )  ;
assign n23132 =  ( n23131 ) ? ( n5165 ) : ( iram_186 ) ;
assign n23133 = wr_addr[7:7] ;
assign n23134 =  ( n23133 ) == ( bv_1_0_n53 )  ;
assign n23135 =  ( wr_addr ) == ( bv_8_186_n441 )  ;
assign n23136 =  ( n23134 ) & (n23135 )  ;
assign n23137 =  ( n23136 ) & (wr )  ;
assign n23138 =  ( n23137 ) ? ( n5204 ) : ( iram_186 ) ;
assign n23139 = wr_addr[7:7] ;
assign n23140 =  ( n23139 ) == ( bv_1_0_n53 )  ;
assign n23141 =  ( wr_addr ) == ( bv_8_186_n441 )  ;
assign n23142 =  ( n23140 ) & (n23141 )  ;
assign n23143 =  ( n23142 ) & (wr )  ;
assign n23144 =  ( n23143 ) ? ( n5262 ) : ( iram_186 ) ;
assign n23145 = wr_addr[7:7] ;
assign n23146 =  ( n23145 ) == ( bv_1_0_n53 )  ;
assign n23147 =  ( wr_addr ) == ( bv_8_186_n441 )  ;
assign n23148 =  ( n23146 ) & (n23147 )  ;
assign n23149 =  ( n23148 ) & (wr )  ;
assign n23150 =  ( n23149 ) ? ( n5298 ) : ( iram_186 ) ;
assign n23151 = wr_addr[7:7] ;
assign n23152 =  ( n23151 ) == ( bv_1_0_n53 )  ;
assign n23153 =  ( wr_addr ) == ( bv_8_186_n441 )  ;
assign n23154 =  ( n23152 ) & (n23153 )  ;
assign n23155 =  ( n23154 ) & (wr )  ;
assign n23156 =  ( n23155 ) ? ( n5325 ) : ( iram_186 ) ;
assign n23157 = wr_addr[7:7] ;
assign n23158 =  ( n23157 ) == ( bv_1_0_n53 )  ;
assign n23159 =  ( wr_addr ) == ( bv_8_187_n443 )  ;
assign n23160 =  ( n23158 ) & (n23159 )  ;
assign n23161 =  ( n23160 ) & (wr )  ;
assign n23162 =  ( n23161 ) ? ( n4782 ) : ( iram_187 ) ;
assign n23163 = wr_addr[7:7] ;
assign n23164 =  ( n23163 ) == ( bv_1_0_n53 )  ;
assign n23165 =  ( wr_addr ) == ( bv_8_187_n443 )  ;
assign n23166 =  ( n23164 ) & (n23165 )  ;
assign n23167 =  ( n23166 ) & (wr )  ;
assign n23168 =  ( n23167 ) ? ( n4841 ) : ( iram_187 ) ;
assign n23169 = wr_addr[7:7] ;
assign n23170 =  ( n23169 ) == ( bv_1_0_n53 )  ;
assign n23171 =  ( wr_addr ) == ( bv_8_187_n443 )  ;
assign n23172 =  ( n23170 ) & (n23171 )  ;
assign n23173 =  ( n23172 ) & (wr )  ;
assign n23174 =  ( n23173 ) ? ( n5449 ) : ( iram_187 ) ;
assign n23175 = wr_addr[7:7] ;
assign n23176 =  ( n23175 ) == ( bv_1_0_n53 )  ;
assign n23177 =  ( wr_addr ) == ( bv_8_187_n443 )  ;
assign n23178 =  ( n23176 ) & (n23177 )  ;
assign n23179 =  ( n23178 ) & (wr )  ;
assign n23180 =  ( n23179 ) ? ( n4906 ) : ( iram_187 ) ;
assign n23181 = wr_addr[7:7] ;
assign n23182 =  ( n23181 ) == ( bv_1_0_n53 )  ;
assign n23183 =  ( wr_addr ) == ( bv_8_187_n443 )  ;
assign n23184 =  ( n23182 ) & (n23183 )  ;
assign n23185 =  ( n23184 ) & (wr )  ;
assign n23186 =  ( n23185 ) ? ( n5485 ) : ( iram_187 ) ;
assign n23187 = wr_addr[7:7] ;
assign n23188 =  ( n23187 ) == ( bv_1_0_n53 )  ;
assign n23189 =  ( wr_addr ) == ( bv_8_187_n443 )  ;
assign n23190 =  ( n23188 ) & (n23189 )  ;
assign n23191 =  ( n23190 ) & (wr )  ;
assign n23192 =  ( n23191 ) ? ( n5512 ) : ( iram_187 ) ;
assign n23193 = wr_addr[7:7] ;
assign n23194 =  ( n23193 ) == ( bv_1_0_n53 )  ;
assign n23195 =  ( wr_addr ) == ( bv_8_187_n443 )  ;
assign n23196 =  ( n23194 ) & (n23195 )  ;
assign n23197 =  ( n23196 ) & (wr )  ;
assign n23198 =  ( n23197 ) ? ( bv_8_0_n69 ) : ( iram_187 ) ;
assign n23199 = wr_addr[7:7] ;
assign n23200 =  ( n23199 ) == ( bv_1_0_n53 )  ;
assign n23201 =  ( wr_addr ) == ( bv_8_187_n443 )  ;
assign n23202 =  ( n23200 ) & (n23201 )  ;
assign n23203 =  ( n23202 ) & (wr )  ;
assign n23204 =  ( n23203 ) ? ( n5071 ) : ( iram_187 ) ;
assign n23205 = wr_addr[7:7] ;
assign n23206 =  ( n23205 ) == ( bv_1_0_n53 )  ;
assign n23207 =  ( wr_addr ) == ( bv_8_187_n443 )  ;
assign n23208 =  ( n23206 ) & (n23207 )  ;
assign n23209 =  ( n23208 ) & (wr )  ;
assign n23210 =  ( n23209 ) ? ( n5096 ) : ( iram_187 ) ;
assign n23211 = wr_addr[7:7] ;
assign n23212 =  ( n23211 ) == ( bv_1_0_n53 )  ;
assign n23213 =  ( wr_addr ) == ( bv_8_187_n443 )  ;
assign n23214 =  ( n23212 ) & (n23213 )  ;
assign n23215 =  ( n23214 ) & (wr )  ;
assign n23216 =  ( n23215 ) ? ( n5123 ) : ( iram_187 ) ;
assign n23217 = wr_addr[7:7] ;
assign n23218 =  ( n23217 ) == ( bv_1_0_n53 )  ;
assign n23219 =  ( wr_addr ) == ( bv_8_187_n443 )  ;
assign n23220 =  ( n23218 ) & (n23219 )  ;
assign n23221 =  ( n23220 ) & (wr )  ;
assign n23222 =  ( n23221 ) ? ( n5165 ) : ( iram_187 ) ;
assign n23223 = wr_addr[7:7] ;
assign n23224 =  ( n23223 ) == ( bv_1_0_n53 )  ;
assign n23225 =  ( wr_addr ) == ( bv_8_187_n443 )  ;
assign n23226 =  ( n23224 ) & (n23225 )  ;
assign n23227 =  ( n23226 ) & (wr )  ;
assign n23228 =  ( n23227 ) ? ( n5204 ) : ( iram_187 ) ;
assign n23229 = wr_addr[7:7] ;
assign n23230 =  ( n23229 ) == ( bv_1_0_n53 )  ;
assign n23231 =  ( wr_addr ) == ( bv_8_187_n443 )  ;
assign n23232 =  ( n23230 ) & (n23231 )  ;
assign n23233 =  ( n23232 ) & (wr )  ;
assign n23234 =  ( n23233 ) ? ( n5262 ) : ( iram_187 ) ;
assign n23235 = wr_addr[7:7] ;
assign n23236 =  ( n23235 ) == ( bv_1_0_n53 )  ;
assign n23237 =  ( wr_addr ) == ( bv_8_187_n443 )  ;
assign n23238 =  ( n23236 ) & (n23237 )  ;
assign n23239 =  ( n23238 ) & (wr )  ;
assign n23240 =  ( n23239 ) ? ( n5298 ) : ( iram_187 ) ;
assign n23241 = wr_addr[7:7] ;
assign n23242 =  ( n23241 ) == ( bv_1_0_n53 )  ;
assign n23243 =  ( wr_addr ) == ( bv_8_187_n443 )  ;
assign n23244 =  ( n23242 ) & (n23243 )  ;
assign n23245 =  ( n23244 ) & (wr )  ;
assign n23246 =  ( n23245 ) ? ( n5325 ) : ( iram_187 ) ;
assign n23247 = wr_addr[7:7] ;
assign n23248 =  ( n23247 ) == ( bv_1_0_n53 )  ;
assign n23249 =  ( wr_addr ) == ( bv_8_188_n445 )  ;
assign n23250 =  ( n23248 ) & (n23249 )  ;
assign n23251 =  ( n23250 ) & (wr )  ;
assign n23252 =  ( n23251 ) ? ( n4782 ) : ( iram_188 ) ;
assign n23253 = wr_addr[7:7] ;
assign n23254 =  ( n23253 ) == ( bv_1_0_n53 )  ;
assign n23255 =  ( wr_addr ) == ( bv_8_188_n445 )  ;
assign n23256 =  ( n23254 ) & (n23255 )  ;
assign n23257 =  ( n23256 ) & (wr )  ;
assign n23258 =  ( n23257 ) ? ( n4841 ) : ( iram_188 ) ;
assign n23259 = wr_addr[7:7] ;
assign n23260 =  ( n23259 ) == ( bv_1_0_n53 )  ;
assign n23261 =  ( wr_addr ) == ( bv_8_188_n445 )  ;
assign n23262 =  ( n23260 ) & (n23261 )  ;
assign n23263 =  ( n23262 ) & (wr )  ;
assign n23264 =  ( n23263 ) ? ( n5449 ) : ( iram_188 ) ;
assign n23265 = wr_addr[7:7] ;
assign n23266 =  ( n23265 ) == ( bv_1_0_n53 )  ;
assign n23267 =  ( wr_addr ) == ( bv_8_188_n445 )  ;
assign n23268 =  ( n23266 ) & (n23267 )  ;
assign n23269 =  ( n23268 ) & (wr )  ;
assign n23270 =  ( n23269 ) ? ( n4906 ) : ( iram_188 ) ;
assign n23271 = wr_addr[7:7] ;
assign n23272 =  ( n23271 ) == ( bv_1_0_n53 )  ;
assign n23273 =  ( wr_addr ) == ( bv_8_188_n445 )  ;
assign n23274 =  ( n23272 ) & (n23273 )  ;
assign n23275 =  ( n23274 ) & (wr )  ;
assign n23276 =  ( n23275 ) ? ( n5485 ) : ( iram_188 ) ;
assign n23277 = wr_addr[7:7] ;
assign n23278 =  ( n23277 ) == ( bv_1_0_n53 )  ;
assign n23279 =  ( wr_addr ) == ( bv_8_188_n445 )  ;
assign n23280 =  ( n23278 ) & (n23279 )  ;
assign n23281 =  ( n23280 ) & (wr )  ;
assign n23282 =  ( n23281 ) ? ( n5512 ) : ( iram_188 ) ;
assign n23283 = wr_addr[7:7] ;
assign n23284 =  ( n23283 ) == ( bv_1_0_n53 )  ;
assign n23285 =  ( wr_addr ) == ( bv_8_188_n445 )  ;
assign n23286 =  ( n23284 ) & (n23285 )  ;
assign n23287 =  ( n23286 ) & (wr )  ;
assign n23288 =  ( n23287 ) ? ( bv_8_0_n69 ) : ( iram_188 ) ;
assign n23289 = wr_addr[7:7] ;
assign n23290 =  ( n23289 ) == ( bv_1_0_n53 )  ;
assign n23291 =  ( wr_addr ) == ( bv_8_188_n445 )  ;
assign n23292 =  ( n23290 ) & (n23291 )  ;
assign n23293 =  ( n23292 ) & (wr )  ;
assign n23294 =  ( n23293 ) ? ( n5071 ) : ( iram_188 ) ;
assign n23295 = wr_addr[7:7] ;
assign n23296 =  ( n23295 ) == ( bv_1_0_n53 )  ;
assign n23297 =  ( wr_addr ) == ( bv_8_188_n445 )  ;
assign n23298 =  ( n23296 ) & (n23297 )  ;
assign n23299 =  ( n23298 ) & (wr )  ;
assign n23300 =  ( n23299 ) ? ( n5096 ) : ( iram_188 ) ;
assign n23301 = wr_addr[7:7] ;
assign n23302 =  ( n23301 ) == ( bv_1_0_n53 )  ;
assign n23303 =  ( wr_addr ) == ( bv_8_188_n445 )  ;
assign n23304 =  ( n23302 ) & (n23303 )  ;
assign n23305 =  ( n23304 ) & (wr )  ;
assign n23306 =  ( n23305 ) ? ( n5123 ) : ( iram_188 ) ;
assign n23307 = wr_addr[7:7] ;
assign n23308 =  ( n23307 ) == ( bv_1_0_n53 )  ;
assign n23309 =  ( wr_addr ) == ( bv_8_188_n445 )  ;
assign n23310 =  ( n23308 ) & (n23309 )  ;
assign n23311 =  ( n23310 ) & (wr )  ;
assign n23312 =  ( n23311 ) ? ( n5165 ) : ( iram_188 ) ;
assign n23313 = wr_addr[7:7] ;
assign n23314 =  ( n23313 ) == ( bv_1_0_n53 )  ;
assign n23315 =  ( wr_addr ) == ( bv_8_188_n445 )  ;
assign n23316 =  ( n23314 ) & (n23315 )  ;
assign n23317 =  ( n23316 ) & (wr )  ;
assign n23318 =  ( n23317 ) ? ( n5204 ) : ( iram_188 ) ;
assign n23319 = wr_addr[7:7] ;
assign n23320 =  ( n23319 ) == ( bv_1_0_n53 )  ;
assign n23321 =  ( wr_addr ) == ( bv_8_188_n445 )  ;
assign n23322 =  ( n23320 ) & (n23321 )  ;
assign n23323 =  ( n23322 ) & (wr )  ;
assign n23324 =  ( n23323 ) ? ( n5262 ) : ( iram_188 ) ;
assign n23325 = wr_addr[7:7] ;
assign n23326 =  ( n23325 ) == ( bv_1_0_n53 )  ;
assign n23327 =  ( wr_addr ) == ( bv_8_188_n445 )  ;
assign n23328 =  ( n23326 ) & (n23327 )  ;
assign n23329 =  ( n23328 ) & (wr )  ;
assign n23330 =  ( n23329 ) ? ( n5298 ) : ( iram_188 ) ;
assign n23331 = wr_addr[7:7] ;
assign n23332 =  ( n23331 ) == ( bv_1_0_n53 )  ;
assign n23333 =  ( wr_addr ) == ( bv_8_188_n445 )  ;
assign n23334 =  ( n23332 ) & (n23333 )  ;
assign n23335 =  ( n23334 ) & (wr )  ;
assign n23336 =  ( n23335 ) ? ( n5325 ) : ( iram_188 ) ;
assign n23337 = wr_addr[7:7] ;
assign n23338 =  ( n23337 ) == ( bv_1_0_n53 )  ;
assign n23339 =  ( wr_addr ) == ( bv_8_189_n447 )  ;
assign n23340 =  ( n23338 ) & (n23339 )  ;
assign n23341 =  ( n23340 ) & (wr )  ;
assign n23342 =  ( n23341 ) ? ( n4782 ) : ( iram_189 ) ;
assign n23343 = wr_addr[7:7] ;
assign n23344 =  ( n23343 ) == ( bv_1_0_n53 )  ;
assign n23345 =  ( wr_addr ) == ( bv_8_189_n447 )  ;
assign n23346 =  ( n23344 ) & (n23345 )  ;
assign n23347 =  ( n23346 ) & (wr )  ;
assign n23348 =  ( n23347 ) ? ( n4841 ) : ( iram_189 ) ;
assign n23349 = wr_addr[7:7] ;
assign n23350 =  ( n23349 ) == ( bv_1_0_n53 )  ;
assign n23351 =  ( wr_addr ) == ( bv_8_189_n447 )  ;
assign n23352 =  ( n23350 ) & (n23351 )  ;
assign n23353 =  ( n23352 ) & (wr )  ;
assign n23354 =  ( n23353 ) ? ( n5449 ) : ( iram_189 ) ;
assign n23355 = wr_addr[7:7] ;
assign n23356 =  ( n23355 ) == ( bv_1_0_n53 )  ;
assign n23357 =  ( wr_addr ) == ( bv_8_189_n447 )  ;
assign n23358 =  ( n23356 ) & (n23357 )  ;
assign n23359 =  ( n23358 ) & (wr )  ;
assign n23360 =  ( n23359 ) ? ( n4906 ) : ( iram_189 ) ;
assign n23361 = wr_addr[7:7] ;
assign n23362 =  ( n23361 ) == ( bv_1_0_n53 )  ;
assign n23363 =  ( wr_addr ) == ( bv_8_189_n447 )  ;
assign n23364 =  ( n23362 ) & (n23363 )  ;
assign n23365 =  ( n23364 ) & (wr )  ;
assign n23366 =  ( n23365 ) ? ( n5485 ) : ( iram_189 ) ;
assign n23367 = wr_addr[7:7] ;
assign n23368 =  ( n23367 ) == ( bv_1_0_n53 )  ;
assign n23369 =  ( wr_addr ) == ( bv_8_189_n447 )  ;
assign n23370 =  ( n23368 ) & (n23369 )  ;
assign n23371 =  ( n23370 ) & (wr )  ;
assign n23372 =  ( n23371 ) ? ( n5512 ) : ( iram_189 ) ;
assign n23373 = wr_addr[7:7] ;
assign n23374 =  ( n23373 ) == ( bv_1_0_n53 )  ;
assign n23375 =  ( wr_addr ) == ( bv_8_189_n447 )  ;
assign n23376 =  ( n23374 ) & (n23375 )  ;
assign n23377 =  ( n23376 ) & (wr )  ;
assign n23378 =  ( n23377 ) ? ( bv_8_0_n69 ) : ( iram_189 ) ;
assign n23379 = wr_addr[7:7] ;
assign n23380 =  ( n23379 ) == ( bv_1_0_n53 )  ;
assign n23381 =  ( wr_addr ) == ( bv_8_189_n447 )  ;
assign n23382 =  ( n23380 ) & (n23381 )  ;
assign n23383 =  ( n23382 ) & (wr )  ;
assign n23384 =  ( n23383 ) ? ( n5071 ) : ( iram_189 ) ;
assign n23385 = wr_addr[7:7] ;
assign n23386 =  ( n23385 ) == ( bv_1_0_n53 )  ;
assign n23387 =  ( wr_addr ) == ( bv_8_189_n447 )  ;
assign n23388 =  ( n23386 ) & (n23387 )  ;
assign n23389 =  ( n23388 ) & (wr )  ;
assign n23390 =  ( n23389 ) ? ( n5096 ) : ( iram_189 ) ;
assign n23391 = wr_addr[7:7] ;
assign n23392 =  ( n23391 ) == ( bv_1_0_n53 )  ;
assign n23393 =  ( wr_addr ) == ( bv_8_189_n447 )  ;
assign n23394 =  ( n23392 ) & (n23393 )  ;
assign n23395 =  ( n23394 ) & (wr )  ;
assign n23396 =  ( n23395 ) ? ( n5123 ) : ( iram_189 ) ;
assign n23397 = wr_addr[7:7] ;
assign n23398 =  ( n23397 ) == ( bv_1_0_n53 )  ;
assign n23399 =  ( wr_addr ) == ( bv_8_189_n447 )  ;
assign n23400 =  ( n23398 ) & (n23399 )  ;
assign n23401 =  ( n23400 ) & (wr )  ;
assign n23402 =  ( n23401 ) ? ( n5165 ) : ( iram_189 ) ;
assign n23403 = wr_addr[7:7] ;
assign n23404 =  ( n23403 ) == ( bv_1_0_n53 )  ;
assign n23405 =  ( wr_addr ) == ( bv_8_189_n447 )  ;
assign n23406 =  ( n23404 ) & (n23405 )  ;
assign n23407 =  ( n23406 ) & (wr )  ;
assign n23408 =  ( n23407 ) ? ( n5204 ) : ( iram_189 ) ;
assign n23409 = wr_addr[7:7] ;
assign n23410 =  ( n23409 ) == ( bv_1_0_n53 )  ;
assign n23411 =  ( wr_addr ) == ( bv_8_189_n447 )  ;
assign n23412 =  ( n23410 ) & (n23411 )  ;
assign n23413 =  ( n23412 ) & (wr )  ;
assign n23414 =  ( n23413 ) ? ( n5262 ) : ( iram_189 ) ;
assign n23415 = wr_addr[7:7] ;
assign n23416 =  ( n23415 ) == ( bv_1_0_n53 )  ;
assign n23417 =  ( wr_addr ) == ( bv_8_189_n447 )  ;
assign n23418 =  ( n23416 ) & (n23417 )  ;
assign n23419 =  ( n23418 ) & (wr )  ;
assign n23420 =  ( n23419 ) ? ( n5298 ) : ( iram_189 ) ;
assign n23421 = wr_addr[7:7] ;
assign n23422 =  ( n23421 ) == ( bv_1_0_n53 )  ;
assign n23423 =  ( wr_addr ) == ( bv_8_189_n447 )  ;
assign n23424 =  ( n23422 ) & (n23423 )  ;
assign n23425 =  ( n23424 ) & (wr )  ;
assign n23426 =  ( n23425 ) ? ( n5325 ) : ( iram_189 ) ;
assign n23427 = wr_addr[7:7] ;
assign n23428 =  ( n23427 ) == ( bv_1_0_n53 )  ;
assign n23429 =  ( wr_addr ) == ( bv_8_190_n449 )  ;
assign n23430 =  ( n23428 ) & (n23429 )  ;
assign n23431 =  ( n23430 ) & (wr )  ;
assign n23432 =  ( n23431 ) ? ( n4782 ) : ( iram_190 ) ;
assign n23433 = wr_addr[7:7] ;
assign n23434 =  ( n23433 ) == ( bv_1_0_n53 )  ;
assign n23435 =  ( wr_addr ) == ( bv_8_190_n449 )  ;
assign n23436 =  ( n23434 ) & (n23435 )  ;
assign n23437 =  ( n23436 ) & (wr )  ;
assign n23438 =  ( n23437 ) ? ( n4841 ) : ( iram_190 ) ;
assign n23439 = wr_addr[7:7] ;
assign n23440 =  ( n23439 ) == ( bv_1_0_n53 )  ;
assign n23441 =  ( wr_addr ) == ( bv_8_190_n449 )  ;
assign n23442 =  ( n23440 ) & (n23441 )  ;
assign n23443 =  ( n23442 ) & (wr )  ;
assign n23444 =  ( n23443 ) ? ( n5449 ) : ( iram_190 ) ;
assign n23445 = wr_addr[7:7] ;
assign n23446 =  ( n23445 ) == ( bv_1_0_n53 )  ;
assign n23447 =  ( wr_addr ) == ( bv_8_190_n449 )  ;
assign n23448 =  ( n23446 ) & (n23447 )  ;
assign n23449 =  ( n23448 ) & (wr )  ;
assign n23450 =  ( n23449 ) ? ( n4906 ) : ( iram_190 ) ;
assign n23451 = wr_addr[7:7] ;
assign n23452 =  ( n23451 ) == ( bv_1_0_n53 )  ;
assign n23453 =  ( wr_addr ) == ( bv_8_190_n449 )  ;
assign n23454 =  ( n23452 ) & (n23453 )  ;
assign n23455 =  ( n23454 ) & (wr )  ;
assign n23456 =  ( n23455 ) ? ( n5485 ) : ( iram_190 ) ;
assign n23457 = wr_addr[7:7] ;
assign n23458 =  ( n23457 ) == ( bv_1_0_n53 )  ;
assign n23459 =  ( wr_addr ) == ( bv_8_190_n449 )  ;
assign n23460 =  ( n23458 ) & (n23459 )  ;
assign n23461 =  ( n23460 ) & (wr )  ;
assign n23462 =  ( n23461 ) ? ( n5512 ) : ( iram_190 ) ;
assign n23463 = wr_addr[7:7] ;
assign n23464 =  ( n23463 ) == ( bv_1_0_n53 )  ;
assign n23465 =  ( wr_addr ) == ( bv_8_190_n449 )  ;
assign n23466 =  ( n23464 ) & (n23465 )  ;
assign n23467 =  ( n23466 ) & (wr )  ;
assign n23468 =  ( n23467 ) ? ( bv_8_0_n69 ) : ( iram_190 ) ;
assign n23469 = wr_addr[7:7] ;
assign n23470 =  ( n23469 ) == ( bv_1_0_n53 )  ;
assign n23471 =  ( wr_addr ) == ( bv_8_190_n449 )  ;
assign n23472 =  ( n23470 ) & (n23471 )  ;
assign n23473 =  ( n23472 ) & (wr )  ;
assign n23474 =  ( n23473 ) ? ( n5071 ) : ( iram_190 ) ;
assign n23475 = wr_addr[7:7] ;
assign n23476 =  ( n23475 ) == ( bv_1_0_n53 )  ;
assign n23477 =  ( wr_addr ) == ( bv_8_190_n449 )  ;
assign n23478 =  ( n23476 ) & (n23477 )  ;
assign n23479 =  ( n23478 ) & (wr )  ;
assign n23480 =  ( n23479 ) ? ( n5096 ) : ( iram_190 ) ;
assign n23481 = wr_addr[7:7] ;
assign n23482 =  ( n23481 ) == ( bv_1_0_n53 )  ;
assign n23483 =  ( wr_addr ) == ( bv_8_190_n449 )  ;
assign n23484 =  ( n23482 ) & (n23483 )  ;
assign n23485 =  ( n23484 ) & (wr )  ;
assign n23486 =  ( n23485 ) ? ( n5123 ) : ( iram_190 ) ;
assign n23487 = wr_addr[7:7] ;
assign n23488 =  ( n23487 ) == ( bv_1_0_n53 )  ;
assign n23489 =  ( wr_addr ) == ( bv_8_190_n449 )  ;
assign n23490 =  ( n23488 ) & (n23489 )  ;
assign n23491 =  ( n23490 ) & (wr )  ;
assign n23492 =  ( n23491 ) ? ( n5165 ) : ( iram_190 ) ;
assign n23493 = wr_addr[7:7] ;
assign n23494 =  ( n23493 ) == ( bv_1_0_n53 )  ;
assign n23495 =  ( wr_addr ) == ( bv_8_190_n449 )  ;
assign n23496 =  ( n23494 ) & (n23495 )  ;
assign n23497 =  ( n23496 ) & (wr )  ;
assign n23498 =  ( n23497 ) ? ( n5204 ) : ( iram_190 ) ;
assign n23499 = wr_addr[7:7] ;
assign n23500 =  ( n23499 ) == ( bv_1_0_n53 )  ;
assign n23501 =  ( wr_addr ) == ( bv_8_190_n449 )  ;
assign n23502 =  ( n23500 ) & (n23501 )  ;
assign n23503 =  ( n23502 ) & (wr )  ;
assign n23504 =  ( n23503 ) ? ( n5262 ) : ( iram_190 ) ;
assign n23505 = wr_addr[7:7] ;
assign n23506 =  ( n23505 ) == ( bv_1_0_n53 )  ;
assign n23507 =  ( wr_addr ) == ( bv_8_190_n449 )  ;
assign n23508 =  ( n23506 ) & (n23507 )  ;
assign n23509 =  ( n23508 ) & (wr )  ;
assign n23510 =  ( n23509 ) ? ( n5298 ) : ( iram_190 ) ;
assign n23511 = wr_addr[7:7] ;
assign n23512 =  ( n23511 ) == ( bv_1_0_n53 )  ;
assign n23513 =  ( wr_addr ) == ( bv_8_190_n449 )  ;
assign n23514 =  ( n23512 ) & (n23513 )  ;
assign n23515 =  ( n23514 ) & (wr )  ;
assign n23516 =  ( n23515 ) ? ( n5325 ) : ( iram_190 ) ;
assign n23517 = wr_addr[7:7] ;
assign n23518 =  ( n23517 ) == ( bv_1_0_n53 )  ;
assign n23519 =  ( wr_addr ) == ( bv_8_191_n451 )  ;
assign n23520 =  ( n23518 ) & (n23519 )  ;
assign n23521 =  ( n23520 ) & (wr )  ;
assign n23522 =  ( n23521 ) ? ( n4782 ) : ( iram_191 ) ;
assign n23523 = wr_addr[7:7] ;
assign n23524 =  ( n23523 ) == ( bv_1_0_n53 )  ;
assign n23525 =  ( wr_addr ) == ( bv_8_191_n451 )  ;
assign n23526 =  ( n23524 ) & (n23525 )  ;
assign n23527 =  ( n23526 ) & (wr )  ;
assign n23528 =  ( n23527 ) ? ( n4841 ) : ( iram_191 ) ;
assign n23529 = wr_addr[7:7] ;
assign n23530 =  ( n23529 ) == ( bv_1_0_n53 )  ;
assign n23531 =  ( wr_addr ) == ( bv_8_191_n451 )  ;
assign n23532 =  ( n23530 ) & (n23531 )  ;
assign n23533 =  ( n23532 ) & (wr )  ;
assign n23534 =  ( n23533 ) ? ( n5449 ) : ( iram_191 ) ;
assign n23535 = wr_addr[7:7] ;
assign n23536 =  ( n23535 ) == ( bv_1_0_n53 )  ;
assign n23537 =  ( wr_addr ) == ( bv_8_191_n451 )  ;
assign n23538 =  ( n23536 ) & (n23537 )  ;
assign n23539 =  ( n23538 ) & (wr )  ;
assign n23540 =  ( n23539 ) ? ( n4906 ) : ( iram_191 ) ;
assign n23541 = wr_addr[7:7] ;
assign n23542 =  ( n23541 ) == ( bv_1_0_n53 )  ;
assign n23543 =  ( wr_addr ) == ( bv_8_191_n451 )  ;
assign n23544 =  ( n23542 ) & (n23543 )  ;
assign n23545 =  ( n23544 ) & (wr )  ;
assign n23546 =  ( n23545 ) ? ( n5485 ) : ( iram_191 ) ;
assign n23547 = wr_addr[7:7] ;
assign n23548 =  ( n23547 ) == ( bv_1_0_n53 )  ;
assign n23549 =  ( wr_addr ) == ( bv_8_191_n451 )  ;
assign n23550 =  ( n23548 ) & (n23549 )  ;
assign n23551 =  ( n23550 ) & (wr )  ;
assign n23552 =  ( n23551 ) ? ( n5512 ) : ( iram_191 ) ;
assign n23553 = wr_addr[7:7] ;
assign n23554 =  ( n23553 ) == ( bv_1_0_n53 )  ;
assign n23555 =  ( wr_addr ) == ( bv_8_191_n451 )  ;
assign n23556 =  ( n23554 ) & (n23555 )  ;
assign n23557 =  ( n23556 ) & (wr )  ;
assign n23558 =  ( n23557 ) ? ( bv_8_0_n69 ) : ( iram_191 ) ;
assign n23559 = wr_addr[7:7] ;
assign n23560 =  ( n23559 ) == ( bv_1_0_n53 )  ;
assign n23561 =  ( wr_addr ) == ( bv_8_191_n451 )  ;
assign n23562 =  ( n23560 ) & (n23561 )  ;
assign n23563 =  ( n23562 ) & (wr )  ;
assign n23564 =  ( n23563 ) ? ( n5071 ) : ( iram_191 ) ;
assign n23565 = wr_addr[7:7] ;
assign n23566 =  ( n23565 ) == ( bv_1_0_n53 )  ;
assign n23567 =  ( wr_addr ) == ( bv_8_191_n451 )  ;
assign n23568 =  ( n23566 ) & (n23567 )  ;
assign n23569 =  ( n23568 ) & (wr )  ;
assign n23570 =  ( n23569 ) ? ( n5096 ) : ( iram_191 ) ;
assign n23571 = wr_addr[7:7] ;
assign n23572 =  ( n23571 ) == ( bv_1_0_n53 )  ;
assign n23573 =  ( wr_addr ) == ( bv_8_191_n451 )  ;
assign n23574 =  ( n23572 ) & (n23573 )  ;
assign n23575 =  ( n23574 ) & (wr )  ;
assign n23576 =  ( n23575 ) ? ( n5123 ) : ( iram_191 ) ;
assign n23577 = wr_addr[7:7] ;
assign n23578 =  ( n23577 ) == ( bv_1_0_n53 )  ;
assign n23579 =  ( wr_addr ) == ( bv_8_191_n451 )  ;
assign n23580 =  ( n23578 ) & (n23579 )  ;
assign n23581 =  ( n23580 ) & (wr )  ;
assign n23582 =  ( n23581 ) ? ( n5165 ) : ( iram_191 ) ;
assign n23583 = wr_addr[7:7] ;
assign n23584 =  ( n23583 ) == ( bv_1_0_n53 )  ;
assign n23585 =  ( wr_addr ) == ( bv_8_191_n451 )  ;
assign n23586 =  ( n23584 ) & (n23585 )  ;
assign n23587 =  ( n23586 ) & (wr )  ;
assign n23588 =  ( n23587 ) ? ( n5204 ) : ( iram_191 ) ;
assign n23589 = wr_addr[7:7] ;
assign n23590 =  ( n23589 ) == ( bv_1_0_n53 )  ;
assign n23591 =  ( wr_addr ) == ( bv_8_191_n451 )  ;
assign n23592 =  ( n23590 ) & (n23591 )  ;
assign n23593 =  ( n23592 ) & (wr )  ;
assign n23594 =  ( n23593 ) ? ( n5262 ) : ( iram_191 ) ;
assign n23595 = wr_addr[7:7] ;
assign n23596 =  ( n23595 ) == ( bv_1_0_n53 )  ;
assign n23597 =  ( wr_addr ) == ( bv_8_191_n451 )  ;
assign n23598 =  ( n23596 ) & (n23597 )  ;
assign n23599 =  ( n23598 ) & (wr )  ;
assign n23600 =  ( n23599 ) ? ( n5298 ) : ( iram_191 ) ;
assign n23601 = wr_addr[7:7] ;
assign n23602 =  ( n23601 ) == ( bv_1_0_n53 )  ;
assign n23603 =  ( wr_addr ) == ( bv_8_191_n451 )  ;
assign n23604 =  ( n23602 ) & (n23603 )  ;
assign n23605 =  ( n23604 ) & (wr )  ;
assign n23606 =  ( n23605 ) ? ( n5325 ) : ( iram_191 ) ;
assign n23607 = wr_addr[7:7] ;
assign n23608 =  ( n23607 ) == ( bv_1_0_n53 )  ;
assign n23609 =  ( wr_addr ) == ( bv_8_192_n453 )  ;
assign n23610 =  ( n23608 ) & (n23609 )  ;
assign n23611 =  ( n23610 ) & (wr )  ;
assign n23612 =  ( n23611 ) ? ( n4782 ) : ( iram_192 ) ;
assign n23613 = wr_addr[7:7] ;
assign n23614 =  ( n23613 ) == ( bv_1_0_n53 )  ;
assign n23615 =  ( wr_addr ) == ( bv_8_192_n453 )  ;
assign n23616 =  ( n23614 ) & (n23615 )  ;
assign n23617 =  ( n23616 ) & (wr )  ;
assign n23618 =  ( n23617 ) ? ( n4841 ) : ( iram_192 ) ;
assign n23619 = wr_addr[7:7] ;
assign n23620 =  ( n23619 ) == ( bv_1_0_n53 )  ;
assign n23621 =  ( wr_addr ) == ( bv_8_192_n453 )  ;
assign n23622 =  ( n23620 ) & (n23621 )  ;
assign n23623 =  ( n23622 ) & (wr )  ;
assign n23624 =  ( n23623 ) ? ( n5449 ) : ( iram_192 ) ;
assign n23625 = wr_addr[7:7] ;
assign n23626 =  ( n23625 ) == ( bv_1_0_n53 )  ;
assign n23627 =  ( wr_addr ) == ( bv_8_192_n453 )  ;
assign n23628 =  ( n23626 ) & (n23627 )  ;
assign n23629 =  ( n23628 ) & (wr )  ;
assign n23630 =  ( n23629 ) ? ( n4906 ) : ( iram_192 ) ;
assign n23631 = wr_addr[7:7] ;
assign n23632 =  ( n23631 ) == ( bv_1_0_n53 )  ;
assign n23633 =  ( wr_addr ) == ( bv_8_192_n453 )  ;
assign n23634 =  ( n23632 ) & (n23633 )  ;
assign n23635 =  ( n23634 ) & (wr )  ;
assign n23636 =  ( n23635 ) ? ( n5485 ) : ( iram_192 ) ;
assign n23637 = wr_addr[7:7] ;
assign n23638 =  ( n23637 ) == ( bv_1_0_n53 )  ;
assign n23639 =  ( wr_addr ) == ( bv_8_192_n453 )  ;
assign n23640 =  ( n23638 ) & (n23639 )  ;
assign n23641 =  ( n23640 ) & (wr )  ;
assign n23642 =  ( n23641 ) ? ( n5512 ) : ( iram_192 ) ;
assign n23643 = wr_addr[7:7] ;
assign n23644 =  ( n23643 ) == ( bv_1_0_n53 )  ;
assign n23645 =  ( wr_addr ) == ( bv_8_192_n453 )  ;
assign n23646 =  ( n23644 ) & (n23645 )  ;
assign n23647 =  ( n23646 ) & (wr )  ;
assign n23648 =  ( n23647 ) ? ( bv_8_0_n69 ) : ( iram_192 ) ;
assign n23649 = wr_addr[7:7] ;
assign n23650 =  ( n23649 ) == ( bv_1_0_n53 )  ;
assign n23651 =  ( wr_addr ) == ( bv_8_192_n453 )  ;
assign n23652 =  ( n23650 ) & (n23651 )  ;
assign n23653 =  ( n23652 ) & (wr )  ;
assign n23654 =  ( n23653 ) ? ( n5071 ) : ( iram_192 ) ;
assign n23655 = wr_addr[7:7] ;
assign n23656 =  ( n23655 ) == ( bv_1_0_n53 )  ;
assign n23657 =  ( wr_addr ) == ( bv_8_192_n453 )  ;
assign n23658 =  ( n23656 ) & (n23657 )  ;
assign n23659 =  ( n23658 ) & (wr )  ;
assign n23660 =  ( n23659 ) ? ( n5096 ) : ( iram_192 ) ;
assign n23661 = wr_addr[7:7] ;
assign n23662 =  ( n23661 ) == ( bv_1_0_n53 )  ;
assign n23663 =  ( wr_addr ) == ( bv_8_192_n453 )  ;
assign n23664 =  ( n23662 ) & (n23663 )  ;
assign n23665 =  ( n23664 ) & (wr )  ;
assign n23666 =  ( n23665 ) ? ( n5123 ) : ( iram_192 ) ;
assign n23667 = wr_addr[7:7] ;
assign n23668 =  ( n23667 ) == ( bv_1_0_n53 )  ;
assign n23669 =  ( wr_addr ) == ( bv_8_192_n453 )  ;
assign n23670 =  ( n23668 ) & (n23669 )  ;
assign n23671 =  ( n23670 ) & (wr )  ;
assign n23672 =  ( n23671 ) ? ( n5165 ) : ( iram_192 ) ;
assign n23673 = wr_addr[7:7] ;
assign n23674 =  ( n23673 ) == ( bv_1_0_n53 )  ;
assign n23675 =  ( wr_addr ) == ( bv_8_192_n453 )  ;
assign n23676 =  ( n23674 ) & (n23675 )  ;
assign n23677 =  ( n23676 ) & (wr )  ;
assign n23678 =  ( n23677 ) ? ( n5204 ) : ( iram_192 ) ;
assign n23679 = wr_addr[7:7] ;
assign n23680 =  ( n23679 ) == ( bv_1_0_n53 )  ;
assign n23681 =  ( wr_addr ) == ( bv_8_192_n453 )  ;
assign n23682 =  ( n23680 ) & (n23681 )  ;
assign n23683 =  ( n23682 ) & (wr )  ;
assign n23684 =  ( n23683 ) ? ( n5262 ) : ( iram_192 ) ;
assign n23685 = wr_addr[7:7] ;
assign n23686 =  ( n23685 ) == ( bv_1_0_n53 )  ;
assign n23687 =  ( wr_addr ) == ( bv_8_192_n453 )  ;
assign n23688 =  ( n23686 ) & (n23687 )  ;
assign n23689 =  ( n23688 ) & (wr )  ;
assign n23690 =  ( n23689 ) ? ( n5298 ) : ( iram_192 ) ;
assign n23691 = wr_addr[7:7] ;
assign n23692 =  ( n23691 ) == ( bv_1_0_n53 )  ;
assign n23693 =  ( wr_addr ) == ( bv_8_192_n453 )  ;
assign n23694 =  ( n23692 ) & (n23693 )  ;
assign n23695 =  ( n23694 ) & (wr )  ;
assign n23696 =  ( n23695 ) ? ( n5325 ) : ( iram_192 ) ;
assign n23697 = wr_addr[7:7] ;
assign n23698 =  ( n23697 ) == ( bv_1_0_n53 )  ;
assign n23699 =  ( wr_addr ) == ( bv_8_193_n455 )  ;
assign n23700 =  ( n23698 ) & (n23699 )  ;
assign n23701 =  ( n23700 ) & (wr )  ;
assign n23702 =  ( n23701 ) ? ( n4782 ) : ( iram_193 ) ;
assign n23703 = wr_addr[7:7] ;
assign n23704 =  ( n23703 ) == ( bv_1_0_n53 )  ;
assign n23705 =  ( wr_addr ) == ( bv_8_193_n455 )  ;
assign n23706 =  ( n23704 ) & (n23705 )  ;
assign n23707 =  ( n23706 ) & (wr )  ;
assign n23708 =  ( n23707 ) ? ( n4841 ) : ( iram_193 ) ;
assign n23709 = wr_addr[7:7] ;
assign n23710 =  ( n23709 ) == ( bv_1_0_n53 )  ;
assign n23711 =  ( wr_addr ) == ( bv_8_193_n455 )  ;
assign n23712 =  ( n23710 ) & (n23711 )  ;
assign n23713 =  ( n23712 ) & (wr )  ;
assign n23714 =  ( n23713 ) ? ( n5449 ) : ( iram_193 ) ;
assign n23715 = wr_addr[7:7] ;
assign n23716 =  ( n23715 ) == ( bv_1_0_n53 )  ;
assign n23717 =  ( wr_addr ) == ( bv_8_193_n455 )  ;
assign n23718 =  ( n23716 ) & (n23717 )  ;
assign n23719 =  ( n23718 ) & (wr )  ;
assign n23720 =  ( n23719 ) ? ( n4906 ) : ( iram_193 ) ;
assign n23721 = wr_addr[7:7] ;
assign n23722 =  ( n23721 ) == ( bv_1_0_n53 )  ;
assign n23723 =  ( wr_addr ) == ( bv_8_193_n455 )  ;
assign n23724 =  ( n23722 ) & (n23723 )  ;
assign n23725 =  ( n23724 ) & (wr )  ;
assign n23726 =  ( n23725 ) ? ( n5485 ) : ( iram_193 ) ;
assign n23727 = wr_addr[7:7] ;
assign n23728 =  ( n23727 ) == ( bv_1_0_n53 )  ;
assign n23729 =  ( wr_addr ) == ( bv_8_193_n455 )  ;
assign n23730 =  ( n23728 ) & (n23729 )  ;
assign n23731 =  ( n23730 ) & (wr )  ;
assign n23732 =  ( n23731 ) ? ( n5512 ) : ( iram_193 ) ;
assign n23733 = wr_addr[7:7] ;
assign n23734 =  ( n23733 ) == ( bv_1_0_n53 )  ;
assign n23735 =  ( wr_addr ) == ( bv_8_193_n455 )  ;
assign n23736 =  ( n23734 ) & (n23735 )  ;
assign n23737 =  ( n23736 ) & (wr )  ;
assign n23738 =  ( n23737 ) ? ( bv_8_0_n69 ) : ( iram_193 ) ;
assign n23739 = wr_addr[7:7] ;
assign n23740 =  ( n23739 ) == ( bv_1_0_n53 )  ;
assign n23741 =  ( wr_addr ) == ( bv_8_193_n455 )  ;
assign n23742 =  ( n23740 ) & (n23741 )  ;
assign n23743 =  ( n23742 ) & (wr )  ;
assign n23744 =  ( n23743 ) ? ( n5071 ) : ( iram_193 ) ;
assign n23745 = wr_addr[7:7] ;
assign n23746 =  ( n23745 ) == ( bv_1_0_n53 )  ;
assign n23747 =  ( wr_addr ) == ( bv_8_193_n455 )  ;
assign n23748 =  ( n23746 ) & (n23747 )  ;
assign n23749 =  ( n23748 ) & (wr )  ;
assign n23750 =  ( n23749 ) ? ( n5096 ) : ( iram_193 ) ;
assign n23751 = wr_addr[7:7] ;
assign n23752 =  ( n23751 ) == ( bv_1_0_n53 )  ;
assign n23753 =  ( wr_addr ) == ( bv_8_193_n455 )  ;
assign n23754 =  ( n23752 ) & (n23753 )  ;
assign n23755 =  ( n23754 ) & (wr )  ;
assign n23756 =  ( n23755 ) ? ( n5123 ) : ( iram_193 ) ;
assign n23757 = wr_addr[7:7] ;
assign n23758 =  ( n23757 ) == ( bv_1_0_n53 )  ;
assign n23759 =  ( wr_addr ) == ( bv_8_193_n455 )  ;
assign n23760 =  ( n23758 ) & (n23759 )  ;
assign n23761 =  ( n23760 ) & (wr )  ;
assign n23762 =  ( n23761 ) ? ( n5165 ) : ( iram_193 ) ;
assign n23763 = wr_addr[7:7] ;
assign n23764 =  ( n23763 ) == ( bv_1_0_n53 )  ;
assign n23765 =  ( wr_addr ) == ( bv_8_193_n455 )  ;
assign n23766 =  ( n23764 ) & (n23765 )  ;
assign n23767 =  ( n23766 ) & (wr )  ;
assign n23768 =  ( n23767 ) ? ( n5204 ) : ( iram_193 ) ;
assign n23769 = wr_addr[7:7] ;
assign n23770 =  ( n23769 ) == ( bv_1_0_n53 )  ;
assign n23771 =  ( wr_addr ) == ( bv_8_193_n455 )  ;
assign n23772 =  ( n23770 ) & (n23771 )  ;
assign n23773 =  ( n23772 ) & (wr )  ;
assign n23774 =  ( n23773 ) ? ( n5262 ) : ( iram_193 ) ;
assign n23775 = wr_addr[7:7] ;
assign n23776 =  ( n23775 ) == ( bv_1_0_n53 )  ;
assign n23777 =  ( wr_addr ) == ( bv_8_193_n455 )  ;
assign n23778 =  ( n23776 ) & (n23777 )  ;
assign n23779 =  ( n23778 ) & (wr )  ;
assign n23780 =  ( n23779 ) ? ( n5298 ) : ( iram_193 ) ;
assign n23781 = wr_addr[7:7] ;
assign n23782 =  ( n23781 ) == ( bv_1_0_n53 )  ;
assign n23783 =  ( wr_addr ) == ( bv_8_193_n455 )  ;
assign n23784 =  ( n23782 ) & (n23783 )  ;
assign n23785 =  ( n23784 ) & (wr )  ;
assign n23786 =  ( n23785 ) ? ( n5325 ) : ( iram_193 ) ;
assign n23787 = wr_addr[7:7] ;
assign n23788 =  ( n23787 ) == ( bv_1_0_n53 )  ;
assign n23789 =  ( wr_addr ) == ( bv_8_194_n457 )  ;
assign n23790 =  ( n23788 ) & (n23789 )  ;
assign n23791 =  ( n23790 ) & (wr )  ;
assign n23792 =  ( n23791 ) ? ( n4782 ) : ( iram_194 ) ;
assign n23793 = wr_addr[7:7] ;
assign n23794 =  ( n23793 ) == ( bv_1_0_n53 )  ;
assign n23795 =  ( wr_addr ) == ( bv_8_194_n457 )  ;
assign n23796 =  ( n23794 ) & (n23795 )  ;
assign n23797 =  ( n23796 ) & (wr )  ;
assign n23798 =  ( n23797 ) ? ( n4841 ) : ( iram_194 ) ;
assign n23799 = wr_addr[7:7] ;
assign n23800 =  ( n23799 ) == ( bv_1_0_n53 )  ;
assign n23801 =  ( wr_addr ) == ( bv_8_194_n457 )  ;
assign n23802 =  ( n23800 ) & (n23801 )  ;
assign n23803 =  ( n23802 ) & (wr )  ;
assign n23804 =  ( n23803 ) ? ( n5449 ) : ( iram_194 ) ;
assign n23805 = wr_addr[7:7] ;
assign n23806 =  ( n23805 ) == ( bv_1_0_n53 )  ;
assign n23807 =  ( wr_addr ) == ( bv_8_194_n457 )  ;
assign n23808 =  ( n23806 ) & (n23807 )  ;
assign n23809 =  ( n23808 ) & (wr )  ;
assign n23810 =  ( n23809 ) ? ( n4906 ) : ( iram_194 ) ;
assign n23811 = wr_addr[7:7] ;
assign n23812 =  ( n23811 ) == ( bv_1_0_n53 )  ;
assign n23813 =  ( wr_addr ) == ( bv_8_194_n457 )  ;
assign n23814 =  ( n23812 ) & (n23813 )  ;
assign n23815 =  ( n23814 ) & (wr )  ;
assign n23816 =  ( n23815 ) ? ( n5485 ) : ( iram_194 ) ;
assign n23817 = wr_addr[7:7] ;
assign n23818 =  ( n23817 ) == ( bv_1_0_n53 )  ;
assign n23819 =  ( wr_addr ) == ( bv_8_194_n457 )  ;
assign n23820 =  ( n23818 ) & (n23819 )  ;
assign n23821 =  ( n23820 ) & (wr )  ;
assign n23822 =  ( n23821 ) ? ( n5512 ) : ( iram_194 ) ;
assign n23823 = wr_addr[7:7] ;
assign n23824 =  ( n23823 ) == ( bv_1_0_n53 )  ;
assign n23825 =  ( wr_addr ) == ( bv_8_194_n457 )  ;
assign n23826 =  ( n23824 ) & (n23825 )  ;
assign n23827 =  ( n23826 ) & (wr )  ;
assign n23828 =  ( n23827 ) ? ( bv_8_0_n69 ) : ( iram_194 ) ;
assign n23829 = wr_addr[7:7] ;
assign n23830 =  ( n23829 ) == ( bv_1_0_n53 )  ;
assign n23831 =  ( wr_addr ) == ( bv_8_194_n457 )  ;
assign n23832 =  ( n23830 ) & (n23831 )  ;
assign n23833 =  ( n23832 ) & (wr )  ;
assign n23834 =  ( n23833 ) ? ( n5071 ) : ( iram_194 ) ;
assign n23835 = wr_addr[7:7] ;
assign n23836 =  ( n23835 ) == ( bv_1_0_n53 )  ;
assign n23837 =  ( wr_addr ) == ( bv_8_194_n457 )  ;
assign n23838 =  ( n23836 ) & (n23837 )  ;
assign n23839 =  ( n23838 ) & (wr )  ;
assign n23840 =  ( n23839 ) ? ( n5096 ) : ( iram_194 ) ;
assign n23841 = wr_addr[7:7] ;
assign n23842 =  ( n23841 ) == ( bv_1_0_n53 )  ;
assign n23843 =  ( wr_addr ) == ( bv_8_194_n457 )  ;
assign n23844 =  ( n23842 ) & (n23843 )  ;
assign n23845 =  ( n23844 ) & (wr )  ;
assign n23846 =  ( n23845 ) ? ( n5123 ) : ( iram_194 ) ;
assign n23847 = wr_addr[7:7] ;
assign n23848 =  ( n23847 ) == ( bv_1_0_n53 )  ;
assign n23849 =  ( wr_addr ) == ( bv_8_194_n457 )  ;
assign n23850 =  ( n23848 ) & (n23849 )  ;
assign n23851 =  ( n23850 ) & (wr )  ;
assign n23852 =  ( n23851 ) ? ( n5165 ) : ( iram_194 ) ;
assign n23853 = wr_addr[7:7] ;
assign n23854 =  ( n23853 ) == ( bv_1_0_n53 )  ;
assign n23855 =  ( wr_addr ) == ( bv_8_194_n457 )  ;
assign n23856 =  ( n23854 ) & (n23855 )  ;
assign n23857 =  ( n23856 ) & (wr )  ;
assign n23858 =  ( n23857 ) ? ( n5204 ) : ( iram_194 ) ;
assign n23859 = wr_addr[7:7] ;
assign n23860 =  ( n23859 ) == ( bv_1_0_n53 )  ;
assign n23861 =  ( wr_addr ) == ( bv_8_194_n457 )  ;
assign n23862 =  ( n23860 ) & (n23861 )  ;
assign n23863 =  ( n23862 ) & (wr )  ;
assign n23864 =  ( n23863 ) ? ( n5262 ) : ( iram_194 ) ;
assign n23865 = wr_addr[7:7] ;
assign n23866 =  ( n23865 ) == ( bv_1_0_n53 )  ;
assign n23867 =  ( wr_addr ) == ( bv_8_194_n457 )  ;
assign n23868 =  ( n23866 ) & (n23867 )  ;
assign n23869 =  ( n23868 ) & (wr )  ;
assign n23870 =  ( n23869 ) ? ( n5298 ) : ( iram_194 ) ;
assign n23871 = wr_addr[7:7] ;
assign n23872 =  ( n23871 ) == ( bv_1_0_n53 )  ;
assign n23873 =  ( wr_addr ) == ( bv_8_194_n457 )  ;
assign n23874 =  ( n23872 ) & (n23873 )  ;
assign n23875 =  ( n23874 ) & (wr )  ;
assign n23876 =  ( n23875 ) ? ( n5325 ) : ( iram_194 ) ;
assign n23877 = wr_addr[7:7] ;
assign n23878 =  ( n23877 ) == ( bv_1_0_n53 )  ;
assign n23879 =  ( wr_addr ) == ( bv_8_195_n459 )  ;
assign n23880 =  ( n23878 ) & (n23879 )  ;
assign n23881 =  ( n23880 ) & (wr )  ;
assign n23882 =  ( n23881 ) ? ( n4782 ) : ( iram_195 ) ;
assign n23883 = wr_addr[7:7] ;
assign n23884 =  ( n23883 ) == ( bv_1_0_n53 )  ;
assign n23885 =  ( wr_addr ) == ( bv_8_195_n459 )  ;
assign n23886 =  ( n23884 ) & (n23885 )  ;
assign n23887 =  ( n23886 ) & (wr )  ;
assign n23888 =  ( n23887 ) ? ( n4841 ) : ( iram_195 ) ;
assign n23889 = wr_addr[7:7] ;
assign n23890 =  ( n23889 ) == ( bv_1_0_n53 )  ;
assign n23891 =  ( wr_addr ) == ( bv_8_195_n459 )  ;
assign n23892 =  ( n23890 ) & (n23891 )  ;
assign n23893 =  ( n23892 ) & (wr )  ;
assign n23894 =  ( n23893 ) ? ( n5449 ) : ( iram_195 ) ;
assign n23895 = wr_addr[7:7] ;
assign n23896 =  ( n23895 ) == ( bv_1_0_n53 )  ;
assign n23897 =  ( wr_addr ) == ( bv_8_195_n459 )  ;
assign n23898 =  ( n23896 ) & (n23897 )  ;
assign n23899 =  ( n23898 ) & (wr )  ;
assign n23900 =  ( n23899 ) ? ( n4906 ) : ( iram_195 ) ;
assign n23901 = wr_addr[7:7] ;
assign n23902 =  ( n23901 ) == ( bv_1_0_n53 )  ;
assign n23903 =  ( wr_addr ) == ( bv_8_195_n459 )  ;
assign n23904 =  ( n23902 ) & (n23903 )  ;
assign n23905 =  ( n23904 ) & (wr )  ;
assign n23906 =  ( n23905 ) ? ( n5485 ) : ( iram_195 ) ;
assign n23907 = wr_addr[7:7] ;
assign n23908 =  ( n23907 ) == ( bv_1_0_n53 )  ;
assign n23909 =  ( wr_addr ) == ( bv_8_195_n459 )  ;
assign n23910 =  ( n23908 ) & (n23909 )  ;
assign n23911 =  ( n23910 ) & (wr )  ;
assign n23912 =  ( n23911 ) ? ( n5512 ) : ( iram_195 ) ;
assign n23913 = wr_addr[7:7] ;
assign n23914 =  ( n23913 ) == ( bv_1_0_n53 )  ;
assign n23915 =  ( wr_addr ) == ( bv_8_195_n459 )  ;
assign n23916 =  ( n23914 ) & (n23915 )  ;
assign n23917 =  ( n23916 ) & (wr )  ;
assign n23918 =  ( n23917 ) ? ( bv_8_0_n69 ) : ( iram_195 ) ;
assign n23919 = wr_addr[7:7] ;
assign n23920 =  ( n23919 ) == ( bv_1_0_n53 )  ;
assign n23921 =  ( wr_addr ) == ( bv_8_195_n459 )  ;
assign n23922 =  ( n23920 ) & (n23921 )  ;
assign n23923 =  ( n23922 ) & (wr )  ;
assign n23924 =  ( n23923 ) ? ( n5071 ) : ( iram_195 ) ;
assign n23925 = wr_addr[7:7] ;
assign n23926 =  ( n23925 ) == ( bv_1_0_n53 )  ;
assign n23927 =  ( wr_addr ) == ( bv_8_195_n459 )  ;
assign n23928 =  ( n23926 ) & (n23927 )  ;
assign n23929 =  ( n23928 ) & (wr )  ;
assign n23930 =  ( n23929 ) ? ( n5096 ) : ( iram_195 ) ;
assign n23931 = wr_addr[7:7] ;
assign n23932 =  ( n23931 ) == ( bv_1_0_n53 )  ;
assign n23933 =  ( wr_addr ) == ( bv_8_195_n459 )  ;
assign n23934 =  ( n23932 ) & (n23933 )  ;
assign n23935 =  ( n23934 ) & (wr )  ;
assign n23936 =  ( n23935 ) ? ( n5123 ) : ( iram_195 ) ;
assign n23937 = wr_addr[7:7] ;
assign n23938 =  ( n23937 ) == ( bv_1_0_n53 )  ;
assign n23939 =  ( wr_addr ) == ( bv_8_195_n459 )  ;
assign n23940 =  ( n23938 ) & (n23939 )  ;
assign n23941 =  ( n23940 ) & (wr )  ;
assign n23942 =  ( n23941 ) ? ( n5165 ) : ( iram_195 ) ;
assign n23943 = wr_addr[7:7] ;
assign n23944 =  ( n23943 ) == ( bv_1_0_n53 )  ;
assign n23945 =  ( wr_addr ) == ( bv_8_195_n459 )  ;
assign n23946 =  ( n23944 ) & (n23945 )  ;
assign n23947 =  ( n23946 ) & (wr )  ;
assign n23948 =  ( n23947 ) ? ( n5204 ) : ( iram_195 ) ;
assign n23949 = wr_addr[7:7] ;
assign n23950 =  ( n23949 ) == ( bv_1_0_n53 )  ;
assign n23951 =  ( wr_addr ) == ( bv_8_195_n459 )  ;
assign n23952 =  ( n23950 ) & (n23951 )  ;
assign n23953 =  ( n23952 ) & (wr )  ;
assign n23954 =  ( n23953 ) ? ( n5262 ) : ( iram_195 ) ;
assign n23955 = wr_addr[7:7] ;
assign n23956 =  ( n23955 ) == ( bv_1_0_n53 )  ;
assign n23957 =  ( wr_addr ) == ( bv_8_195_n459 )  ;
assign n23958 =  ( n23956 ) & (n23957 )  ;
assign n23959 =  ( n23958 ) & (wr )  ;
assign n23960 =  ( n23959 ) ? ( n5298 ) : ( iram_195 ) ;
assign n23961 = wr_addr[7:7] ;
assign n23962 =  ( n23961 ) == ( bv_1_0_n53 )  ;
assign n23963 =  ( wr_addr ) == ( bv_8_195_n459 )  ;
assign n23964 =  ( n23962 ) & (n23963 )  ;
assign n23965 =  ( n23964 ) & (wr )  ;
assign n23966 =  ( n23965 ) ? ( n5325 ) : ( iram_195 ) ;
assign n23967 = wr_addr[7:7] ;
assign n23968 =  ( n23967 ) == ( bv_1_0_n53 )  ;
assign n23969 =  ( wr_addr ) == ( bv_8_196_n461 )  ;
assign n23970 =  ( n23968 ) & (n23969 )  ;
assign n23971 =  ( n23970 ) & (wr )  ;
assign n23972 =  ( n23971 ) ? ( n4782 ) : ( iram_196 ) ;
assign n23973 = wr_addr[7:7] ;
assign n23974 =  ( n23973 ) == ( bv_1_0_n53 )  ;
assign n23975 =  ( wr_addr ) == ( bv_8_196_n461 )  ;
assign n23976 =  ( n23974 ) & (n23975 )  ;
assign n23977 =  ( n23976 ) & (wr )  ;
assign n23978 =  ( n23977 ) ? ( n4841 ) : ( iram_196 ) ;
assign n23979 = wr_addr[7:7] ;
assign n23980 =  ( n23979 ) == ( bv_1_0_n53 )  ;
assign n23981 =  ( wr_addr ) == ( bv_8_196_n461 )  ;
assign n23982 =  ( n23980 ) & (n23981 )  ;
assign n23983 =  ( n23982 ) & (wr )  ;
assign n23984 =  ( n23983 ) ? ( n5449 ) : ( iram_196 ) ;
assign n23985 = wr_addr[7:7] ;
assign n23986 =  ( n23985 ) == ( bv_1_0_n53 )  ;
assign n23987 =  ( wr_addr ) == ( bv_8_196_n461 )  ;
assign n23988 =  ( n23986 ) & (n23987 )  ;
assign n23989 =  ( n23988 ) & (wr )  ;
assign n23990 =  ( n23989 ) ? ( n4906 ) : ( iram_196 ) ;
assign n23991 = wr_addr[7:7] ;
assign n23992 =  ( n23991 ) == ( bv_1_0_n53 )  ;
assign n23993 =  ( wr_addr ) == ( bv_8_196_n461 )  ;
assign n23994 =  ( n23992 ) & (n23993 )  ;
assign n23995 =  ( n23994 ) & (wr )  ;
assign n23996 =  ( n23995 ) ? ( n5485 ) : ( iram_196 ) ;
assign n23997 = wr_addr[7:7] ;
assign n23998 =  ( n23997 ) == ( bv_1_0_n53 )  ;
assign n23999 =  ( wr_addr ) == ( bv_8_196_n461 )  ;
assign n24000 =  ( n23998 ) & (n23999 )  ;
assign n24001 =  ( n24000 ) & (wr )  ;
assign n24002 =  ( n24001 ) ? ( n5512 ) : ( iram_196 ) ;
assign n24003 = wr_addr[7:7] ;
assign n24004 =  ( n24003 ) == ( bv_1_0_n53 )  ;
assign n24005 =  ( wr_addr ) == ( bv_8_196_n461 )  ;
assign n24006 =  ( n24004 ) & (n24005 )  ;
assign n24007 =  ( n24006 ) & (wr )  ;
assign n24008 =  ( n24007 ) ? ( bv_8_0_n69 ) : ( iram_196 ) ;
assign n24009 = wr_addr[7:7] ;
assign n24010 =  ( n24009 ) == ( bv_1_0_n53 )  ;
assign n24011 =  ( wr_addr ) == ( bv_8_196_n461 )  ;
assign n24012 =  ( n24010 ) & (n24011 )  ;
assign n24013 =  ( n24012 ) & (wr )  ;
assign n24014 =  ( n24013 ) ? ( n5071 ) : ( iram_196 ) ;
assign n24015 = wr_addr[7:7] ;
assign n24016 =  ( n24015 ) == ( bv_1_0_n53 )  ;
assign n24017 =  ( wr_addr ) == ( bv_8_196_n461 )  ;
assign n24018 =  ( n24016 ) & (n24017 )  ;
assign n24019 =  ( n24018 ) & (wr )  ;
assign n24020 =  ( n24019 ) ? ( n5096 ) : ( iram_196 ) ;
assign n24021 = wr_addr[7:7] ;
assign n24022 =  ( n24021 ) == ( bv_1_0_n53 )  ;
assign n24023 =  ( wr_addr ) == ( bv_8_196_n461 )  ;
assign n24024 =  ( n24022 ) & (n24023 )  ;
assign n24025 =  ( n24024 ) & (wr )  ;
assign n24026 =  ( n24025 ) ? ( n5123 ) : ( iram_196 ) ;
assign n24027 = wr_addr[7:7] ;
assign n24028 =  ( n24027 ) == ( bv_1_0_n53 )  ;
assign n24029 =  ( wr_addr ) == ( bv_8_196_n461 )  ;
assign n24030 =  ( n24028 ) & (n24029 )  ;
assign n24031 =  ( n24030 ) & (wr )  ;
assign n24032 =  ( n24031 ) ? ( n5165 ) : ( iram_196 ) ;
assign n24033 = wr_addr[7:7] ;
assign n24034 =  ( n24033 ) == ( bv_1_0_n53 )  ;
assign n24035 =  ( wr_addr ) == ( bv_8_196_n461 )  ;
assign n24036 =  ( n24034 ) & (n24035 )  ;
assign n24037 =  ( n24036 ) & (wr )  ;
assign n24038 =  ( n24037 ) ? ( n5204 ) : ( iram_196 ) ;
assign n24039 = wr_addr[7:7] ;
assign n24040 =  ( n24039 ) == ( bv_1_0_n53 )  ;
assign n24041 =  ( wr_addr ) == ( bv_8_196_n461 )  ;
assign n24042 =  ( n24040 ) & (n24041 )  ;
assign n24043 =  ( n24042 ) & (wr )  ;
assign n24044 =  ( n24043 ) ? ( n5262 ) : ( iram_196 ) ;
assign n24045 = wr_addr[7:7] ;
assign n24046 =  ( n24045 ) == ( bv_1_0_n53 )  ;
assign n24047 =  ( wr_addr ) == ( bv_8_196_n461 )  ;
assign n24048 =  ( n24046 ) & (n24047 )  ;
assign n24049 =  ( n24048 ) & (wr )  ;
assign n24050 =  ( n24049 ) ? ( n5298 ) : ( iram_196 ) ;
assign n24051 = wr_addr[7:7] ;
assign n24052 =  ( n24051 ) == ( bv_1_0_n53 )  ;
assign n24053 =  ( wr_addr ) == ( bv_8_196_n461 )  ;
assign n24054 =  ( n24052 ) & (n24053 )  ;
assign n24055 =  ( n24054 ) & (wr )  ;
assign n24056 =  ( n24055 ) ? ( n5325 ) : ( iram_196 ) ;
assign n24057 = wr_addr[7:7] ;
assign n24058 =  ( n24057 ) == ( bv_1_0_n53 )  ;
assign n24059 =  ( wr_addr ) == ( bv_8_197_n463 )  ;
assign n24060 =  ( n24058 ) & (n24059 )  ;
assign n24061 =  ( n24060 ) & (wr )  ;
assign n24062 =  ( n24061 ) ? ( n4782 ) : ( iram_197 ) ;
assign n24063 = wr_addr[7:7] ;
assign n24064 =  ( n24063 ) == ( bv_1_0_n53 )  ;
assign n24065 =  ( wr_addr ) == ( bv_8_197_n463 )  ;
assign n24066 =  ( n24064 ) & (n24065 )  ;
assign n24067 =  ( n24066 ) & (wr )  ;
assign n24068 =  ( n24067 ) ? ( n4841 ) : ( iram_197 ) ;
assign n24069 = wr_addr[7:7] ;
assign n24070 =  ( n24069 ) == ( bv_1_0_n53 )  ;
assign n24071 =  ( wr_addr ) == ( bv_8_197_n463 )  ;
assign n24072 =  ( n24070 ) & (n24071 )  ;
assign n24073 =  ( n24072 ) & (wr )  ;
assign n24074 =  ( n24073 ) ? ( n5449 ) : ( iram_197 ) ;
assign n24075 = wr_addr[7:7] ;
assign n24076 =  ( n24075 ) == ( bv_1_0_n53 )  ;
assign n24077 =  ( wr_addr ) == ( bv_8_197_n463 )  ;
assign n24078 =  ( n24076 ) & (n24077 )  ;
assign n24079 =  ( n24078 ) & (wr )  ;
assign n24080 =  ( n24079 ) ? ( n4906 ) : ( iram_197 ) ;
assign n24081 = wr_addr[7:7] ;
assign n24082 =  ( n24081 ) == ( bv_1_0_n53 )  ;
assign n24083 =  ( wr_addr ) == ( bv_8_197_n463 )  ;
assign n24084 =  ( n24082 ) & (n24083 )  ;
assign n24085 =  ( n24084 ) & (wr )  ;
assign n24086 =  ( n24085 ) ? ( n5485 ) : ( iram_197 ) ;
assign n24087 = wr_addr[7:7] ;
assign n24088 =  ( n24087 ) == ( bv_1_0_n53 )  ;
assign n24089 =  ( wr_addr ) == ( bv_8_197_n463 )  ;
assign n24090 =  ( n24088 ) & (n24089 )  ;
assign n24091 =  ( n24090 ) & (wr )  ;
assign n24092 =  ( n24091 ) ? ( n5512 ) : ( iram_197 ) ;
assign n24093 = wr_addr[7:7] ;
assign n24094 =  ( n24093 ) == ( bv_1_0_n53 )  ;
assign n24095 =  ( wr_addr ) == ( bv_8_197_n463 )  ;
assign n24096 =  ( n24094 ) & (n24095 )  ;
assign n24097 =  ( n24096 ) & (wr )  ;
assign n24098 =  ( n24097 ) ? ( bv_8_0_n69 ) : ( iram_197 ) ;
assign n24099 = wr_addr[7:7] ;
assign n24100 =  ( n24099 ) == ( bv_1_0_n53 )  ;
assign n24101 =  ( wr_addr ) == ( bv_8_197_n463 )  ;
assign n24102 =  ( n24100 ) & (n24101 )  ;
assign n24103 =  ( n24102 ) & (wr )  ;
assign n24104 =  ( n24103 ) ? ( n5071 ) : ( iram_197 ) ;
assign n24105 = wr_addr[7:7] ;
assign n24106 =  ( n24105 ) == ( bv_1_0_n53 )  ;
assign n24107 =  ( wr_addr ) == ( bv_8_197_n463 )  ;
assign n24108 =  ( n24106 ) & (n24107 )  ;
assign n24109 =  ( n24108 ) & (wr )  ;
assign n24110 =  ( n24109 ) ? ( n5096 ) : ( iram_197 ) ;
assign n24111 = wr_addr[7:7] ;
assign n24112 =  ( n24111 ) == ( bv_1_0_n53 )  ;
assign n24113 =  ( wr_addr ) == ( bv_8_197_n463 )  ;
assign n24114 =  ( n24112 ) & (n24113 )  ;
assign n24115 =  ( n24114 ) & (wr )  ;
assign n24116 =  ( n24115 ) ? ( n5123 ) : ( iram_197 ) ;
assign n24117 = wr_addr[7:7] ;
assign n24118 =  ( n24117 ) == ( bv_1_0_n53 )  ;
assign n24119 =  ( wr_addr ) == ( bv_8_197_n463 )  ;
assign n24120 =  ( n24118 ) & (n24119 )  ;
assign n24121 =  ( n24120 ) & (wr )  ;
assign n24122 =  ( n24121 ) ? ( n5165 ) : ( iram_197 ) ;
assign n24123 = wr_addr[7:7] ;
assign n24124 =  ( n24123 ) == ( bv_1_0_n53 )  ;
assign n24125 =  ( wr_addr ) == ( bv_8_197_n463 )  ;
assign n24126 =  ( n24124 ) & (n24125 )  ;
assign n24127 =  ( n24126 ) & (wr )  ;
assign n24128 =  ( n24127 ) ? ( n5204 ) : ( iram_197 ) ;
assign n24129 = wr_addr[7:7] ;
assign n24130 =  ( n24129 ) == ( bv_1_0_n53 )  ;
assign n24131 =  ( wr_addr ) == ( bv_8_197_n463 )  ;
assign n24132 =  ( n24130 ) & (n24131 )  ;
assign n24133 =  ( n24132 ) & (wr )  ;
assign n24134 =  ( n24133 ) ? ( n5262 ) : ( iram_197 ) ;
assign n24135 = wr_addr[7:7] ;
assign n24136 =  ( n24135 ) == ( bv_1_0_n53 )  ;
assign n24137 =  ( wr_addr ) == ( bv_8_197_n463 )  ;
assign n24138 =  ( n24136 ) & (n24137 )  ;
assign n24139 =  ( n24138 ) & (wr )  ;
assign n24140 =  ( n24139 ) ? ( n5298 ) : ( iram_197 ) ;
assign n24141 = wr_addr[7:7] ;
assign n24142 =  ( n24141 ) == ( bv_1_0_n53 )  ;
assign n24143 =  ( wr_addr ) == ( bv_8_197_n463 )  ;
assign n24144 =  ( n24142 ) & (n24143 )  ;
assign n24145 =  ( n24144 ) & (wr )  ;
assign n24146 =  ( n24145 ) ? ( n5325 ) : ( iram_197 ) ;
assign n24147 = wr_addr[7:7] ;
assign n24148 =  ( n24147 ) == ( bv_1_0_n53 )  ;
assign n24149 =  ( wr_addr ) == ( bv_8_198_n465 )  ;
assign n24150 =  ( n24148 ) & (n24149 )  ;
assign n24151 =  ( n24150 ) & (wr )  ;
assign n24152 =  ( n24151 ) ? ( n4782 ) : ( iram_198 ) ;
assign n24153 = wr_addr[7:7] ;
assign n24154 =  ( n24153 ) == ( bv_1_0_n53 )  ;
assign n24155 =  ( wr_addr ) == ( bv_8_198_n465 )  ;
assign n24156 =  ( n24154 ) & (n24155 )  ;
assign n24157 =  ( n24156 ) & (wr )  ;
assign n24158 =  ( n24157 ) ? ( n4841 ) : ( iram_198 ) ;
assign n24159 = wr_addr[7:7] ;
assign n24160 =  ( n24159 ) == ( bv_1_0_n53 )  ;
assign n24161 =  ( wr_addr ) == ( bv_8_198_n465 )  ;
assign n24162 =  ( n24160 ) & (n24161 )  ;
assign n24163 =  ( n24162 ) & (wr )  ;
assign n24164 =  ( n24163 ) ? ( n5449 ) : ( iram_198 ) ;
assign n24165 = wr_addr[7:7] ;
assign n24166 =  ( n24165 ) == ( bv_1_0_n53 )  ;
assign n24167 =  ( wr_addr ) == ( bv_8_198_n465 )  ;
assign n24168 =  ( n24166 ) & (n24167 )  ;
assign n24169 =  ( n24168 ) & (wr )  ;
assign n24170 =  ( n24169 ) ? ( n4906 ) : ( iram_198 ) ;
assign n24171 = wr_addr[7:7] ;
assign n24172 =  ( n24171 ) == ( bv_1_0_n53 )  ;
assign n24173 =  ( wr_addr ) == ( bv_8_198_n465 )  ;
assign n24174 =  ( n24172 ) & (n24173 )  ;
assign n24175 =  ( n24174 ) & (wr )  ;
assign n24176 =  ( n24175 ) ? ( n5485 ) : ( iram_198 ) ;
assign n24177 = wr_addr[7:7] ;
assign n24178 =  ( n24177 ) == ( bv_1_0_n53 )  ;
assign n24179 =  ( wr_addr ) == ( bv_8_198_n465 )  ;
assign n24180 =  ( n24178 ) & (n24179 )  ;
assign n24181 =  ( n24180 ) & (wr )  ;
assign n24182 =  ( n24181 ) ? ( n5512 ) : ( iram_198 ) ;
assign n24183 = wr_addr[7:7] ;
assign n24184 =  ( n24183 ) == ( bv_1_0_n53 )  ;
assign n24185 =  ( wr_addr ) == ( bv_8_198_n465 )  ;
assign n24186 =  ( n24184 ) & (n24185 )  ;
assign n24187 =  ( n24186 ) & (wr )  ;
assign n24188 =  ( n24187 ) ? ( bv_8_0_n69 ) : ( iram_198 ) ;
assign n24189 = wr_addr[7:7] ;
assign n24190 =  ( n24189 ) == ( bv_1_0_n53 )  ;
assign n24191 =  ( wr_addr ) == ( bv_8_198_n465 )  ;
assign n24192 =  ( n24190 ) & (n24191 )  ;
assign n24193 =  ( n24192 ) & (wr )  ;
assign n24194 =  ( n24193 ) ? ( n5071 ) : ( iram_198 ) ;
assign n24195 = wr_addr[7:7] ;
assign n24196 =  ( n24195 ) == ( bv_1_0_n53 )  ;
assign n24197 =  ( wr_addr ) == ( bv_8_198_n465 )  ;
assign n24198 =  ( n24196 ) & (n24197 )  ;
assign n24199 =  ( n24198 ) & (wr )  ;
assign n24200 =  ( n24199 ) ? ( n5096 ) : ( iram_198 ) ;
assign n24201 = wr_addr[7:7] ;
assign n24202 =  ( n24201 ) == ( bv_1_0_n53 )  ;
assign n24203 =  ( wr_addr ) == ( bv_8_198_n465 )  ;
assign n24204 =  ( n24202 ) & (n24203 )  ;
assign n24205 =  ( n24204 ) & (wr )  ;
assign n24206 =  ( n24205 ) ? ( n5123 ) : ( iram_198 ) ;
assign n24207 = wr_addr[7:7] ;
assign n24208 =  ( n24207 ) == ( bv_1_0_n53 )  ;
assign n24209 =  ( wr_addr ) == ( bv_8_198_n465 )  ;
assign n24210 =  ( n24208 ) & (n24209 )  ;
assign n24211 =  ( n24210 ) & (wr )  ;
assign n24212 =  ( n24211 ) ? ( n5165 ) : ( iram_198 ) ;
assign n24213 = wr_addr[7:7] ;
assign n24214 =  ( n24213 ) == ( bv_1_0_n53 )  ;
assign n24215 =  ( wr_addr ) == ( bv_8_198_n465 )  ;
assign n24216 =  ( n24214 ) & (n24215 )  ;
assign n24217 =  ( n24216 ) & (wr )  ;
assign n24218 =  ( n24217 ) ? ( n5204 ) : ( iram_198 ) ;
assign n24219 = wr_addr[7:7] ;
assign n24220 =  ( n24219 ) == ( bv_1_0_n53 )  ;
assign n24221 =  ( wr_addr ) == ( bv_8_198_n465 )  ;
assign n24222 =  ( n24220 ) & (n24221 )  ;
assign n24223 =  ( n24222 ) & (wr )  ;
assign n24224 =  ( n24223 ) ? ( n5262 ) : ( iram_198 ) ;
assign n24225 = wr_addr[7:7] ;
assign n24226 =  ( n24225 ) == ( bv_1_0_n53 )  ;
assign n24227 =  ( wr_addr ) == ( bv_8_198_n465 )  ;
assign n24228 =  ( n24226 ) & (n24227 )  ;
assign n24229 =  ( n24228 ) & (wr )  ;
assign n24230 =  ( n24229 ) ? ( n5298 ) : ( iram_198 ) ;
assign n24231 = wr_addr[7:7] ;
assign n24232 =  ( n24231 ) == ( bv_1_0_n53 )  ;
assign n24233 =  ( wr_addr ) == ( bv_8_198_n465 )  ;
assign n24234 =  ( n24232 ) & (n24233 )  ;
assign n24235 =  ( n24234 ) & (wr )  ;
assign n24236 =  ( n24235 ) ? ( n5325 ) : ( iram_198 ) ;
assign n24237 = wr_addr[7:7] ;
assign n24238 =  ( n24237 ) == ( bv_1_0_n53 )  ;
assign n24239 =  ( wr_addr ) == ( bv_8_199_n467 )  ;
assign n24240 =  ( n24238 ) & (n24239 )  ;
assign n24241 =  ( n24240 ) & (wr )  ;
assign n24242 =  ( n24241 ) ? ( n4782 ) : ( iram_199 ) ;
assign n24243 = wr_addr[7:7] ;
assign n24244 =  ( n24243 ) == ( bv_1_0_n53 )  ;
assign n24245 =  ( wr_addr ) == ( bv_8_199_n467 )  ;
assign n24246 =  ( n24244 ) & (n24245 )  ;
assign n24247 =  ( n24246 ) & (wr )  ;
assign n24248 =  ( n24247 ) ? ( n4841 ) : ( iram_199 ) ;
assign n24249 = wr_addr[7:7] ;
assign n24250 =  ( n24249 ) == ( bv_1_0_n53 )  ;
assign n24251 =  ( wr_addr ) == ( bv_8_199_n467 )  ;
assign n24252 =  ( n24250 ) & (n24251 )  ;
assign n24253 =  ( n24252 ) & (wr )  ;
assign n24254 =  ( n24253 ) ? ( n5449 ) : ( iram_199 ) ;
assign n24255 = wr_addr[7:7] ;
assign n24256 =  ( n24255 ) == ( bv_1_0_n53 )  ;
assign n24257 =  ( wr_addr ) == ( bv_8_199_n467 )  ;
assign n24258 =  ( n24256 ) & (n24257 )  ;
assign n24259 =  ( n24258 ) & (wr )  ;
assign n24260 =  ( n24259 ) ? ( n4906 ) : ( iram_199 ) ;
assign n24261 = wr_addr[7:7] ;
assign n24262 =  ( n24261 ) == ( bv_1_0_n53 )  ;
assign n24263 =  ( wr_addr ) == ( bv_8_199_n467 )  ;
assign n24264 =  ( n24262 ) & (n24263 )  ;
assign n24265 =  ( n24264 ) & (wr )  ;
assign n24266 =  ( n24265 ) ? ( n5485 ) : ( iram_199 ) ;
assign n24267 = wr_addr[7:7] ;
assign n24268 =  ( n24267 ) == ( bv_1_0_n53 )  ;
assign n24269 =  ( wr_addr ) == ( bv_8_199_n467 )  ;
assign n24270 =  ( n24268 ) & (n24269 )  ;
assign n24271 =  ( n24270 ) & (wr )  ;
assign n24272 =  ( n24271 ) ? ( n5512 ) : ( iram_199 ) ;
assign n24273 = wr_addr[7:7] ;
assign n24274 =  ( n24273 ) == ( bv_1_0_n53 )  ;
assign n24275 =  ( wr_addr ) == ( bv_8_199_n467 )  ;
assign n24276 =  ( n24274 ) & (n24275 )  ;
assign n24277 =  ( n24276 ) & (wr )  ;
assign n24278 =  ( n24277 ) ? ( bv_8_0_n69 ) : ( iram_199 ) ;
assign n24279 = wr_addr[7:7] ;
assign n24280 =  ( n24279 ) == ( bv_1_0_n53 )  ;
assign n24281 =  ( wr_addr ) == ( bv_8_199_n467 )  ;
assign n24282 =  ( n24280 ) & (n24281 )  ;
assign n24283 =  ( n24282 ) & (wr )  ;
assign n24284 =  ( n24283 ) ? ( n5071 ) : ( iram_199 ) ;
assign n24285 = wr_addr[7:7] ;
assign n24286 =  ( n24285 ) == ( bv_1_0_n53 )  ;
assign n24287 =  ( wr_addr ) == ( bv_8_199_n467 )  ;
assign n24288 =  ( n24286 ) & (n24287 )  ;
assign n24289 =  ( n24288 ) & (wr )  ;
assign n24290 =  ( n24289 ) ? ( n5096 ) : ( iram_199 ) ;
assign n24291 = wr_addr[7:7] ;
assign n24292 =  ( n24291 ) == ( bv_1_0_n53 )  ;
assign n24293 =  ( wr_addr ) == ( bv_8_199_n467 )  ;
assign n24294 =  ( n24292 ) & (n24293 )  ;
assign n24295 =  ( n24294 ) & (wr )  ;
assign n24296 =  ( n24295 ) ? ( n5123 ) : ( iram_199 ) ;
assign n24297 = wr_addr[7:7] ;
assign n24298 =  ( n24297 ) == ( bv_1_0_n53 )  ;
assign n24299 =  ( wr_addr ) == ( bv_8_199_n467 )  ;
assign n24300 =  ( n24298 ) & (n24299 )  ;
assign n24301 =  ( n24300 ) & (wr )  ;
assign n24302 =  ( n24301 ) ? ( n5165 ) : ( iram_199 ) ;
assign n24303 = wr_addr[7:7] ;
assign n24304 =  ( n24303 ) == ( bv_1_0_n53 )  ;
assign n24305 =  ( wr_addr ) == ( bv_8_199_n467 )  ;
assign n24306 =  ( n24304 ) & (n24305 )  ;
assign n24307 =  ( n24306 ) & (wr )  ;
assign n24308 =  ( n24307 ) ? ( n5204 ) : ( iram_199 ) ;
assign n24309 = wr_addr[7:7] ;
assign n24310 =  ( n24309 ) == ( bv_1_0_n53 )  ;
assign n24311 =  ( wr_addr ) == ( bv_8_199_n467 )  ;
assign n24312 =  ( n24310 ) & (n24311 )  ;
assign n24313 =  ( n24312 ) & (wr )  ;
assign n24314 =  ( n24313 ) ? ( n5262 ) : ( iram_199 ) ;
assign n24315 = wr_addr[7:7] ;
assign n24316 =  ( n24315 ) == ( bv_1_0_n53 )  ;
assign n24317 =  ( wr_addr ) == ( bv_8_199_n467 )  ;
assign n24318 =  ( n24316 ) & (n24317 )  ;
assign n24319 =  ( n24318 ) & (wr )  ;
assign n24320 =  ( n24319 ) ? ( n5298 ) : ( iram_199 ) ;
assign n24321 = wr_addr[7:7] ;
assign n24322 =  ( n24321 ) == ( bv_1_0_n53 )  ;
assign n24323 =  ( wr_addr ) == ( bv_8_199_n467 )  ;
assign n24324 =  ( n24322 ) & (n24323 )  ;
assign n24325 =  ( n24324 ) & (wr )  ;
assign n24326 =  ( n24325 ) ? ( n5325 ) : ( iram_199 ) ;
assign n24327 = wr_addr[7:7] ;
assign n24328 =  ( n24327 ) == ( bv_1_0_n53 )  ;
assign n24329 =  ( wr_addr ) == ( bv_8_200_n469 )  ;
assign n24330 =  ( n24328 ) & (n24329 )  ;
assign n24331 =  ( n24330 ) & (wr )  ;
assign n24332 =  ( n24331 ) ? ( n4782 ) : ( iram_200 ) ;
assign n24333 = wr_addr[7:7] ;
assign n24334 =  ( n24333 ) == ( bv_1_0_n53 )  ;
assign n24335 =  ( wr_addr ) == ( bv_8_200_n469 )  ;
assign n24336 =  ( n24334 ) & (n24335 )  ;
assign n24337 =  ( n24336 ) & (wr )  ;
assign n24338 =  ( n24337 ) ? ( n4841 ) : ( iram_200 ) ;
assign n24339 = wr_addr[7:7] ;
assign n24340 =  ( n24339 ) == ( bv_1_0_n53 )  ;
assign n24341 =  ( wr_addr ) == ( bv_8_200_n469 )  ;
assign n24342 =  ( n24340 ) & (n24341 )  ;
assign n24343 =  ( n24342 ) & (wr )  ;
assign n24344 =  ( n24343 ) ? ( n5449 ) : ( iram_200 ) ;
assign n24345 = wr_addr[7:7] ;
assign n24346 =  ( n24345 ) == ( bv_1_0_n53 )  ;
assign n24347 =  ( wr_addr ) == ( bv_8_200_n469 )  ;
assign n24348 =  ( n24346 ) & (n24347 )  ;
assign n24349 =  ( n24348 ) & (wr )  ;
assign n24350 =  ( n24349 ) ? ( n4906 ) : ( iram_200 ) ;
assign n24351 = wr_addr[7:7] ;
assign n24352 =  ( n24351 ) == ( bv_1_0_n53 )  ;
assign n24353 =  ( wr_addr ) == ( bv_8_200_n469 )  ;
assign n24354 =  ( n24352 ) & (n24353 )  ;
assign n24355 =  ( n24354 ) & (wr )  ;
assign n24356 =  ( n24355 ) ? ( n5485 ) : ( iram_200 ) ;
assign n24357 = wr_addr[7:7] ;
assign n24358 =  ( n24357 ) == ( bv_1_0_n53 )  ;
assign n24359 =  ( wr_addr ) == ( bv_8_200_n469 )  ;
assign n24360 =  ( n24358 ) & (n24359 )  ;
assign n24361 =  ( n24360 ) & (wr )  ;
assign n24362 =  ( n24361 ) ? ( n5512 ) : ( iram_200 ) ;
assign n24363 = wr_addr[7:7] ;
assign n24364 =  ( n24363 ) == ( bv_1_0_n53 )  ;
assign n24365 =  ( wr_addr ) == ( bv_8_200_n469 )  ;
assign n24366 =  ( n24364 ) & (n24365 )  ;
assign n24367 =  ( n24366 ) & (wr )  ;
assign n24368 =  ( n24367 ) ? ( bv_8_0_n69 ) : ( iram_200 ) ;
assign n24369 = wr_addr[7:7] ;
assign n24370 =  ( n24369 ) == ( bv_1_0_n53 )  ;
assign n24371 =  ( wr_addr ) == ( bv_8_200_n469 )  ;
assign n24372 =  ( n24370 ) & (n24371 )  ;
assign n24373 =  ( n24372 ) & (wr )  ;
assign n24374 =  ( n24373 ) ? ( n5071 ) : ( iram_200 ) ;
assign n24375 = wr_addr[7:7] ;
assign n24376 =  ( n24375 ) == ( bv_1_0_n53 )  ;
assign n24377 =  ( wr_addr ) == ( bv_8_200_n469 )  ;
assign n24378 =  ( n24376 ) & (n24377 )  ;
assign n24379 =  ( n24378 ) & (wr )  ;
assign n24380 =  ( n24379 ) ? ( n5096 ) : ( iram_200 ) ;
assign n24381 = wr_addr[7:7] ;
assign n24382 =  ( n24381 ) == ( bv_1_0_n53 )  ;
assign n24383 =  ( wr_addr ) == ( bv_8_200_n469 )  ;
assign n24384 =  ( n24382 ) & (n24383 )  ;
assign n24385 =  ( n24384 ) & (wr )  ;
assign n24386 =  ( n24385 ) ? ( n5123 ) : ( iram_200 ) ;
assign n24387 = wr_addr[7:7] ;
assign n24388 =  ( n24387 ) == ( bv_1_0_n53 )  ;
assign n24389 =  ( wr_addr ) == ( bv_8_200_n469 )  ;
assign n24390 =  ( n24388 ) & (n24389 )  ;
assign n24391 =  ( n24390 ) & (wr )  ;
assign n24392 =  ( n24391 ) ? ( n5165 ) : ( iram_200 ) ;
assign n24393 = wr_addr[7:7] ;
assign n24394 =  ( n24393 ) == ( bv_1_0_n53 )  ;
assign n24395 =  ( wr_addr ) == ( bv_8_200_n469 )  ;
assign n24396 =  ( n24394 ) & (n24395 )  ;
assign n24397 =  ( n24396 ) & (wr )  ;
assign n24398 =  ( n24397 ) ? ( n5204 ) : ( iram_200 ) ;
assign n24399 = wr_addr[7:7] ;
assign n24400 =  ( n24399 ) == ( bv_1_0_n53 )  ;
assign n24401 =  ( wr_addr ) == ( bv_8_200_n469 )  ;
assign n24402 =  ( n24400 ) & (n24401 )  ;
assign n24403 =  ( n24402 ) & (wr )  ;
assign n24404 =  ( n24403 ) ? ( n5262 ) : ( iram_200 ) ;
assign n24405 = wr_addr[7:7] ;
assign n24406 =  ( n24405 ) == ( bv_1_0_n53 )  ;
assign n24407 =  ( wr_addr ) == ( bv_8_200_n469 )  ;
assign n24408 =  ( n24406 ) & (n24407 )  ;
assign n24409 =  ( n24408 ) & (wr )  ;
assign n24410 =  ( n24409 ) ? ( n5298 ) : ( iram_200 ) ;
assign n24411 = wr_addr[7:7] ;
assign n24412 =  ( n24411 ) == ( bv_1_0_n53 )  ;
assign n24413 =  ( wr_addr ) == ( bv_8_200_n469 )  ;
assign n24414 =  ( n24412 ) & (n24413 )  ;
assign n24415 =  ( n24414 ) & (wr )  ;
assign n24416 =  ( n24415 ) ? ( n5325 ) : ( iram_200 ) ;
assign n24417 = wr_addr[7:7] ;
assign n24418 =  ( n24417 ) == ( bv_1_0_n53 )  ;
assign n24419 =  ( wr_addr ) == ( bv_8_201_n471 )  ;
assign n24420 =  ( n24418 ) & (n24419 )  ;
assign n24421 =  ( n24420 ) & (wr )  ;
assign n24422 =  ( n24421 ) ? ( n4782 ) : ( iram_201 ) ;
assign n24423 = wr_addr[7:7] ;
assign n24424 =  ( n24423 ) == ( bv_1_0_n53 )  ;
assign n24425 =  ( wr_addr ) == ( bv_8_201_n471 )  ;
assign n24426 =  ( n24424 ) & (n24425 )  ;
assign n24427 =  ( n24426 ) & (wr )  ;
assign n24428 =  ( n24427 ) ? ( n4841 ) : ( iram_201 ) ;
assign n24429 = wr_addr[7:7] ;
assign n24430 =  ( n24429 ) == ( bv_1_0_n53 )  ;
assign n24431 =  ( wr_addr ) == ( bv_8_201_n471 )  ;
assign n24432 =  ( n24430 ) & (n24431 )  ;
assign n24433 =  ( n24432 ) & (wr )  ;
assign n24434 =  ( n24433 ) ? ( n5449 ) : ( iram_201 ) ;
assign n24435 = wr_addr[7:7] ;
assign n24436 =  ( n24435 ) == ( bv_1_0_n53 )  ;
assign n24437 =  ( wr_addr ) == ( bv_8_201_n471 )  ;
assign n24438 =  ( n24436 ) & (n24437 )  ;
assign n24439 =  ( n24438 ) & (wr )  ;
assign n24440 =  ( n24439 ) ? ( n4906 ) : ( iram_201 ) ;
assign n24441 = wr_addr[7:7] ;
assign n24442 =  ( n24441 ) == ( bv_1_0_n53 )  ;
assign n24443 =  ( wr_addr ) == ( bv_8_201_n471 )  ;
assign n24444 =  ( n24442 ) & (n24443 )  ;
assign n24445 =  ( n24444 ) & (wr )  ;
assign n24446 =  ( n24445 ) ? ( n5485 ) : ( iram_201 ) ;
assign n24447 = wr_addr[7:7] ;
assign n24448 =  ( n24447 ) == ( bv_1_0_n53 )  ;
assign n24449 =  ( wr_addr ) == ( bv_8_201_n471 )  ;
assign n24450 =  ( n24448 ) & (n24449 )  ;
assign n24451 =  ( n24450 ) & (wr )  ;
assign n24452 =  ( n24451 ) ? ( n5512 ) : ( iram_201 ) ;
assign n24453 = wr_addr[7:7] ;
assign n24454 =  ( n24453 ) == ( bv_1_0_n53 )  ;
assign n24455 =  ( wr_addr ) == ( bv_8_201_n471 )  ;
assign n24456 =  ( n24454 ) & (n24455 )  ;
assign n24457 =  ( n24456 ) & (wr )  ;
assign n24458 =  ( n24457 ) ? ( bv_8_0_n69 ) : ( iram_201 ) ;
assign n24459 = wr_addr[7:7] ;
assign n24460 =  ( n24459 ) == ( bv_1_0_n53 )  ;
assign n24461 =  ( wr_addr ) == ( bv_8_201_n471 )  ;
assign n24462 =  ( n24460 ) & (n24461 )  ;
assign n24463 =  ( n24462 ) & (wr )  ;
assign n24464 =  ( n24463 ) ? ( n5071 ) : ( iram_201 ) ;
assign n24465 = wr_addr[7:7] ;
assign n24466 =  ( n24465 ) == ( bv_1_0_n53 )  ;
assign n24467 =  ( wr_addr ) == ( bv_8_201_n471 )  ;
assign n24468 =  ( n24466 ) & (n24467 )  ;
assign n24469 =  ( n24468 ) & (wr )  ;
assign n24470 =  ( n24469 ) ? ( n5096 ) : ( iram_201 ) ;
assign n24471 = wr_addr[7:7] ;
assign n24472 =  ( n24471 ) == ( bv_1_0_n53 )  ;
assign n24473 =  ( wr_addr ) == ( bv_8_201_n471 )  ;
assign n24474 =  ( n24472 ) & (n24473 )  ;
assign n24475 =  ( n24474 ) & (wr )  ;
assign n24476 =  ( n24475 ) ? ( n5123 ) : ( iram_201 ) ;
assign n24477 = wr_addr[7:7] ;
assign n24478 =  ( n24477 ) == ( bv_1_0_n53 )  ;
assign n24479 =  ( wr_addr ) == ( bv_8_201_n471 )  ;
assign n24480 =  ( n24478 ) & (n24479 )  ;
assign n24481 =  ( n24480 ) & (wr )  ;
assign n24482 =  ( n24481 ) ? ( n5165 ) : ( iram_201 ) ;
assign n24483 = wr_addr[7:7] ;
assign n24484 =  ( n24483 ) == ( bv_1_0_n53 )  ;
assign n24485 =  ( wr_addr ) == ( bv_8_201_n471 )  ;
assign n24486 =  ( n24484 ) & (n24485 )  ;
assign n24487 =  ( n24486 ) & (wr )  ;
assign n24488 =  ( n24487 ) ? ( n5204 ) : ( iram_201 ) ;
assign n24489 = wr_addr[7:7] ;
assign n24490 =  ( n24489 ) == ( bv_1_0_n53 )  ;
assign n24491 =  ( wr_addr ) == ( bv_8_201_n471 )  ;
assign n24492 =  ( n24490 ) & (n24491 )  ;
assign n24493 =  ( n24492 ) & (wr )  ;
assign n24494 =  ( n24493 ) ? ( n5262 ) : ( iram_201 ) ;
assign n24495 = wr_addr[7:7] ;
assign n24496 =  ( n24495 ) == ( bv_1_0_n53 )  ;
assign n24497 =  ( wr_addr ) == ( bv_8_201_n471 )  ;
assign n24498 =  ( n24496 ) & (n24497 )  ;
assign n24499 =  ( n24498 ) & (wr )  ;
assign n24500 =  ( n24499 ) ? ( n5298 ) : ( iram_201 ) ;
assign n24501 = wr_addr[7:7] ;
assign n24502 =  ( n24501 ) == ( bv_1_0_n53 )  ;
assign n24503 =  ( wr_addr ) == ( bv_8_201_n471 )  ;
assign n24504 =  ( n24502 ) & (n24503 )  ;
assign n24505 =  ( n24504 ) & (wr )  ;
assign n24506 =  ( n24505 ) ? ( n5325 ) : ( iram_201 ) ;
assign n24507 = wr_addr[7:7] ;
assign n24508 =  ( n24507 ) == ( bv_1_0_n53 )  ;
assign n24509 =  ( wr_addr ) == ( bv_8_202_n473 )  ;
assign n24510 =  ( n24508 ) & (n24509 )  ;
assign n24511 =  ( n24510 ) & (wr )  ;
assign n24512 =  ( n24511 ) ? ( n4782 ) : ( iram_202 ) ;
assign n24513 = wr_addr[7:7] ;
assign n24514 =  ( n24513 ) == ( bv_1_0_n53 )  ;
assign n24515 =  ( wr_addr ) == ( bv_8_202_n473 )  ;
assign n24516 =  ( n24514 ) & (n24515 )  ;
assign n24517 =  ( n24516 ) & (wr )  ;
assign n24518 =  ( n24517 ) ? ( n4841 ) : ( iram_202 ) ;
assign n24519 = wr_addr[7:7] ;
assign n24520 =  ( n24519 ) == ( bv_1_0_n53 )  ;
assign n24521 =  ( wr_addr ) == ( bv_8_202_n473 )  ;
assign n24522 =  ( n24520 ) & (n24521 )  ;
assign n24523 =  ( n24522 ) & (wr )  ;
assign n24524 =  ( n24523 ) ? ( n5449 ) : ( iram_202 ) ;
assign n24525 = wr_addr[7:7] ;
assign n24526 =  ( n24525 ) == ( bv_1_0_n53 )  ;
assign n24527 =  ( wr_addr ) == ( bv_8_202_n473 )  ;
assign n24528 =  ( n24526 ) & (n24527 )  ;
assign n24529 =  ( n24528 ) & (wr )  ;
assign n24530 =  ( n24529 ) ? ( n4906 ) : ( iram_202 ) ;
assign n24531 = wr_addr[7:7] ;
assign n24532 =  ( n24531 ) == ( bv_1_0_n53 )  ;
assign n24533 =  ( wr_addr ) == ( bv_8_202_n473 )  ;
assign n24534 =  ( n24532 ) & (n24533 )  ;
assign n24535 =  ( n24534 ) & (wr )  ;
assign n24536 =  ( n24535 ) ? ( n5485 ) : ( iram_202 ) ;
assign n24537 = wr_addr[7:7] ;
assign n24538 =  ( n24537 ) == ( bv_1_0_n53 )  ;
assign n24539 =  ( wr_addr ) == ( bv_8_202_n473 )  ;
assign n24540 =  ( n24538 ) & (n24539 )  ;
assign n24541 =  ( n24540 ) & (wr )  ;
assign n24542 =  ( n24541 ) ? ( n5512 ) : ( iram_202 ) ;
assign n24543 = wr_addr[7:7] ;
assign n24544 =  ( n24543 ) == ( bv_1_0_n53 )  ;
assign n24545 =  ( wr_addr ) == ( bv_8_202_n473 )  ;
assign n24546 =  ( n24544 ) & (n24545 )  ;
assign n24547 =  ( n24546 ) & (wr )  ;
assign n24548 =  ( n24547 ) ? ( bv_8_0_n69 ) : ( iram_202 ) ;
assign n24549 = wr_addr[7:7] ;
assign n24550 =  ( n24549 ) == ( bv_1_0_n53 )  ;
assign n24551 =  ( wr_addr ) == ( bv_8_202_n473 )  ;
assign n24552 =  ( n24550 ) & (n24551 )  ;
assign n24553 =  ( n24552 ) & (wr )  ;
assign n24554 =  ( n24553 ) ? ( n5071 ) : ( iram_202 ) ;
assign n24555 = wr_addr[7:7] ;
assign n24556 =  ( n24555 ) == ( bv_1_0_n53 )  ;
assign n24557 =  ( wr_addr ) == ( bv_8_202_n473 )  ;
assign n24558 =  ( n24556 ) & (n24557 )  ;
assign n24559 =  ( n24558 ) & (wr )  ;
assign n24560 =  ( n24559 ) ? ( n5096 ) : ( iram_202 ) ;
assign n24561 = wr_addr[7:7] ;
assign n24562 =  ( n24561 ) == ( bv_1_0_n53 )  ;
assign n24563 =  ( wr_addr ) == ( bv_8_202_n473 )  ;
assign n24564 =  ( n24562 ) & (n24563 )  ;
assign n24565 =  ( n24564 ) & (wr )  ;
assign n24566 =  ( n24565 ) ? ( n5123 ) : ( iram_202 ) ;
assign n24567 = wr_addr[7:7] ;
assign n24568 =  ( n24567 ) == ( bv_1_0_n53 )  ;
assign n24569 =  ( wr_addr ) == ( bv_8_202_n473 )  ;
assign n24570 =  ( n24568 ) & (n24569 )  ;
assign n24571 =  ( n24570 ) & (wr )  ;
assign n24572 =  ( n24571 ) ? ( n5165 ) : ( iram_202 ) ;
assign n24573 = wr_addr[7:7] ;
assign n24574 =  ( n24573 ) == ( bv_1_0_n53 )  ;
assign n24575 =  ( wr_addr ) == ( bv_8_202_n473 )  ;
assign n24576 =  ( n24574 ) & (n24575 )  ;
assign n24577 =  ( n24576 ) & (wr )  ;
assign n24578 =  ( n24577 ) ? ( n5204 ) : ( iram_202 ) ;
assign n24579 = wr_addr[7:7] ;
assign n24580 =  ( n24579 ) == ( bv_1_0_n53 )  ;
assign n24581 =  ( wr_addr ) == ( bv_8_202_n473 )  ;
assign n24582 =  ( n24580 ) & (n24581 )  ;
assign n24583 =  ( n24582 ) & (wr )  ;
assign n24584 =  ( n24583 ) ? ( n5262 ) : ( iram_202 ) ;
assign n24585 = wr_addr[7:7] ;
assign n24586 =  ( n24585 ) == ( bv_1_0_n53 )  ;
assign n24587 =  ( wr_addr ) == ( bv_8_202_n473 )  ;
assign n24588 =  ( n24586 ) & (n24587 )  ;
assign n24589 =  ( n24588 ) & (wr )  ;
assign n24590 =  ( n24589 ) ? ( n5298 ) : ( iram_202 ) ;
assign n24591 = wr_addr[7:7] ;
assign n24592 =  ( n24591 ) == ( bv_1_0_n53 )  ;
assign n24593 =  ( wr_addr ) == ( bv_8_202_n473 )  ;
assign n24594 =  ( n24592 ) & (n24593 )  ;
assign n24595 =  ( n24594 ) & (wr )  ;
assign n24596 =  ( n24595 ) ? ( n5325 ) : ( iram_202 ) ;
assign n24597 = wr_addr[7:7] ;
assign n24598 =  ( n24597 ) == ( bv_1_0_n53 )  ;
assign n24599 =  ( wr_addr ) == ( bv_8_203_n475 )  ;
assign n24600 =  ( n24598 ) & (n24599 )  ;
assign n24601 =  ( n24600 ) & (wr )  ;
assign n24602 =  ( n24601 ) ? ( n4782 ) : ( iram_203 ) ;
assign n24603 = wr_addr[7:7] ;
assign n24604 =  ( n24603 ) == ( bv_1_0_n53 )  ;
assign n24605 =  ( wr_addr ) == ( bv_8_203_n475 )  ;
assign n24606 =  ( n24604 ) & (n24605 )  ;
assign n24607 =  ( n24606 ) & (wr )  ;
assign n24608 =  ( n24607 ) ? ( n4841 ) : ( iram_203 ) ;
assign n24609 = wr_addr[7:7] ;
assign n24610 =  ( n24609 ) == ( bv_1_0_n53 )  ;
assign n24611 =  ( wr_addr ) == ( bv_8_203_n475 )  ;
assign n24612 =  ( n24610 ) & (n24611 )  ;
assign n24613 =  ( n24612 ) & (wr )  ;
assign n24614 =  ( n24613 ) ? ( n5449 ) : ( iram_203 ) ;
assign n24615 = wr_addr[7:7] ;
assign n24616 =  ( n24615 ) == ( bv_1_0_n53 )  ;
assign n24617 =  ( wr_addr ) == ( bv_8_203_n475 )  ;
assign n24618 =  ( n24616 ) & (n24617 )  ;
assign n24619 =  ( n24618 ) & (wr )  ;
assign n24620 =  ( n24619 ) ? ( n4906 ) : ( iram_203 ) ;
assign n24621 = wr_addr[7:7] ;
assign n24622 =  ( n24621 ) == ( bv_1_0_n53 )  ;
assign n24623 =  ( wr_addr ) == ( bv_8_203_n475 )  ;
assign n24624 =  ( n24622 ) & (n24623 )  ;
assign n24625 =  ( n24624 ) & (wr )  ;
assign n24626 =  ( n24625 ) ? ( n5485 ) : ( iram_203 ) ;
assign n24627 = wr_addr[7:7] ;
assign n24628 =  ( n24627 ) == ( bv_1_0_n53 )  ;
assign n24629 =  ( wr_addr ) == ( bv_8_203_n475 )  ;
assign n24630 =  ( n24628 ) & (n24629 )  ;
assign n24631 =  ( n24630 ) & (wr )  ;
assign n24632 =  ( n24631 ) ? ( n5512 ) : ( iram_203 ) ;
assign n24633 = wr_addr[7:7] ;
assign n24634 =  ( n24633 ) == ( bv_1_0_n53 )  ;
assign n24635 =  ( wr_addr ) == ( bv_8_203_n475 )  ;
assign n24636 =  ( n24634 ) & (n24635 )  ;
assign n24637 =  ( n24636 ) & (wr )  ;
assign n24638 =  ( n24637 ) ? ( bv_8_0_n69 ) : ( iram_203 ) ;
assign n24639 = wr_addr[7:7] ;
assign n24640 =  ( n24639 ) == ( bv_1_0_n53 )  ;
assign n24641 =  ( wr_addr ) == ( bv_8_203_n475 )  ;
assign n24642 =  ( n24640 ) & (n24641 )  ;
assign n24643 =  ( n24642 ) & (wr )  ;
assign n24644 =  ( n24643 ) ? ( n5071 ) : ( iram_203 ) ;
assign n24645 = wr_addr[7:7] ;
assign n24646 =  ( n24645 ) == ( bv_1_0_n53 )  ;
assign n24647 =  ( wr_addr ) == ( bv_8_203_n475 )  ;
assign n24648 =  ( n24646 ) & (n24647 )  ;
assign n24649 =  ( n24648 ) & (wr )  ;
assign n24650 =  ( n24649 ) ? ( n5096 ) : ( iram_203 ) ;
assign n24651 = wr_addr[7:7] ;
assign n24652 =  ( n24651 ) == ( bv_1_0_n53 )  ;
assign n24653 =  ( wr_addr ) == ( bv_8_203_n475 )  ;
assign n24654 =  ( n24652 ) & (n24653 )  ;
assign n24655 =  ( n24654 ) & (wr )  ;
assign n24656 =  ( n24655 ) ? ( n5123 ) : ( iram_203 ) ;
assign n24657 = wr_addr[7:7] ;
assign n24658 =  ( n24657 ) == ( bv_1_0_n53 )  ;
assign n24659 =  ( wr_addr ) == ( bv_8_203_n475 )  ;
assign n24660 =  ( n24658 ) & (n24659 )  ;
assign n24661 =  ( n24660 ) & (wr )  ;
assign n24662 =  ( n24661 ) ? ( n5165 ) : ( iram_203 ) ;
assign n24663 = wr_addr[7:7] ;
assign n24664 =  ( n24663 ) == ( bv_1_0_n53 )  ;
assign n24665 =  ( wr_addr ) == ( bv_8_203_n475 )  ;
assign n24666 =  ( n24664 ) & (n24665 )  ;
assign n24667 =  ( n24666 ) & (wr )  ;
assign n24668 =  ( n24667 ) ? ( n5204 ) : ( iram_203 ) ;
assign n24669 = wr_addr[7:7] ;
assign n24670 =  ( n24669 ) == ( bv_1_0_n53 )  ;
assign n24671 =  ( wr_addr ) == ( bv_8_203_n475 )  ;
assign n24672 =  ( n24670 ) & (n24671 )  ;
assign n24673 =  ( n24672 ) & (wr )  ;
assign n24674 =  ( n24673 ) ? ( n5262 ) : ( iram_203 ) ;
assign n24675 = wr_addr[7:7] ;
assign n24676 =  ( n24675 ) == ( bv_1_0_n53 )  ;
assign n24677 =  ( wr_addr ) == ( bv_8_203_n475 )  ;
assign n24678 =  ( n24676 ) & (n24677 )  ;
assign n24679 =  ( n24678 ) & (wr )  ;
assign n24680 =  ( n24679 ) ? ( n5298 ) : ( iram_203 ) ;
assign n24681 = wr_addr[7:7] ;
assign n24682 =  ( n24681 ) == ( bv_1_0_n53 )  ;
assign n24683 =  ( wr_addr ) == ( bv_8_203_n475 )  ;
assign n24684 =  ( n24682 ) & (n24683 )  ;
assign n24685 =  ( n24684 ) & (wr )  ;
assign n24686 =  ( n24685 ) ? ( n5325 ) : ( iram_203 ) ;
assign n24687 = wr_addr[7:7] ;
assign n24688 =  ( n24687 ) == ( bv_1_0_n53 )  ;
assign n24689 =  ( wr_addr ) == ( bv_8_204_n477 )  ;
assign n24690 =  ( n24688 ) & (n24689 )  ;
assign n24691 =  ( n24690 ) & (wr )  ;
assign n24692 =  ( n24691 ) ? ( n4782 ) : ( iram_204 ) ;
assign n24693 = wr_addr[7:7] ;
assign n24694 =  ( n24693 ) == ( bv_1_0_n53 )  ;
assign n24695 =  ( wr_addr ) == ( bv_8_204_n477 )  ;
assign n24696 =  ( n24694 ) & (n24695 )  ;
assign n24697 =  ( n24696 ) & (wr )  ;
assign n24698 =  ( n24697 ) ? ( n4841 ) : ( iram_204 ) ;
assign n24699 = wr_addr[7:7] ;
assign n24700 =  ( n24699 ) == ( bv_1_0_n53 )  ;
assign n24701 =  ( wr_addr ) == ( bv_8_204_n477 )  ;
assign n24702 =  ( n24700 ) & (n24701 )  ;
assign n24703 =  ( n24702 ) & (wr )  ;
assign n24704 =  ( n24703 ) ? ( n5449 ) : ( iram_204 ) ;
assign n24705 = wr_addr[7:7] ;
assign n24706 =  ( n24705 ) == ( bv_1_0_n53 )  ;
assign n24707 =  ( wr_addr ) == ( bv_8_204_n477 )  ;
assign n24708 =  ( n24706 ) & (n24707 )  ;
assign n24709 =  ( n24708 ) & (wr )  ;
assign n24710 =  ( n24709 ) ? ( n4906 ) : ( iram_204 ) ;
assign n24711 = wr_addr[7:7] ;
assign n24712 =  ( n24711 ) == ( bv_1_0_n53 )  ;
assign n24713 =  ( wr_addr ) == ( bv_8_204_n477 )  ;
assign n24714 =  ( n24712 ) & (n24713 )  ;
assign n24715 =  ( n24714 ) & (wr )  ;
assign n24716 =  ( n24715 ) ? ( n5485 ) : ( iram_204 ) ;
assign n24717 = wr_addr[7:7] ;
assign n24718 =  ( n24717 ) == ( bv_1_0_n53 )  ;
assign n24719 =  ( wr_addr ) == ( bv_8_204_n477 )  ;
assign n24720 =  ( n24718 ) & (n24719 )  ;
assign n24721 =  ( n24720 ) & (wr )  ;
assign n24722 =  ( n24721 ) ? ( n5512 ) : ( iram_204 ) ;
assign n24723 = wr_addr[7:7] ;
assign n24724 =  ( n24723 ) == ( bv_1_0_n53 )  ;
assign n24725 =  ( wr_addr ) == ( bv_8_204_n477 )  ;
assign n24726 =  ( n24724 ) & (n24725 )  ;
assign n24727 =  ( n24726 ) & (wr )  ;
assign n24728 =  ( n24727 ) ? ( bv_8_0_n69 ) : ( iram_204 ) ;
assign n24729 = wr_addr[7:7] ;
assign n24730 =  ( n24729 ) == ( bv_1_0_n53 )  ;
assign n24731 =  ( wr_addr ) == ( bv_8_204_n477 )  ;
assign n24732 =  ( n24730 ) & (n24731 )  ;
assign n24733 =  ( n24732 ) & (wr )  ;
assign n24734 =  ( n24733 ) ? ( n5071 ) : ( iram_204 ) ;
assign n24735 = wr_addr[7:7] ;
assign n24736 =  ( n24735 ) == ( bv_1_0_n53 )  ;
assign n24737 =  ( wr_addr ) == ( bv_8_204_n477 )  ;
assign n24738 =  ( n24736 ) & (n24737 )  ;
assign n24739 =  ( n24738 ) & (wr )  ;
assign n24740 =  ( n24739 ) ? ( n5096 ) : ( iram_204 ) ;
assign n24741 = wr_addr[7:7] ;
assign n24742 =  ( n24741 ) == ( bv_1_0_n53 )  ;
assign n24743 =  ( wr_addr ) == ( bv_8_204_n477 )  ;
assign n24744 =  ( n24742 ) & (n24743 )  ;
assign n24745 =  ( n24744 ) & (wr )  ;
assign n24746 =  ( n24745 ) ? ( n5123 ) : ( iram_204 ) ;
assign n24747 = wr_addr[7:7] ;
assign n24748 =  ( n24747 ) == ( bv_1_0_n53 )  ;
assign n24749 =  ( wr_addr ) == ( bv_8_204_n477 )  ;
assign n24750 =  ( n24748 ) & (n24749 )  ;
assign n24751 =  ( n24750 ) & (wr )  ;
assign n24752 =  ( n24751 ) ? ( n5165 ) : ( iram_204 ) ;
assign n24753 = wr_addr[7:7] ;
assign n24754 =  ( n24753 ) == ( bv_1_0_n53 )  ;
assign n24755 =  ( wr_addr ) == ( bv_8_204_n477 )  ;
assign n24756 =  ( n24754 ) & (n24755 )  ;
assign n24757 =  ( n24756 ) & (wr )  ;
assign n24758 =  ( n24757 ) ? ( n5204 ) : ( iram_204 ) ;
assign n24759 = wr_addr[7:7] ;
assign n24760 =  ( n24759 ) == ( bv_1_0_n53 )  ;
assign n24761 =  ( wr_addr ) == ( bv_8_204_n477 )  ;
assign n24762 =  ( n24760 ) & (n24761 )  ;
assign n24763 =  ( n24762 ) & (wr )  ;
assign n24764 =  ( n24763 ) ? ( n5262 ) : ( iram_204 ) ;
assign n24765 = wr_addr[7:7] ;
assign n24766 =  ( n24765 ) == ( bv_1_0_n53 )  ;
assign n24767 =  ( wr_addr ) == ( bv_8_204_n477 )  ;
assign n24768 =  ( n24766 ) & (n24767 )  ;
assign n24769 =  ( n24768 ) & (wr )  ;
assign n24770 =  ( n24769 ) ? ( n5298 ) : ( iram_204 ) ;
assign n24771 = wr_addr[7:7] ;
assign n24772 =  ( n24771 ) == ( bv_1_0_n53 )  ;
assign n24773 =  ( wr_addr ) == ( bv_8_204_n477 )  ;
assign n24774 =  ( n24772 ) & (n24773 )  ;
assign n24775 =  ( n24774 ) & (wr )  ;
assign n24776 =  ( n24775 ) ? ( n5325 ) : ( iram_204 ) ;
assign n24777 = wr_addr[7:7] ;
assign n24778 =  ( n24777 ) == ( bv_1_0_n53 )  ;
assign n24779 =  ( wr_addr ) == ( bv_8_205_n479 )  ;
assign n24780 =  ( n24778 ) & (n24779 )  ;
assign n24781 =  ( n24780 ) & (wr )  ;
assign n24782 =  ( n24781 ) ? ( n4782 ) : ( iram_205 ) ;
assign n24783 = wr_addr[7:7] ;
assign n24784 =  ( n24783 ) == ( bv_1_0_n53 )  ;
assign n24785 =  ( wr_addr ) == ( bv_8_205_n479 )  ;
assign n24786 =  ( n24784 ) & (n24785 )  ;
assign n24787 =  ( n24786 ) & (wr )  ;
assign n24788 =  ( n24787 ) ? ( n4841 ) : ( iram_205 ) ;
assign n24789 = wr_addr[7:7] ;
assign n24790 =  ( n24789 ) == ( bv_1_0_n53 )  ;
assign n24791 =  ( wr_addr ) == ( bv_8_205_n479 )  ;
assign n24792 =  ( n24790 ) & (n24791 )  ;
assign n24793 =  ( n24792 ) & (wr )  ;
assign n24794 =  ( n24793 ) ? ( n5449 ) : ( iram_205 ) ;
assign n24795 = wr_addr[7:7] ;
assign n24796 =  ( n24795 ) == ( bv_1_0_n53 )  ;
assign n24797 =  ( wr_addr ) == ( bv_8_205_n479 )  ;
assign n24798 =  ( n24796 ) & (n24797 )  ;
assign n24799 =  ( n24798 ) & (wr )  ;
assign n24800 =  ( n24799 ) ? ( n4906 ) : ( iram_205 ) ;
assign n24801 = wr_addr[7:7] ;
assign n24802 =  ( n24801 ) == ( bv_1_0_n53 )  ;
assign n24803 =  ( wr_addr ) == ( bv_8_205_n479 )  ;
assign n24804 =  ( n24802 ) & (n24803 )  ;
assign n24805 =  ( n24804 ) & (wr )  ;
assign n24806 =  ( n24805 ) ? ( n5485 ) : ( iram_205 ) ;
assign n24807 = wr_addr[7:7] ;
assign n24808 =  ( n24807 ) == ( bv_1_0_n53 )  ;
assign n24809 =  ( wr_addr ) == ( bv_8_205_n479 )  ;
assign n24810 =  ( n24808 ) & (n24809 )  ;
assign n24811 =  ( n24810 ) & (wr )  ;
assign n24812 =  ( n24811 ) ? ( n5512 ) : ( iram_205 ) ;
assign n24813 = wr_addr[7:7] ;
assign n24814 =  ( n24813 ) == ( bv_1_0_n53 )  ;
assign n24815 =  ( wr_addr ) == ( bv_8_205_n479 )  ;
assign n24816 =  ( n24814 ) & (n24815 )  ;
assign n24817 =  ( n24816 ) & (wr )  ;
assign n24818 =  ( n24817 ) ? ( bv_8_0_n69 ) : ( iram_205 ) ;
assign n24819 = wr_addr[7:7] ;
assign n24820 =  ( n24819 ) == ( bv_1_0_n53 )  ;
assign n24821 =  ( wr_addr ) == ( bv_8_205_n479 )  ;
assign n24822 =  ( n24820 ) & (n24821 )  ;
assign n24823 =  ( n24822 ) & (wr )  ;
assign n24824 =  ( n24823 ) ? ( n5071 ) : ( iram_205 ) ;
assign n24825 = wr_addr[7:7] ;
assign n24826 =  ( n24825 ) == ( bv_1_0_n53 )  ;
assign n24827 =  ( wr_addr ) == ( bv_8_205_n479 )  ;
assign n24828 =  ( n24826 ) & (n24827 )  ;
assign n24829 =  ( n24828 ) & (wr )  ;
assign n24830 =  ( n24829 ) ? ( n5096 ) : ( iram_205 ) ;
assign n24831 = wr_addr[7:7] ;
assign n24832 =  ( n24831 ) == ( bv_1_0_n53 )  ;
assign n24833 =  ( wr_addr ) == ( bv_8_205_n479 )  ;
assign n24834 =  ( n24832 ) & (n24833 )  ;
assign n24835 =  ( n24834 ) & (wr )  ;
assign n24836 =  ( n24835 ) ? ( n5123 ) : ( iram_205 ) ;
assign n24837 = wr_addr[7:7] ;
assign n24838 =  ( n24837 ) == ( bv_1_0_n53 )  ;
assign n24839 =  ( wr_addr ) == ( bv_8_205_n479 )  ;
assign n24840 =  ( n24838 ) & (n24839 )  ;
assign n24841 =  ( n24840 ) & (wr )  ;
assign n24842 =  ( n24841 ) ? ( n5165 ) : ( iram_205 ) ;
assign n24843 = wr_addr[7:7] ;
assign n24844 =  ( n24843 ) == ( bv_1_0_n53 )  ;
assign n24845 =  ( wr_addr ) == ( bv_8_205_n479 )  ;
assign n24846 =  ( n24844 ) & (n24845 )  ;
assign n24847 =  ( n24846 ) & (wr )  ;
assign n24848 =  ( n24847 ) ? ( n5204 ) : ( iram_205 ) ;
assign n24849 = wr_addr[7:7] ;
assign n24850 =  ( n24849 ) == ( bv_1_0_n53 )  ;
assign n24851 =  ( wr_addr ) == ( bv_8_205_n479 )  ;
assign n24852 =  ( n24850 ) & (n24851 )  ;
assign n24853 =  ( n24852 ) & (wr )  ;
assign n24854 =  ( n24853 ) ? ( n5262 ) : ( iram_205 ) ;
assign n24855 = wr_addr[7:7] ;
assign n24856 =  ( n24855 ) == ( bv_1_0_n53 )  ;
assign n24857 =  ( wr_addr ) == ( bv_8_205_n479 )  ;
assign n24858 =  ( n24856 ) & (n24857 )  ;
assign n24859 =  ( n24858 ) & (wr )  ;
assign n24860 =  ( n24859 ) ? ( n5298 ) : ( iram_205 ) ;
assign n24861 = wr_addr[7:7] ;
assign n24862 =  ( n24861 ) == ( bv_1_0_n53 )  ;
assign n24863 =  ( wr_addr ) == ( bv_8_205_n479 )  ;
assign n24864 =  ( n24862 ) & (n24863 )  ;
assign n24865 =  ( n24864 ) & (wr )  ;
assign n24866 =  ( n24865 ) ? ( n5325 ) : ( iram_205 ) ;
assign n24867 = wr_addr[7:7] ;
assign n24868 =  ( n24867 ) == ( bv_1_0_n53 )  ;
assign n24869 =  ( wr_addr ) == ( bv_8_206_n481 )  ;
assign n24870 =  ( n24868 ) & (n24869 )  ;
assign n24871 =  ( n24870 ) & (wr )  ;
assign n24872 =  ( n24871 ) ? ( n4782 ) : ( iram_206 ) ;
assign n24873 = wr_addr[7:7] ;
assign n24874 =  ( n24873 ) == ( bv_1_0_n53 )  ;
assign n24875 =  ( wr_addr ) == ( bv_8_206_n481 )  ;
assign n24876 =  ( n24874 ) & (n24875 )  ;
assign n24877 =  ( n24876 ) & (wr )  ;
assign n24878 =  ( n24877 ) ? ( n4841 ) : ( iram_206 ) ;
assign n24879 = wr_addr[7:7] ;
assign n24880 =  ( n24879 ) == ( bv_1_0_n53 )  ;
assign n24881 =  ( wr_addr ) == ( bv_8_206_n481 )  ;
assign n24882 =  ( n24880 ) & (n24881 )  ;
assign n24883 =  ( n24882 ) & (wr )  ;
assign n24884 =  ( n24883 ) ? ( n5449 ) : ( iram_206 ) ;
assign n24885 = wr_addr[7:7] ;
assign n24886 =  ( n24885 ) == ( bv_1_0_n53 )  ;
assign n24887 =  ( wr_addr ) == ( bv_8_206_n481 )  ;
assign n24888 =  ( n24886 ) & (n24887 )  ;
assign n24889 =  ( n24888 ) & (wr )  ;
assign n24890 =  ( n24889 ) ? ( n4906 ) : ( iram_206 ) ;
assign n24891 = wr_addr[7:7] ;
assign n24892 =  ( n24891 ) == ( bv_1_0_n53 )  ;
assign n24893 =  ( wr_addr ) == ( bv_8_206_n481 )  ;
assign n24894 =  ( n24892 ) & (n24893 )  ;
assign n24895 =  ( n24894 ) & (wr )  ;
assign n24896 =  ( n24895 ) ? ( n5485 ) : ( iram_206 ) ;
assign n24897 = wr_addr[7:7] ;
assign n24898 =  ( n24897 ) == ( bv_1_0_n53 )  ;
assign n24899 =  ( wr_addr ) == ( bv_8_206_n481 )  ;
assign n24900 =  ( n24898 ) & (n24899 )  ;
assign n24901 =  ( n24900 ) & (wr )  ;
assign n24902 =  ( n24901 ) ? ( n5512 ) : ( iram_206 ) ;
assign n24903 = wr_addr[7:7] ;
assign n24904 =  ( n24903 ) == ( bv_1_0_n53 )  ;
assign n24905 =  ( wr_addr ) == ( bv_8_206_n481 )  ;
assign n24906 =  ( n24904 ) & (n24905 )  ;
assign n24907 =  ( n24906 ) & (wr )  ;
assign n24908 =  ( n24907 ) ? ( bv_8_0_n69 ) : ( iram_206 ) ;
assign n24909 = wr_addr[7:7] ;
assign n24910 =  ( n24909 ) == ( bv_1_0_n53 )  ;
assign n24911 =  ( wr_addr ) == ( bv_8_206_n481 )  ;
assign n24912 =  ( n24910 ) & (n24911 )  ;
assign n24913 =  ( n24912 ) & (wr )  ;
assign n24914 =  ( n24913 ) ? ( n5071 ) : ( iram_206 ) ;
assign n24915 = wr_addr[7:7] ;
assign n24916 =  ( n24915 ) == ( bv_1_0_n53 )  ;
assign n24917 =  ( wr_addr ) == ( bv_8_206_n481 )  ;
assign n24918 =  ( n24916 ) & (n24917 )  ;
assign n24919 =  ( n24918 ) & (wr )  ;
assign n24920 =  ( n24919 ) ? ( n5096 ) : ( iram_206 ) ;
assign n24921 = wr_addr[7:7] ;
assign n24922 =  ( n24921 ) == ( bv_1_0_n53 )  ;
assign n24923 =  ( wr_addr ) == ( bv_8_206_n481 )  ;
assign n24924 =  ( n24922 ) & (n24923 )  ;
assign n24925 =  ( n24924 ) & (wr )  ;
assign n24926 =  ( n24925 ) ? ( n5123 ) : ( iram_206 ) ;
assign n24927 = wr_addr[7:7] ;
assign n24928 =  ( n24927 ) == ( bv_1_0_n53 )  ;
assign n24929 =  ( wr_addr ) == ( bv_8_206_n481 )  ;
assign n24930 =  ( n24928 ) & (n24929 )  ;
assign n24931 =  ( n24930 ) & (wr )  ;
assign n24932 =  ( n24931 ) ? ( n5165 ) : ( iram_206 ) ;
assign n24933 = wr_addr[7:7] ;
assign n24934 =  ( n24933 ) == ( bv_1_0_n53 )  ;
assign n24935 =  ( wr_addr ) == ( bv_8_206_n481 )  ;
assign n24936 =  ( n24934 ) & (n24935 )  ;
assign n24937 =  ( n24936 ) & (wr )  ;
assign n24938 =  ( n24937 ) ? ( n5204 ) : ( iram_206 ) ;
assign n24939 = wr_addr[7:7] ;
assign n24940 =  ( n24939 ) == ( bv_1_0_n53 )  ;
assign n24941 =  ( wr_addr ) == ( bv_8_206_n481 )  ;
assign n24942 =  ( n24940 ) & (n24941 )  ;
assign n24943 =  ( n24942 ) & (wr )  ;
assign n24944 =  ( n24943 ) ? ( n5262 ) : ( iram_206 ) ;
assign n24945 = wr_addr[7:7] ;
assign n24946 =  ( n24945 ) == ( bv_1_0_n53 )  ;
assign n24947 =  ( wr_addr ) == ( bv_8_206_n481 )  ;
assign n24948 =  ( n24946 ) & (n24947 )  ;
assign n24949 =  ( n24948 ) & (wr )  ;
assign n24950 =  ( n24949 ) ? ( n5298 ) : ( iram_206 ) ;
assign n24951 = wr_addr[7:7] ;
assign n24952 =  ( n24951 ) == ( bv_1_0_n53 )  ;
assign n24953 =  ( wr_addr ) == ( bv_8_206_n481 )  ;
assign n24954 =  ( n24952 ) & (n24953 )  ;
assign n24955 =  ( n24954 ) & (wr )  ;
assign n24956 =  ( n24955 ) ? ( n5325 ) : ( iram_206 ) ;
assign n24957 = wr_addr[7:7] ;
assign n24958 =  ( n24957 ) == ( bv_1_0_n53 )  ;
assign n24959 =  ( wr_addr ) == ( bv_8_207_n483 )  ;
assign n24960 =  ( n24958 ) & (n24959 )  ;
assign n24961 =  ( n24960 ) & (wr )  ;
assign n24962 =  ( n24961 ) ? ( n4782 ) : ( iram_207 ) ;
assign n24963 = wr_addr[7:7] ;
assign n24964 =  ( n24963 ) == ( bv_1_0_n53 )  ;
assign n24965 =  ( wr_addr ) == ( bv_8_207_n483 )  ;
assign n24966 =  ( n24964 ) & (n24965 )  ;
assign n24967 =  ( n24966 ) & (wr )  ;
assign n24968 =  ( n24967 ) ? ( n4841 ) : ( iram_207 ) ;
assign n24969 = wr_addr[7:7] ;
assign n24970 =  ( n24969 ) == ( bv_1_0_n53 )  ;
assign n24971 =  ( wr_addr ) == ( bv_8_207_n483 )  ;
assign n24972 =  ( n24970 ) & (n24971 )  ;
assign n24973 =  ( n24972 ) & (wr )  ;
assign n24974 =  ( n24973 ) ? ( n5449 ) : ( iram_207 ) ;
assign n24975 = wr_addr[7:7] ;
assign n24976 =  ( n24975 ) == ( bv_1_0_n53 )  ;
assign n24977 =  ( wr_addr ) == ( bv_8_207_n483 )  ;
assign n24978 =  ( n24976 ) & (n24977 )  ;
assign n24979 =  ( n24978 ) & (wr )  ;
assign n24980 =  ( n24979 ) ? ( n4906 ) : ( iram_207 ) ;
assign n24981 = wr_addr[7:7] ;
assign n24982 =  ( n24981 ) == ( bv_1_0_n53 )  ;
assign n24983 =  ( wr_addr ) == ( bv_8_207_n483 )  ;
assign n24984 =  ( n24982 ) & (n24983 )  ;
assign n24985 =  ( n24984 ) & (wr )  ;
assign n24986 =  ( n24985 ) ? ( n5485 ) : ( iram_207 ) ;
assign n24987 = wr_addr[7:7] ;
assign n24988 =  ( n24987 ) == ( bv_1_0_n53 )  ;
assign n24989 =  ( wr_addr ) == ( bv_8_207_n483 )  ;
assign n24990 =  ( n24988 ) & (n24989 )  ;
assign n24991 =  ( n24990 ) & (wr )  ;
assign n24992 =  ( n24991 ) ? ( n5512 ) : ( iram_207 ) ;
assign n24993 = wr_addr[7:7] ;
assign n24994 =  ( n24993 ) == ( bv_1_0_n53 )  ;
assign n24995 =  ( wr_addr ) == ( bv_8_207_n483 )  ;
assign n24996 =  ( n24994 ) & (n24995 )  ;
assign n24997 =  ( n24996 ) & (wr )  ;
assign n24998 =  ( n24997 ) ? ( bv_8_0_n69 ) : ( iram_207 ) ;
assign n24999 = wr_addr[7:7] ;
assign n25000 =  ( n24999 ) == ( bv_1_0_n53 )  ;
assign n25001 =  ( wr_addr ) == ( bv_8_207_n483 )  ;
assign n25002 =  ( n25000 ) & (n25001 )  ;
assign n25003 =  ( n25002 ) & (wr )  ;
assign n25004 =  ( n25003 ) ? ( n5071 ) : ( iram_207 ) ;
assign n25005 = wr_addr[7:7] ;
assign n25006 =  ( n25005 ) == ( bv_1_0_n53 )  ;
assign n25007 =  ( wr_addr ) == ( bv_8_207_n483 )  ;
assign n25008 =  ( n25006 ) & (n25007 )  ;
assign n25009 =  ( n25008 ) & (wr )  ;
assign n25010 =  ( n25009 ) ? ( n5096 ) : ( iram_207 ) ;
assign n25011 = wr_addr[7:7] ;
assign n25012 =  ( n25011 ) == ( bv_1_0_n53 )  ;
assign n25013 =  ( wr_addr ) == ( bv_8_207_n483 )  ;
assign n25014 =  ( n25012 ) & (n25013 )  ;
assign n25015 =  ( n25014 ) & (wr )  ;
assign n25016 =  ( n25015 ) ? ( n5123 ) : ( iram_207 ) ;
assign n25017 = wr_addr[7:7] ;
assign n25018 =  ( n25017 ) == ( bv_1_0_n53 )  ;
assign n25019 =  ( wr_addr ) == ( bv_8_207_n483 )  ;
assign n25020 =  ( n25018 ) & (n25019 )  ;
assign n25021 =  ( n25020 ) & (wr )  ;
assign n25022 =  ( n25021 ) ? ( n5165 ) : ( iram_207 ) ;
assign n25023 = wr_addr[7:7] ;
assign n25024 =  ( n25023 ) == ( bv_1_0_n53 )  ;
assign n25025 =  ( wr_addr ) == ( bv_8_207_n483 )  ;
assign n25026 =  ( n25024 ) & (n25025 )  ;
assign n25027 =  ( n25026 ) & (wr )  ;
assign n25028 =  ( n25027 ) ? ( n5204 ) : ( iram_207 ) ;
assign n25029 = wr_addr[7:7] ;
assign n25030 =  ( n25029 ) == ( bv_1_0_n53 )  ;
assign n25031 =  ( wr_addr ) == ( bv_8_207_n483 )  ;
assign n25032 =  ( n25030 ) & (n25031 )  ;
assign n25033 =  ( n25032 ) & (wr )  ;
assign n25034 =  ( n25033 ) ? ( n5262 ) : ( iram_207 ) ;
assign n25035 = wr_addr[7:7] ;
assign n25036 =  ( n25035 ) == ( bv_1_0_n53 )  ;
assign n25037 =  ( wr_addr ) == ( bv_8_207_n483 )  ;
assign n25038 =  ( n25036 ) & (n25037 )  ;
assign n25039 =  ( n25038 ) & (wr )  ;
assign n25040 =  ( n25039 ) ? ( n5298 ) : ( iram_207 ) ;
assign n25041 = wr_addr[7:7] ;
assign n25042 =  ( n25041 ) == ( bv_1_0_n53 )  ;
assign n25043 =  ( wr_addr ) == ( bv_8_207_n483 )  ;
assign n25044 =  ( n25042 ) & (n25043 )  ;
assign n25045 =  ( n25044 ) & (wr )  ;
assign n25046 =  ( n25045 ) ? ( n5325 ) : ( iram_207 ) ;
assign n25047 = wr_addr[7:7] ;
assign n25048 =  ( n25047 ) == ( bv_1_0_n53 )  ;
assign n25049 =  ( wr_addr ) == ( bv_8_208_n485 )  ;
assign n25050 =  ( n25048 ) & (n25049 )  ;
assign n25051 =  ( n25050 ) & (wr )  ;
assign n25052 =  ( n25051 ) ? ( n4782 ) : ( iram_208 ) ;
assign n25053 = wr_addr[7:7] ;
assign n25054 =  ( n25053 ) == ( bv_1_0_n53 )  ;
assign n25055 =  ( wr_addr ) == ( bv_8_208_n485 )  ;
assign n25056 =  ( n25054 ) & (n25055 )  ;
assign n25057 =  ( n25056 ) & (wr )  ;
assign n25058 =  ( n25057 ) ? ( n4841 ) : ( iram_208 ) ;
assign n25059 = wr_addr[7:7] ;
assign n25060 =  ( n25059 ) == ( bv_1_0_n53 )  ;
assign n25061 =  ( wr_addr ) == ( bv_8_208_n485 )  ;
assign n25062 =  ( n25060 ) & (n25061 )  ;
assign n25063 =  ( n25062 ) & (wr )  ;
assign n25064 =  ( n25063 ) ? ( n5449 ) : ( iram_208 ) ;
assign n25065 = wr_addr[7:7] ;
assign n25066 =  ( n25065 ) == ( bv_1_0_n53 )  ;
assign n25067 =  ( wr_addr ) == ( bv_8_208_n485 )  ;
assign n25068 =  ( n25066 ) & (n25067 )  ;
assign n25069 =  ( n25068 ) & (wr )  ;
assign n25070 =  ( n25069 ) ? ( n4906 ) : ( iram_208 ) ;
assign n25071 = wr_addr[7:7] ;
assign n25072 =  ( n25071 ) == ( bv_1_0_n53 )  ;
assign n25073 =  ( wr_addr ) == ( bv_8_208_n485 )  ;
assign n25074 =  ( n25072 ) & (n25073 )  ;
assign n25075 =  ( n25074 ) & (wr )  ;
assign n25076 =  ( n25075 ) ? ( n5485 ) : ( iram_208 ) ;
assign n25077 = wr_addr[7:7] ;
assign n25078 =  ( n25077 ) == ( bv_1_0_n53 )  ;
assign n25079 =  ( wr_addr ) == ( bv_8_208_n485 )  ;
assign n25080 =  ( n25078 ) & (n25079 )  ;
assign n25081 =  ( n25080 ) & (wr )  ;
assign n25082 =  ( n25081 ) ? ( n5512 ) : ( iram_208 ) ;
assign n25083 = wr_addr[7:7] ;
assign n25084 =  ( n25083 ) == ( bv_1_0_n53 )  ;
assign n25085 =  ( wr_addr ) == ( bv_8_208_n485 )  ;
assign n25086 =  ( n25084 ) & (n25085 )  ;
assign n25087 =  ( n25086 ) & (wr )  ;
assign n25088 =  ( n25087 ) ? ( bv_8_0_n69 ) : ( iram_208 ) ;
assign n25089 = wr_addr[7:7] ;
assign n25090 =  ( n25089 ) == ( bv_1_0_n53 )  ;
assign n25091 =  ( wr_addr ) == ( bv_8_208_n485 )  ;
assign n25092 =  ( n25090 ) & (n25091 )  ;
assign n25093 =  ( n25092 ) & (wr )  ;
assign n25094 =  ( n25093 ) ? ( n5071 ) : ( iram_208 ) ;
assign n25095 = wr_addr[7:7] ;
assign n25096 =  ( n25095 ) == ( bv_1_0_n53 )  ;
assign n25097 =  ( wr_addr ) == ( bv_8_208_n485 )  ;
assign n25098 =  ( n25096 ) & (n25097 )  ;
assign n25099 =  ( n25098 ) & (wr )  ;
assign n25100 =  ( n25099 ) ? ( n5096 ) : ( iram_208 ) ;
assign n25101 = wr_addr[7:7] ;
assign n25102 =  ( n25101 ) == ( bv_1_0_n53 )  ;
assign n25103 =  ( wr_addr ) == ( bv_8_208_n485 )  ;
assign n25104 =  ( n25102 ) & (n25103 )  ;
assign n25105 =  ( n25104 ) & (wr )  ;
assign n25106 =  ( n25105 ) ? ( n5123 ) : ( iram_208 ) ;
assign n25107 = wr_addr[7:7] ;
assign n25108 =  ( n25107 ) == ( bv_1_0_n53 )  ;
assign n25109 =  ( wr_addr ) == ( bv_8_208_n485 )  ;
assign n25110 =  ( n25108 ) & (n25109 )  ;
assign n25111 =  ( n25110 ) & (wr )  ;
assign n25112 =  ( n25111 ) ? ( n5165 ) : ( iram_208 ) ;
assign n25113 = wr_addr[7:7] ;
assign n25114 =  ( n25113 ) == ( bv_1_0_n53 )  ;
assign n25115 =  ( wr_addr ) == ( bv_8_208_n485 )  ;
assign n25116 =  ( n25114 ) & (n25115 )  ;
assign n25117 =  ( n25116 ) & (wr )  ;
assign n25118 =  ( n25117 ) ? ( n5204 ) : ( iram_208 ) ;
assign n25119 = wr_addr[7:7] ;
assign n25120 =  ( n25119 ) == ( bv_1_0_n53 )  ;
assign n25121 =  ( wr_addr ) == ( bv_8_208_n485 )  ;
assign n25122 =  ( n25120 ) & (n25121 )  ;
assign n25123 =  ( n25122 ) & (wr )  ;
assign n25124 =  ( n25123 ) ? ( n5262 ) : ( iram_208 ) ;
assign n25125 = wr_addr[7:7] ;
assign n25126 =  ( n25125 ) == ( bv_1_0_n53 )  ;
assign n25127 =  ( wr_addr ) == ( bv_8_208_n485 )  ;
assign n25128 =  ( n25126 ) & (n25127 )  ;
assign n25129 =  ( n25128 ) & (wr )  ;
assign n25130 =  ( n25129 ) ? ( n5298 ) : ( iram_208 ) ;
assign n25131 = wr_addr[7:7] ;
assign n25132 =  ( n25131 ) == ( bv_1_0_n53 )  ;
assign n25133 =  ( wr_addr ) == ( bv_8_208_n485 )  ;
assign n25134 =  ( n25132 ) & (n25133 )  ;
assign n25135 =  ( n25134 ) & (wr )  ;
assign n25136 =  ( n25135 ) ? ( n5325 ) : ( iram_208 ) ;
assign n25137 = wr_addr[7:7] ;
assign n25138 =  ( n25137 ) == ( bv_1_0_n53 )  ;
assign n25139 =  ( wr_addr ) == ( bv_8_209_n487 )  ;
assign n25140 =  ( n25138 ) & (n25139 )  ;
assign n25141 =  ( n25140 ) & (wr )  ;
assign n25142 =  ( n25141 ) ? ( n4782 ) : ( iram_209 ) ;
assign n25143 = wr_addr[7:7] ;
assign n25144 =  ( n25143 ) == ( bv_1_0_n53 )  ;
assign n25145 =  ( wr_addr ) == ( bv_8_209_n487 )  ;
assign n25146 =  ( n25144 ) & (n25145 )  ;
assign n25147 =  ( n25146 ) & (wr )  ;
assign n25148 =  ( n25147 ) ? ( n4841 ) : ( iram_209 ) ;
assign n25149 = wr_addr[7:7] ;
assign n25150 =  ( n25149 ) == ( bv_1_0_n53 )  ;
assign n25151 =  ( wr_addr ) == ( bv_8_209_n487 )  ;
assign n25152 =  ( n25150 ) & (n25151 )  ;
assign n25153 =  ( n25152 ) & (wr )  ;
assign n25154 =  ( n25153 ) ? ( n5449 ) : ( iram_209 ) ;
assign n25155 = wr_addr[7:7] ;
assign n25156 =  ( n25155 ) == ( bv_1_0_n53 )  ;
assign n25157 =  ( wr_addr ) == ( bv_8_209_n487 )  ;
assign n25158 =  ( n25156 ) & (n25157 )  ;
assign n25159 =  ( n25158 ) & (wr )  ;
assign n25160 =  ( n25159 ) ? ( n4906 ) : ( iram_209 ) ;
assign n25161 = wr_addr[7:7] ;
assign n25162 =  ( n25161 ) == ( bv_1_0_n53 )  ;
assign n25163 =  ( wr_addr ) == ( bv_8_209_n487 )  ;
assign n25164 =  ( n25162 ) & (n25163 )  ;
assign n25165 =  ( n25164 ) & (wr )  ;
assign n25166 =  ( n25165 ) ? ( n5485 ) : ( iram_209 ) ;
assign n25167 = wr_addr[7:7] ;
assign n25168 =  ( n25167 ) == ( bv_1_0_n53 )  ;
assign n25169 =  ( wr_addr ) == ( bv_8_209_n487 )  ;
assign n25170 =  ( n25168 ) & (n25169 )  ;
assign n25171 =  ( n25170 ) & (wr )  ;
assign n25172 =  ( n25171 ) ? ( n5512 ) : ( iram_209 ) ;
assign n25173 = wr_addr[7:7] ;
assign n25174 =  ( n25173 ) == ( bv_1_0_n53 )  ;
assign n25175 =  ( wr_addr ) == ( bv_8_209_n487 )  ;
assign n25176 =  ( n25174 ) & (n25175 )  ;
assign n25177 =  ( n25176 ) & (wr )  ;
assign n25178 =  ( n25177 ) ? ( bv_8_0_n69 ) : ( iram_209 ) ;
assign n25179 = wr_addr[7:7] ;
assign n25180 =  ( n25179 ) == ( bv_1_0_n53 )  ;
assign n25181 =  ( wr_addr ) == ( bv_8_209_n487 )  ;
assign n25182 =  ( n25180 ) & (n25181 )  ;
assign n25183 =  ( n25182 ) & (wr )  ;
assign n25184 =  ( n25183 ) ? ( n5071 ) : ( iram_209 ) ;
assign n25185 = wr_addr[7:7] ;
assign n25186 =  ( n25185 ) == ( bv_1_0_n53 )  ;
assign n25187 =  ( wr_addr ) == ( bv_8_209_n487 )  ;
assign n25188 =  ( n25186 ) & (n25187 )  ;
assign n25189 =  ( n25188 ) & (wr )  ;
assign n25190 =  ( n25189 ) ? ( n5096 ) : ( iram_209 ) ;
assign n25191 = wr_addr[7:7] ;
assign n25192 =  ( n25191 ) == ( bv_1_0_n53 )  ;
assign n25193 =  ( wr_addr ) == ( bv_8_209_n487 )  ;
assign n25194 =  ( n25192 ) & (n25193 )  ;
assign n25195 =  ( n25194 ) & (wr )  ;
assign n25196 =  ( n25195 ) ? ( n5123 ) : ( iram_209 ) ;
assign n25197 = wr_addr[7:7] ;
assign n25198 =  ( n25197 ) == ( bv_1_0_n53 )  ;
assign n25199 =  ( wr_addr ) == ( bv_8_209_n487 )  ;
assign n25200 =  ( n25198 ) & (n25199 )  ;
assign n25201 =  ( n25200 ) & (wr )  ;
assign n25202 =  ( n25201 ) ? ( n5165 ) : ( iram_209 ) ;
assign n25203 = wr_addr[7:7] ;
assign n25204 =  ( n25203 ) == ( bv_1_0_n53 )  ;
assign n25205 =  ( wr_addr ) == ( bv_8_209_n487 )  ;
assign n25206 =  ( n25204 ) & (n25205 )  ;
assign n25207 =  ( n25206 ) & (wr )  ;
assign n25208 =  ( n25207 ) ? ( n5204 ) : ( iram_209 ) ;
assign n25209 = wr_addr[7:7] ;
assign n25210 =  ( n25209 ) == ( bv_1_0_n53 )  ;
assign n25211 =  ( wr_addr ) == ( bv_8_209_n487 )  ;
assign n25212 =  ( n25210 ) & (n25211 )  ;
assign n25213 =  ( n25212 ) & (wr )  ;
assign n25214 =  ( n25213 ) ? ( n5262 ) : ( iram_209 ) ;
assign n25215 = wr_addr[7:7] ;
assign n25216 =  ( n25215 ) == ( bv_1_0_n53 )  ;
assign n25217 =  ( wr_addr ) == ( bv_8_209_n487 )  ;
assign n25218 =  ( n25216 ) & (n25217 )  ;
assign n25219 =  ( n25218 ) & (wr )  ;
assign n25220 =  ( n25219 ) ? ( n5298 ) : ( iram_209 ) ;
assign n25221 = wr_addr[7:7] ;
assign n25222 =  ( n25221 ) == ( bv_1_0_n53 )  ;
assign n25223 =  ( wr_addr ) == ( bv_8_209_n487 )  ;
assign n25224 =  ( n25222 ) & (n25223 )  ;
assign n25225 =  ( n25224 ) & (wr )  ;
assign n25226 =  ( n25225 ) ? ( n5325 ) : ( iram_209 ) ;
assign n25227 = wr_addr[7:7] ;
assign n25228 =  ( n25227 ) == ( bv_1_0_n53 )  ;
assign n25229 =  ( wr_addr ) == ( bv_8_210_n489 )  ;
assign n25230 =  ( n25228 ) & (n25229 )  ;
assign n25231 =  ( n25230 ) & (wr )  ;
assign n25232 =  ( n25231 ) ? ( n4782 ) : ( iram_210 ) ;
assign n25233 = wr_addr[7:7] ;
assign n25234 =  ( n25233 ) == ( bv_1_0_n53 )  ;
assign n25235 =  ( wr_addr ) == ( bv_8_210_n489 )  ;
assign n25236 =  ( n25234 ) & (n25235 )  ;
assign n25237 =  ( n25236 ) & (wr )  ;
assign n25238 =  ( n25237 ) ? ( n4841 ) : ( iram_210 ) ;
assign n25239 = wr_addr[7:7] ;
assign n25240 =  ( n25239 ) == ( bv_1_0_n53 )  ;
assign n25241 =  ( wr_addr ) == ( bv_8_210_n489 )  ;
assign n25242 =  ( n25240 ) & (n25241 )  ;
assign n25243 =  ( n25242 ) & (wr )  ;
assign n25244 =  ( n25243 ) ? ( n5449 ) : ( iram_210 ) ;
assign n25245 = wr_addr[7:7] ;
assign n25246 =  ( n25245 ) == ( bv_1_0_n53 )  ;
assign n25247 =  ( wr_addr ) == ( bv_8_210_n489 )  ;
assign n25248 =  ( n25246 ) & (n25247 )  ;
assign n25249 =  ( n25248 ) & (wr )  ;
assign n25250 =  ( n25249 ) ? ( n4906 ) : ( iram_210 ) ;
assign n25251 = wr_addr[7:7] ;
assign n25252 =  ( n25251 ) == ( bv_1_0_n53 )  ;
assign n25253 =  ( wr_addr ) == ( bv_8_210_n489 )  ;
assign n25254 =  ( n25252 ) & (n25253 )  ;
assign n25255 =  ( n25254 ) & (wr )  ;
assign n25256 =  ( n25255 ) ? ( n5485 ) : ( iram_210 ) ;
assign n25257 = wr_addr[7:7] ;
assign n25258 =  ( n25257 ) == ( bv_1_0_n53 )  ;
assign n25259 =  ( wr_addr ) == ( bv_8_210_n489 )  ;
assign n25260 =  ( n25258 ) & (n25259 )  ;
assign n25261 =  ( n25260 ) & (wr )  ;
assign n25262 =  ( n25261 ) ? ( n5512 ) : ( iram_210 ) ;
assign n25263 = wr_addr[7:7] ;
assign n25264 =  ( n25263 ) == ( bv_1_0_n53 )  ;
assign n25265 =  ( wr_addr ) == ( bv_8_210_n489 )  ;
assign n25266 =  ( n25264 ) & (n25265 )  ;
assign n25267 =  ( n25266 ) & (wr )  ;
assign n25268 =  ( n25267 ) ? ( bv_8_0_n69 ) : ( iram_210 ) ;
assign n25269 = wr_addr[7:7] ;
assign n25270 =  ( n25269 ) == ( bv_1_0_n53 )  ;
assign n25271 =  ( wr_addr ) == ( bv_8_210_n489 )  ;
assign n25272 =  ( n25270 ) & (n25271 )  ;
assign n25273 =  ( n25272 ) & (wr )  ;
assign n25274 =  ( n25273 ) ? ( n5071 ) : ( iram_210 ) ;
assign n25275 = wr_addr[7:7] ;
assign n25276 =  ( n25275 ) == ( bv_1_0_n53 )  ;
assign n25277 =  ( wr_addr ) == ( bv_8_210_n489 )  ;
assign n25278 =  ( n25276 ) & (n25277 )  ;
assign n25279 =  ( n25278 ) & (wr )  ;
assign n25280 =  ( n25279 ) ? ( n5096 ) : ( iram_210 ) ;
assign n25281 = wr_addr[7:7] ;
assign n25282 =  ( n25281 ) == ( bv_1_0_n53 )  ;
assign n25283 =  ( wr_addr ) == ( bv_8_210_n489 )  ;
assign n25284 =  ( n25282 ) & (n25283 )  ;
assign n25285 =  ( n25284 ) & (wr )  ;
assign n25286 =  ( n25285 ) ? ( n5123 ) : ( iram_210 ) ;
assign n25287 = wr_addr[7:7] ;
assign n25288 =  ( n25287 ) == ( bv_1_0_n53 )  ;
assign n25289 =  ( wr_addr ) == ( bv_8_210_n489 )  ;
assign n25290 =  ( n25288 ) & (n25289 )  ;
assign n25291 =  ( n25290 ) & (wr )  ;
assign n25292 =  ( n25291 ) ? ( n5165 ) : ( iram_210 ) ;
assign n25293 = wr_addr[7:7] ;
assign n25294 =  ( n25293 ) == ( bv_1_0_n53 )  ;
assign n25295 =  ( wr_addr ) == ( bv_8_210_n489 )  ;
assign n25296 =  ( n25294 ) & (n25295 )  ;
assign n25297 =  ( n25296 ) & (wr )  ;
assign n25298 =  ( n25297 ) ? ( n5204 ) : ( iram_210 ) ;
assign n25299 = wr_addr[7:7] ;
assign n25300 =  ( n25299 ) == ( bv_1_0_n53 )  ;
assign n25301 =  ( wr_addr ) == ( bv_8_210_n489 )  ;
assign n25302 =  ( n25300 ) & (n25301 )  ;
assign n25303 =  ( n25302 ) & (wr )  ;
assign n25304 =  ( n25303 ) ? ( n5262 ) : ( iram_210 ) ;
assign n25305 = wr_addr[7:7] ;
assign n25306 =  ( n25305 ) == ( bv_1_0_n53 )  ;
assign n25307 =  ( wr_addr ) == ( bv_8_210_n489 )  ;
assign n25308 =  ( n25306 ) & (n25307 )  ;
assign n25309 =  ( n25308 ) & (wr )  ;
assign n25310 =  ( n25309 ) ? ( n5298 ) : ( iram_210 ) ;
assign n25311 = wr_addr[7:7] ;
assign n25312 =  ( n25311 ) == ( bv_1_0_n53 )  ;
assign n25313 =  ( wr_addr ) == ( bv_8_210_n489 )  ;
assign n25314 =  ( n25312 ) & (n25313 )  ;
assign n25315 =  ( n25314 ) & (wr )  ;
assign n25316 =  ( n25315 ) ? ( n5325 ) : ( iram_210 ) ;
assign n25317 = wr_addr[7:7] ;
assign n25318 =  ( n25317 ) == ( bv_1_0_n53 )  ;
assign n25319 =  ( wr_addr ) == ( bv_8_211_n491 )  ;
assign n25320 =  ( n25318 ) & (n25319 )  ;
assign n25321 =  ( n25320 ) & (wr )  ;
assign n25322 =  ( n25321 ) ? ( n4782 ) : ( iram_211 ) ;
assign n25323 = wr_addr[7:7] ;
assign n25324 =  ( n25323 ) == ( bv_1_0_n53 )  ;
assign n25325 =  ( wr_addr ) == ( bv_8_211_n491 )  ;
assign n25326 =  ( n25324 ) & (n25325 )  ;
assign n25327 =  ( n25326 ) & (wr )  ;
assign n25328 =  ( n25327 ) ? ( n4841 ) : ( iram_211 ) ;
assign n25329 = wr_addr[7:7] ;
assign n25330 =  ( n25329 ) == ( bv_1_0_n53 )  ;
assign n25331 =  ( wr_addr ) == ( bv_8_211_n491 )  ;
assign n25332 =  ( n25330 ) & (n25331 )  ;
assign n25333 =  ( n25332 ) & (wr )  ;
assign n25334 =  ( n25333 ) ? ( n5449 ) : ( iram_211 ) ;
assign n25335 = wr_addr[7:7] ;
assign n25336 =  ( n25335 ) == ( bv_1_0_n53 )  ;
assign n25337 =  ( wr_addr ) == ( bv_8_211_n491 )  ;
assign n25338 =  ( n25336 ) & (n25337 )  ;
assign n25339 =  ( n25338 ) & (wr )  ;
assign n25340 =  ( n25339 ) ? ( n4906 ) : ( iram_211 ) ;
assign n25341 = wr_addr[7:7] ;
assign n25342 =  ( n25341 ) == ( bv_1_0_n53 )  ;
assign n25343 =  ( wr_addr ) == ( bv_8_211_n491 )  ;
assign n25344 =  ( n25342 ) & (n25343 )  ;
assign n25345 =  ( n25344 ) & (wr )  ;
assign n25346 =  ( n25345 ) ? ( n5485 ) : ( iram_211 ) ;
assign n25347 = wr_addr[7:7] ;
assign n25348 =  ( n25347 ) == ( bv_1_0_n53 )  ;
assign n25349 =  ( wr_addr ) == ( bv_8_211_n491 )  ;
assign n25350 =  ( n25348 ) & (n25349 )  ;
assign n25351 =  ( n25350 ) & (wr )  ;
assign n25352 =  ( n25351 ) ? ( n5512 ) : ( iram_211 ) ;
assign n25353 = wr_addr[7:7] ;
assign n25354 =  ( n25353 ) == ( bv_1_0_n53 )  ;
assign n25355 =  ( wr_addr ) == ( bv_8_211_n491 )  ;
assign n25356 =  ( n25354 ) & (n25355 )  ;
assign n25357 =  ( n25356 ) & (wr )  ;
assign n25358 =  ( n25357 ) ? ( bv_8_0_n69 ) : ( iram_211 ) ;
assign n25359 = wr_addr[7:7] ;
assign n25360 =  ( n25359 ) == ( bv_1_0_n53 )  ;
assign n25361 =  ( wr_addr ) == ( bv_8_211_n491 )  ;
assign n25362 =  ( n25360 ) & (n25361 )  ;
assign n25363 =  ( n25362 ) & (wr )  ;
assign n25364 =  ( n25363 ) ? ( n5071 ) : ( iram_211 ) ;
assign n25365 = wr_addr[7:7] ;
assign n25366 =  ( n25365 ) == ( bv_1_0_n53 )  ;
assign n25367 =  ( wr_addr ) == ( bv_8_211_n491 )  ;
assign n25368 =  ( n25366 ) & (n25367 )  ;
assign n25369 =  ( n25368 ) & (wr )  ;
assign n25370 =  ( n25369 ) ? ( n5096 ) : ( iram_211 ) ;
assign n25371 = wr_addr[7:7] ;
assign n25372 =  ( n25371 ) == ( bv_1_0_n53 )  ;
assign n25373 =  ( wr_addr ) == ( bv_8_211_n491 )  ;
assign n25374 =  ( n25372 ) & (n25373 )  ;
assign n25375 =  ( n25374 ) & (wr )  ;
assign n25376 =  ( n25375 ) ? ( n5123 ) : ( iram_211 ) ;
assign n25377 = wr_addr[7:7] ;
assign n25378 =  ( n25377 ) == ( bv_1_0_n53 )  ;
assign n25379 =  ( wr_addr ) == ( bv_8_211_n491 )  ;
assign n25380 =  ( n25378 ) & (n25379 )  ;
assign n25381 =  ( n25380 ) & (wr )  ;
assign n25382 =  ( n25381 ) ? ( n5165 ) : ( iram_211 ) ;
assign n25383 = wr_addr[7:7] ;
assign n25384 =  ( n25383 ) == ( bv_1_0_n53 )  ;
assign n25385 =  ( wr_addr ) == ( bv_8_211_n491 )  ;
assign n25386 =  ( n25384 ) & (n25385 )  ;
assign n25387 =  ( n25386 ) & (wr )  ;
assign n25388 =  ( n25387 ) ? ( n5204 ) : ( iram_211 ) ;
assign n25389 = wr_addr[7:7] ;
assign n25390 =  ( n25389 ) == ( bv_1_0_n53 )  ;
assign n25391 =  ( wr_addr ) == ( bv_8_211_n491 )  ;
assign n25392 =  ( n25390 ) & (n25391 )  ;
assign n25393 =  ( n25392 ) & (wr )  ;
assign n25394 =  ( n25393 ) ? ( n5262 ) : ( iram_211 ) ;
assign n25395 = wr_addr[7:7] ;
assign n25396 =  ( n25395 ) == ( bv_1_0_n53 )  ;
assign n25397 =  ( wr_addr ) == ( bv_8_211_n491 )  ;
assign n25398 =  ( n25396 ) & (n25397 )  ;
assign n25399 =  ( n25398 ) & (wr )  ;
assign n25400 =  ( n25399 ) ? ( n5298 ) : ( iram_211 ) ;
assign n25401 = wr_addr[7:7] ;
assign n25402 =  ( n25401 ) == ( bv_1_0_n53 )  ;
assign n25403 =  ( wr_addr ) == ( bv_8_211_n491 )  ;
assign n25404 =  ( n25402 ) & (n25403 )  ;
assign n25405 =  ( n25404 ) & (wr )  ;
assign n25406 =  ( n25405 ) ? ( n5325 ) : ( iram_211 ) ;
assign n25407 = wr_addr[7:7] ;
assign n25408 =  ( n25407 ) == ( bv_1_0_n53 )  ;
assign n25409 =  ( wr_addr ) == ( bv_8_212_n493 )  ;
assign n25410 =  ( n25408 ) & (n25409 )  ;
assign n25411 =  ( n25410 ) & (wr )  ;
assign n25412 =  ( n25411 ) ? ( n4782 ) : ( iram_212 ) ;
assign n25413 = wr_addr[7:7] ;
assign n25414 =  ( n25413 ) == ( bv_1_0_n53 )  ;
assign n25415 =  ( wr_addr ) == ( bv_8_212_n493 )  ;
assign n25416 =  ( n25414 ) & (n25415 )  ;
assign n25417 =  ( n25416 ) & (wr )  ;
assign n25418 =  ( n25417 ) ? ( n4841 ) : ( iram_212 ) ;
assign n25419 = wr_addr[7:7] ;
assign n25420 =  ( n25419 ) == ( bv_1_0_n53 )  ;
assign n25421 =  ( wr_addr ) == ( bv_8_212_n493 )  ;
assign n25422 =  ( n25420 ) & (n25421 )  ;
assign n25423 =  ( n25422 ) & (wr )  ;
assign n25424 =  ( n25423 ) ? ( n5449 ) : ( iram_212 ) ;
assign n25425 = wr_addr[7:7] ;
assign n25426 =  ( n25425 ) == ( bv_1_0_n53 )  ;
assign n25427 =  ( wr_addr ) == ( bv_8_212_n493 )  ;
assign n25428 =  ( n25426 ) & (n25427 )  ;
assign n25429 =  ( n25428 ) & (wr )  ;
assign n25430 =  ( n25429 ) ? ( n4906 ) : ( iram_212 ) ;
assign n25431 = wr_addr[7:7] ;
assign n25432 =  ( n25431 ) == ( bv_1_0_n53 )  ;
assign n25433 =  ( wr_addr ) == ( bv_8_212_n493 )  ;
assign n25434 =  ( n25432 ) & (n25433 )  ;
assign n25435 =  ( n25434 ) & (wr )  ;
assign n25436 =  ( n25435 ) ? ( n5485 ) : ( iram_212 ) ;
assign n25437 = wr_addr[7:7] ;
assign n25438 =  ( n25437 ) == ( bv_1_0_n53 )  ;
assign n25439 =  ( wr_addr ) == ( bv_8_212_n493 )  ;
assign n25440 =  ( n25438 ) & (n25439 )  ;
assign n25441 =  ( n25440 ) & (wr )  ;
assign n25442 =  ( n25441 ) ? ( n5512 ) : ( iram_212 ) ;
assign n25443 = wr_addr[7:7] ;
assign n25444 =  ( n25443 ) == ( bv_1_0_n53 )  ;
assign n25445 =  ( wr_addr ) == ( bv_8_212_n493 )  ;
assign n25446 =  ( n25444 ) & (n25445 )  ;
assign n25447 =  ( n25446 ) & (wr )  ;
assign n25448 =  ( n25447 ) ? ( bv_8_0_n69 ) : ( iram_212 ) ;
assign n25449 = wr_addr[7:7] ;
assign n25450 =  ( n25449 ) == ( bv_1_0_n53 )  ;
assign n25451 =  ( wr_addr ) == ( bv_8_212_n493 )  ;
assign n25452 =  ( n25450 ) & (n25451 )  ;
assign n25453 =  ( n25452 ) & (wr )  ;
assign n25454 =  ( n25453 ) ? ( n5071 ) : ( iram_212 ) ;
assign n25455 = wr_addr[7:7] ;
assign n25456 =  ( n25455 ) == ( bv_1_0_n53 )  ;
assign n25457 =  ( wr_addr ) == ( bv_8_212_n493 )  ;
assign n25458 =  ( n25456 ) & (n25457 )  ;
assign n25459 =  ( n25458 ) & (wr )  ;
assign n25460 =  ( n25459 ) ? ( n5096 ) : ( iram_212 ) ;
assign n25461 = wr_addr[7:7] ;
assign n25462 =  ( n25461 ) == ( bv_1_0_n53 )  ;
assign n25463 =  ( wr_addr ) == ( bv_8_212_n493 )  ;
assign n25464 =  ( n25462 ) & (n25463 )  ;
assign n25465 =  ( n25464 ) & (wr )  ;
assign n25466 =  ( n25465 ) ? ( n5123 ) : ( iram_212 ) ;
assign n25467 = wr_addr[7:7] ;
assign n25468 =  ( n25467 ) == ( bv_1_0_n53 )  ;
assign n25469 =  ( wr_addr ) == ( bv_8_212_n493 )  ;
assign n25470 =  ( n25468 ) & (n25469 )  ;
assign n25471 =  ( n25470 ) & (wr )  ;
assign n25472 =  ( n25471 ) ? ( n5165 ) : ( iram_212 ) ;
assign n25473 = wr_addr[7:7] ;
assign n25474 =  ( n25473 ) == ( bv_1_0_n53 )  ;
assign n25475 =  ( wr_addr ) == ( bv_8_212_n493 )  ;
assign n25476 =  ( n25474 ) & (n25475 )  ;
assign n25477 =  ( n25476 ) & (wr )  ;
assign n25478 =  ( n25477 ) ? ( n5204 ) : ( iram_212 ) ;
assign n25479 = wr_addr[7:7] ;
assign n25480 =  ( n25479 ) == ( bv_1_0_n53 )  ;
assign n25481 =  ( wr_addr ) == ( bv_8_212_n493 )  ;
assign n25482 =  ( n25480 ) & (n25481 )  ;
assign n25483 =  ( n25482 ) & (wr )  ;
assign n25484 =  ( n25483 ) ? ( n5262 ) : ( iram_212 ) ;
assign n25485 = wr_addr[7:7] ;
assign n25486 =  ( n25485 ) == ( bv_1_0_n53 )  ;
assign n25487 =  ( wr_addr ) == ( bv_8_212_n493 )  ;
assign n25488 =  ( n25486 ) & (n25487 )  ;
assign n25489 =  ( n25488 ) & (wr )  ;
assign n25490 =  ( n25489 ) ? ( n5298 ) : ( iram_212 ) ;
assign n25491 = wr_addr[7:7] ;
assign n25492 =  ( n25491 ) == ( bv_1_0_n53 )  ;
assign n25493 =  ( wr_addr ) == ( bv_8_212_n493 )  ;
assign n25494 =  ( n25492 ) & (n25493 )  ;
assign n25495 =  ( n25494 ) & (wr )  ;
assign n25496 =  ( n25495 ) ? ( n5325 ) : ( iram_212 ) ;
assign n25497 = wr_addr[7:7] ;
assign n25498 =  ( n25497 ) == ( bv_1_0_n53 )  ;
assign n25499 =  ( wr_addr ) == ( bv_8_213_n495 )  ;
assign n25500 =  ( n25498 ) & (n25499 )  ;
assign n25501 =  ( n25500 ) & (wr )  ;
assign n25502 =  ( n25501 ) ? ( n4782 ) : ( iram_213 ) ;
assign n25503 = wr_addr[7:7] ;
assign n25504 =  ( n25503 ) == ( bv_1_0_n53 )  ;
assign n25505 =  ( wr_addr ) == ( bv_8_213_n495 )  ;
assign n25506 =  ( n25504 ) & (n25505 )  ;
assign n25507 =  ( n25506 ) & (wr )  ;
assign n25508 =  ( n25507 ) ? ( n4841 ) : ( iram_213 ) ;
assign n25509 = wr_addr[7:7] ;
assign n25510 =  ( n25509 ) == ( bv_1_0_n53 )  ;
assign n25511 =  ( wr_addr ) == ( bv_8_213_n495 )  ;
assign n25512 =  ( n25510 ) & (n25511 )  ;
assign n25513 =  ( n25512 ) & (wr )  ;
assign n25514 =  ( n25513 ) ? ( n5449 ) : ( iram_213 ) ;
assign n25515 = wr_addr[7:7] ;
assign n25516 =  ( n25515 ) == ( bv_1_0_n53 )  ;
assign n25517 =  ( wr_addr ) == ( bv_8_213_n495 )  ;
assign n25518 =  ( n25516 ) & (n25517 )  ;
assign n25519 =  ( n25518 ) & (wr )  ;
assign n25520 =  ( n25519 ) ? ( n4906 ) : ( iram_213 ) ;
assign n25521 = wr_addr[7:7] ;
assign n25522 =  ( n25521 ) == ( bv_1_0_n53 )  ;
assign n25523 =  ( wr_addr ) == ( bv_8_213_n495 )  ;
assign n25524 =  ( n25522 ) & (n25523 )  ;
assign n25525 =  ( n25524 ) & (wr )  ;
assign n25526 =  ( n25525 ) ? ( n5485 ) : ( iram_213 ) ;
assign n25527 = wr_addr[7:7] ;
assign n25528 =  ( n25527 ) == ( bv_1_0_n53 )  ;
assign n25529 =  ( wr_addr ) == ( bv_8_213_n495 )  ;
assign n25530 =  ( n25528 ) & (n25529 )  ;
assign n25531 =  ( n25530 ) & (wr )  ;
assign n25532 =  ( n25531 ) ? ( n5512 ) : ( iram_213 ) ;
assign n25533 = wr_addr[7:7] ;
assign n25534 =  ( n25533 ) == ( bv_1_0_n53 )  ;
assign n25535 =  ( wr_addr ) == ( bv_8_213_n495 )  ;
assign n25536 =  ( n25534 ) & (n25535 )  ;
assign n25537 =  ( n25536 ) & (wr )  ;
assign n25538 =  ( n25537 ) ? ( bv_8_0_n69 ) : ( iram_213 ) ;
assign n25539 = wr_addr[7:7] ;
assign n25540 =  ( n25539 ) == ( bv_1_0_n53 )  ;
assign n25541 =  ( wr_addr ) == ( bv_8_213_n495 )  ;
assign n25542 =  ( n25540 ) & (n25541 )  ;
assign n25543 =  ( n25542 ) & (wr )  ;
assign n25544 =  ( n25543 ) ? ( n5071 ) : ( iram_213 ) ;
assign n25545 = wr_addr[7:7] ;
assign n25546 =  ( n25545 ) == ( bv_1_0_n53 )  ;
assign n25547 =  ( wr_addr ) == ( bv_8_213_n495 )  ;
assign n25548 =  ( n25546 ) & (n25547 )  ;
assign n25549 =  ( n25548 ) & (wr )  ;
assign n25550 =  ( n25549 ) ? ( n5096 ) : ( iram_213 ) ;
assign n25551 = wr_addr[7:7] ;
assign n25552 =  ( n25551 ) == ( bv_1_0_n53 )  ;
assign n25553 =  ( wr_addr ) == ( bv_8_213_n495 )  ;
assign n25554 =  ( n25552 ) & (n25553 )  ;
assign n25555 =  ( n25554 ) & (wr )  ;
assign n25556 =  ( n25555 ) ? ( n5123 ) : ( iram_213 ) ;
assign n25557 = wr_addr[7:7] ;
assign n25558 =  ( n25557 ) == ( bv_1_0_n53 )  ;
assign n25559 =  ( wr_addr ) == ( bv_8_213_n495 )  ;
assign n25560 =  ( n25558 ) & (n25559 )  ;
assign n25561 =  ( n25560 ) & (wr )  ;
assign n25562 =  ( n25561 ) ? ( n5165 ) : ( iram_213 ) ;
assign n25563 = wr_addr[7:7] ;
assign n25564 =  ( n25563 ) == ( bv_1_0_n53 )  ;
assign n25565 =  ( wr_addr ) == ( bv_8_213_n495 )  ;
assign n25566 =  ( n25564 ) & (n25565 )  ;
assign n25567 =  ( n25566 ) & (wr )  ;
assign n25568 =  ( n25567 ) ? ( n5204 ) : ( iram_213 ) ;
assign n25569 = wr_addr[7:7] ;
assign n25570 =  ( n25569 ) == ( bv_1_0_n53 )  ;
assign n25571 =  ( wr_addr ) == ( bv_8_213_n495 )  ;
assign n25572 =  ( n25570 ) & (n25571 )  ;
assign n25573 =  ( n25572 ) & (wr )  ;
assign n25574 =  ( n25573 ) ? ( n5262 ) : ( iram_213 ) ;
assign n25575 = wr_addr[7:7] ;
assign n25576 =  ( n25575 ) == ( bv_1_0_n53 )  ;
assign n25577 =  ( wr_addr ) == ( bv_8_213_n495 )  ;
assign n25578 =  ( n25576 ) & (n25577 )  ;
assign n25579 =  ( n25578 ) & (wr )  ;
assign n25580 =  ( n25579 ) ? ( n5298 ) : ( iram_213 ) ;
assign n25581 = wr_addr[7:7] ;
assign n25582 =  ( n25581 ) == ( bv_1_0_n53 )  ;
assign n25583 =  ( wr_addr ) == ( bv_8_213_n495 )  ;
assign n25584 =  ( n25582 ) & (n25583 )  ;
assign n25585 =  ( n25584 ) & (wr )  ;
assign n25586 =  ( n25585 ) ? ( n5325 ) : ( iram_213 ) ;
assign n25587 = wr_addr[7:7] ;
assign n25588 =  ( n25587 ) == ( bv_1_0_n53 )  ;
assign n25589 =  ( wr_addr ) == ( bv_8_214_n497 )  ;
assign n25590 =  ( n25588 ) & (n25589 )  ;
assign n25591 =  ( n25590 ) & (wr )  ;
assign n25592 =  ( n25591 ) ? ( n4782 ) : ( iram_214 ) ;
assign n25593 = wr_addr[7:7] ;
assign n25594 =  ( n25593 ) == ( bv_1_0_n53 )  ;
assign n25595 =  ( wr_addr ) == ( bv_8_214_n497 )  ;
assign n25596 =  ( n25594 ) & (n25595 )  ;
assign n25597 =  ( n25596 ) & (wr )  ;
assign n25598 =  ( n25597 ) ? ( n4841 ) : ( iram_214 ) ;
assign n25599 = wr_addr[7:7] ;
assign n25600 =  ( n25599 ) == ( bv_1_0_n53 )  ;
assign n25601 =  ( wr_addr ) == ( bv_8_214_n497 )  ;
assign n25602 =  ( n25600 ) & (n25601 )  ;
assign n25603 =  ( n25602 ) & (wr )  ;
assign n25604 =  ( n25603 ) ? ( n5449 ) : ( iram_214 ) ;
assign n25605 = wr_addr[7:7] ;
assign n25606 =  ( n25605 ) == ( bv_1_0_n53 )  ;
assign n25607 =  ( wr_addr ) == ( bv_8_214_n497 )  ;
assign n25608 =  ( n25606 ) & (n25607 )  ;
assign n25609 =  ( n25608 ) & (wr )  ;
assign n25610 =  ( n25609 ) ? ( n4906 ) : ( iram_214 ) ;
assign n25611 = wr_addr[7:7] ;
assign n25612 =  ( n25611 ) == ( bv_1_0_n53 )  ;
assign n25613 =  ( wr_addr ) == ( bv_8_214_n497 )  ;
assign n25614 =  ( n25612 ) & (n25613 )  ;
assign n25615 =  ( n25614 ) & (wr )  ;
assign n25616 =  ( n25615 ) ? ( n5485 ) : ( iram_214 ) ;
assign n25617 = wr_addr[7:7] ;
assign n25618 =  ( n25617 ) == ( bv_1_0_n53 )  ;
assign n25619 =  ( wr_addr ) == ( bv_8_214_n497 )  ;
assign n25620 =  ( n25618 ) & (n25619 )  ;
assign n25621 =  ( n25620 ) & (wr )  ;
assign n25622 =  ( n25621 ) ? ( n5512 ) : ( iram_214 ) ;
assign n25623 = wr_addr[7:7] ;
assign n25624 =  ( n25623 ) == ( bv_1_0_n53 )  ;
assign n25625 =  ( wr_addr ) == ( bv_8_214_n497 )  ;
assign n25626 =  ( n25624 ) & (n25625 )  ;
assign n25627 =  ( n25626 ) & (wr )  ;
assign n25628 =  ( n25627 ) ? ( bv_8_0_n69 ) : ( iram_214 ) ;
assign n25629 = wr_addr[7:7] ;
assign n25630 =  ( n25629 ) == ( bv_1_0_n53 )  ;
assign n25631 =  ( wr_addr ) == ( bv_8_214_n497 )  ;
assign n25632 =  ( n25630 ) & (n25631 )  ;
assign n25633 =  ( n25632 ) & (wr )  ;
assign n25634 =  ( n25633 ) ? ( n5071 ) : ( iram_214 ) ;
assign n25635 = wr_addr[7:7] ;
assign n25636 =  ( n25635 ) == ( bv_1_0_n53 )  ;
assign n25637 =  ( wr_addr ) == ( bv_8_214_n497 )  ;
assign n25638 =  ( n25636 ) & (n25637 )  ;
assign n25639 =  ( n25638 ) & (wr )  ;
assign n25640 =  ( n25639 ) ? ( n5096 ) : ( iram_214 ) ;
assign n25641 = wr_addr[7:7] ;
assign n25642 =  ( n25641 ) == ( bv_1_0_n53 )  ;
assign n25643 =  ( wr_addr ) == ( bv_8_214_n497 )  ;
assign n25644 =  ( n25642 ) & (n25643 )  ;
assign n25645 =  ( n25644 ) & (wr )  ;
assign n25646 =  ( n25645 ) ? ( n5123 ) : ( iram_214 ) ;
assign n25647 = wr_addr[7:7] ;
assign n25648 =  ( n25647 ) == ( bv_1_0_n53 )  ;
assign n25649 =  ( wr_addr ) == ( bv_8_214_n497 )  ;
assign n25650 =  ( n25648 ) & (n25649 )  ;
assign n25651 =  ( n25650 ) & (wr )  ;
assign n25652 =  ( n25651 ) ? ( n5165 ) : ( iram_214 ) ;
assign n25653 = wr_addr[7:7] ;
assign n25654 =  ( n25653 ) == ( bv_1_0_n53 )  ;
assign n25655 =  ( wr_addr ) == ( bv_8_214_n497 )  ;
assign n25656 =  ( n25654 ) & (n25655 )  ;
assign n25657 =  ( n25656 ) & (wr )  ;
assign n25658 =  ( n25657 ) ? ( n5204 ) : ( iram_214 ) ;
assign n25659 = wr_addr[7:7] ;
assign n25660 =  ( n25659 ) == ( bv_1_0_n53 )  ;
assign n25661 =  ( wr_addr ) == ( bv_8_214_n497 )  ;
assign n25662 =  ( n25660 ) & (n25661 )  ;
assign n25663 =  ( n25662 ) & (wr )  ;
assign n25664 =  ( n25663 ) ? ( n5262 ) : ( iram_214 ) ;
assign n25665 = wr_addr[7:7] ;
assign n25666 =  ( n25665 ) == ( bv_1_0_n53 )  ;
assign n25667 =  ( wr_addr ) == ( bv_8_214_n497 )  ;
assign n25668 =  ( n25666 ) & (n25667 )  ;
assign n25669 =  ( n25668 ) & (wr )  ;
assign n25670 =  ( n25669 ) ? ( n5298 ) : ( iram_214 ) ;
assign n25671 = wr_addr[7:7] ;
assign n25672 =  ( n25671 ) == ( bv_1_0_n53 )  ;
assign n25673 =  ( wr_addr ) == ( bv_8_214_n497 )  ;
assign n25674 =  ( n25672 ) & (n25673 )  ;
assign n25675 =  ( n25674 ) & (wr )  ;
assign n25676 =  ( n25675 ) ? ( n5325 ) : ( iram_214 ) ;
assign n25677 = wr_addr[7:7] ;
assign n25678 =  ( n25677 ) == ( bv_1_0_n53 )  ;
assign n25679 =  ( wr_addr ) == ( bv_8_215_n499 )  ;
assign n25680 =  ( n25678 ) & (n25679 )  ;
assign n25681 =  ( n25680 ) & (wr )  ;
assign n25682 =  ( n25681 ) ? ( n4782 ) : ( iram_215 ) ;
assign n25683 = wr_addr[7:7] ;
assign n25684 =  ( n25683 ) == ( bv_1_0_n53 )  ;
assign n25685 =  ( wr_addr ) == ( bv_8_215_n499 )  ;
assign n25686 =  ( n25684 ) & (n25685 )  ;
assign n25687 =  ( n25686 ) & (wr )  ;
assign n25688 =  ( n25687 ) ? ( n4841 ) : ( iram_215 ) ;
assign n25689 = wr_addr[7:7] ;
assign n25690 =  ( n25689 ) == ( bv_1_0_n53 )  ;
assign n25691 =  ( wr_addr ) == ( bv_8_215_n499 )  ;
assign n25692 =  ( n25690 ) & (n25691 )  ;
assign n25693 =  ( n25692 ) & (wr )  ;
assign n25694 =  ( n25693 ) ? ( n5449 ) : ( iram_215 ) ;
assign n25695 = wr_addr[7:7] ;
assign n25696 =  ( n25695 ) == ( bv_1_0_n53 )  ;
assign n25697 =  ( wr_addr ) == ( bv_8_215_n499 )  ;
assign n25698 =  ( n25696 ) & (n25697 )  ;
assign n25699 =  ( n25698 ) & (wr )  ;
assign n25700 =  ( n25699 ) ? ( n4906 ) : ( iram_215 ) ;
assign n25701 = wr_addr[7:7] ;
assign n25702 =  ( n25701 ) == ( bv_1_0_n53 )  ;
assign n25703 =  ( wr_addr ) == ( bv_8_215_n499 )  ;
assign n25704 =  ( n25702 ) & (n25703 )  ;
assign n25705 =  ( n25704 ) & (wr )  ;
assign n25706 =  ( n25705 ) ? ( n5485 ) : ( iram_215 ) ;
assign n25707 = wr_addr[7:7] ;
assign n25708 =  ( n25707 ) == ( bv_1_0_n53 )  ;
assign n25709 =  ( wr_addr ) == ( bv_8_215_n499 )  ;
assign n25710 =  ( n25708 ) & (n25709 )  ;
assign n25711 =  ( n25710 ) & (wr )  ;
assign n25712 =  ( n25711 ) ? ( n5512 ) : ( iram_215 ) ;
assign n25713 = wr_addr[7:7] ;
assign n25714 =  ( n25713 ) == ( bv_1_0_n53 )  ;
assign n25715 =  ( wr_addr ) == ( bv_8_215_n499 )  ;
assign n25716 =  ( n25714 ) & (n25715 )  ;
assign n25717 =  ( n25716 ) & (wr )  ;
assign n25718 =  ( n25717 ) ? ( bv_8_0_n69 ) : ( iram_215 ) ;
assign n25719 = wr_addr[7:7] ;
assign n25720 =  ( n25719 ) == ( bv_1_0_n53 )  ;
assign n25721 =  ( wr_addr ) == ( bv_8_215_n499 )  ;
assign n25722 =  ( n25720 ) & (n25721 )  ;
assign n25723 =  ( n25722 ) & (wr )  ;
assign n25724 =  ( n25723 ) ? ( n5071 ) : ( iram_215 ) ;
assign n25725 = wr_addr[7:7] ;
assign n25726 =  ( n25725 ) == ( bv_1_0_n53 )  ;
assign n25727 =  ( wr_addr ) == ( bv_8_215_n499 )  ;
assign n25728 =  ( n25726 ) & (n25727 )  ;
assign n25729 =  ( n25728 ) & (wr )  ;
assign n25730 =  ( n25729 ) ? ( n5096 ) : ( iram_215 ) ;
assign n25731 = wr_addr[7:7] ;
assign n25732 =  ( n25731 ) == ( bv_1_0_n53 )  ;
assign n25733 =  ( wr_addr ) == ( bv_8_215_n499 )  ;
assign n25734 =  ( n25732 ) & (n25733 )  ;
assign n25735 =  ( n25734 ) & (wr )  ;
assign n25736 =  ( n25735 ) ? ( n5123 ) : ( iram_215 ) ;
assign n25737 = wr_addr[7:7] ;
assign n25738 =  ( n25737 ) == ( bv_1_0_n53 )  ;
assign n25739 =  ( wr_addr ) == ( bv_8_215_n499 )  ;
assign n25740 =  ( n25738 ) & (n25739 )  ;
assign n25741 =  ( n25740 ) & (wr )  ;
assign n25742 =  ( n25741 ) ? ( n5165 ) : ( iram_215 ) ;
assign n25743 = wr_addr[7:7] ;
assign n25744 =  ( n25743 ) == ( bv_1_0_n53 )  ;
assign n25745 =  ( wr_addr ) == ( bv_8_215_n499 )  ;
assign n25746 =  ( n25744 ) & (n25745 )  ;
assign n25747 =  ( n25746 ) & (wr )  ;
assign n25748 =  ( n25747 ) ? ( n5204 ) : ( iram_215 ) ;
assign n25749 = wr_addr[7:7] ;
assign n25750 =  ( n25749 ) == ( bv_1_0_n53 )  ;
assign n25751 =  ( wr_addr ) == ( bv_8_215_n499 )  ;
assign n25752 =  ( n25750 ) & (n25751 )  ;
assign n25753 =  ( n25752 ) & (wr )  ;
assign n25754 =  ( n25753 ) ? ( n5262 ) : ( iram_215 ) ;
assign n25755 = wr_addr[7:7] ;
assign n25756 =  ( n25755 ) == ( bv_1_0_n53 )  ;
assign n25757 =  ( wr_addr ) == ( bv_8_215_n499 )  ;
assign n25758 =  ( n25756 ) & (n25757 )  ;
assign n25759 =  ( n25758 ) & (wr )  ;
assign n25760 =  ( n25759 ) ? ( n5298 ) : ( iram_215 ) ;
assign n25761 = wr_addr[7:7] ;
assign n25762 =  ( n25761 ) == ( bv_1_0_n53 )  ;
assign n25763 =  ( wr_addr ) == ( bv_8_215_n499 )  ;
assign n25764 =  ( n25762 ) & (n25763 )  ;
assign n25765 =  ( n25764 ) & (wr )  ;
assign n25766 =  ( n25765 ) ? ( n5325 ) : ( iram_215 ) ;
assign n25767 = wr_addr[7:7] ;
assign n25768 =  ( n25767 ) == ( bv_1_0_n53 )  ;
assign n25769 =  ( wr_addr ) == ( bv_8_216_n501 )  ;
assign n25770 =  ( n25768 ) & (n25769 )  ;
assign n25771 =  ( n25770 ) & (wr )  ;
assign n25772 =  ( n25771 ) ? ( n4782 ) : ( iram_216 ) ;
assign n25773 = wr_addr[7:7] ;
assign n25774 =  ( n25773 ) == ( bv_1_0_n53 )  ;
assign n25775 =  ( wr_addr ) == ( bv_8_216_n501 )  ;
assign n25776 =  ( n25774 ) & (n25775 )  ;
assign n25777 =  ( n25776 ) & (wr )  ;
assign n25778 =  ( n25777 ) ? ( n4841 ) : ( iram_216 ) ;
assign n25779 = wr_addr[7:7] ;
assign n25780 =  ( n25779 ) == ( bv_1_0_n53 )  ;
assign n25781 =  ( wr_addr ) == ( bv_8_216_n501 )  ;
assign n25782 =  ( n25780 ) & (n25781 )  ;
assign n25783 =  ( n25782 ) & (wr )  ;
assign n25784 =  ( n25783 ) ? ( n5449 ) : ( iram_216 ) ;
assign n25785 = wr_addr[7:7] ;
assign n25786 =  ( n25785 ) == ( bv_1_0_n53 )  ;
assign n25787 =  ( wr_addr ) == ( bv_8_216_n501 )  ;
assign n25788 =  ( n25786 ) & (n25787 )  ;
assign n25789 =  ( n25788 ) & (wr )  ;
assign n25790 =  ( n25789 ) ? ( n4906 ) : ( iram_216 ) ;
assign n25791 = wr_addr[7:7] ;
assign n25792 =  ( n25791 ) == ( bv_1_0_n53 )  ;
assign n25793 =  ( wr_addr ) == ( bv_8_216_n501 )  ;
assign n25794 =  ( n25792 ) & (n25793 )  ;
assign n25795 =  ( n25794 ) & (wr )  ;
assign n25796 =  ( n25795 ) ? ( n5485 ) : ( iram_216 ) ;
assign n25797 = wr_addr[7:7] ;
assign n25798 =  ( n25797 ) == ( bv_1_0_n53 )  ;
assign n25799 =  ( wr_addr ) == ( bv_8_216_n501 )  ;
assign n25800 =  ( n25798 ) & (n25799 )  ;
assign n25801 =  ( n25800 ) & (wr )  ;
assign n25802 =  ( n25801 ) ? ( n5512 ) : ( iram_216 ) ;
assign n25803 = wr_addr[7:7] ;
assign n25804 =  ( n25803 ) == ( bv_1_0_n53 )  ;
assign n25805 =  ( wr_addr ) == ( bv_8_216_n501 )  ;
assign n25806 =  ( n25804 ) & (n25805 )  ;
assign n25807 =  ( n25806 ) & (wr )  ;
assign n25808 =  ( n25807 ) ? ( bv_8_0_n69 ) : ( iram_216 ) ;
assign n25809 = wr_addr[7:7] ;
assign n25810 =  ( n25809 ) == ( bv_1_0_n53 )  ;
assign n25811 =  ( wr_addr ) == ( bv_8_216_n501 )  ;
assign n25812 =  ( n25810 ) & (n25811 )  ;
assign n25813 =  ( n25812 ) & (wr )  ;
assign n25814 =  ( n25813 ) ? ( n5071 ) : ( iram_216 ) ;
assign n25815 = wr_addr[7:7] ;
assign n25816 =  ( n25815 ) == ( bv_1_0_n53 )  ;
assign n25817 =  ( wr_addr ) == ( bv_8_216_n501 )  ;
assign n25818 =  ( n25816 ) & (n25817 )  ;
assign n25819 =  ( n25818 ) & (wr )  ;
assign n25820 =  ( n25819 ) ? ( n5096 ) : ( iram_216 ) ;
assign n25821 = wr_addr[7:7] ;
assign n25822 =  ( n25821 ) == ( bv_1_0_n53 )  ;
assign n25823 =  ( wr_addr ) == ( bv_8_216_n501 )  ;
assign n25824 =  ( n25822 ) & (n25823 )  ;
assign n25825 =  ( n25824 ) & (wr )  ;
assign n25826 =  ( n25825 ) ? ( n5123 ) : ( iram_216 ) ;
assign n25827 = wr_addr[7:7] ;
assign n25828 =  ( n25827 ) == ( bv_1_0_n53 )  ;
assign n25829 =  ( wr_addr ) == ( bv_8_216_n501 )  ;
assign n25830 =  ( n25828 ) & (n25829 )  ;
assign n25831 =  ( n25830 ) & (wr )  ;
assign n25832 =  ( n25831 ) ? ( n5165 ) : ( iram_216 ) ;
assign n25833 = wr_addr[7:7] ;
assign n25834 =  ( n25833 ) == ( bv_1_0_n53 )  ;
assign n25835 =  ( wr_addr ) == ( bv_8_216_n501 )  ;
assign n25836 =  ( n25834 ) & (n25835 )  ;
assign n25837 =  ( n25836 ) & (wr )  ;
assign n25838 =  ( n25837 ) ? ( n5204 ) : ( iram_216 ) ;
assign n25839 = wr_addr[7:7] ;
assign n25840 =  ( n25839 ) == ( bv_1_0_n53 )  ;
assign n25841 =  ( wr_addr ) == ( bv_8_216_n501 )  ;
assign n25842 =  ( n25840 ) & (n25841 )  ;
assign n25843 =  ( n25842 ) & (wr )  ;
assign n25844 =  ( n25843 ) ? ( n5262 ) : ( iram_216 ) ;
assign n25845 = wr_addr[7:7] ;
assign n25846 =  ( n25845 ) == ( bv_1_0_n53 )  ;
assign n25847 =  ( wr_addr ) == ( bv_8_216_n501 )  ;
assign n25848 =  ( n25846 ) & (n25847 )  ;
assign n25849 =  ( n25848 ) & (wr )  ;
assign n25850 =  ( n25849 ) ? ( n5298 ) : ( iram_216 ) ;
assign n25851 = wr_addr[7:7] ;
assign n25852 =  ( n25851 ) == ( bv_1_0_n53 )  ;
assign n25853 =  ( wr_addr ) == ( bv_8_216_n501 )  ;
assign n25854 =  ( n25852 ) & (n25853 )  ;
assign n25855 =  ( n25854 ) & (wr )  ;
assign n25856 =  ( n25855 ) ? ( n5325 ) : ( iram_216 ) ;
assign n25857 = wr_addr[7:7] ;
assign n25858 =  ( n25857 ) == ( bv_1_0_n53 )  ;
assign n25859 =  ( wr_addr ) == ( bv_8_217_n503 )  ;
assign n25860 =  ( n25858 ) & (n25859 )  ;
assign n25861 =  ( n25860 ) & (wr )  ;
assign n25862 =  ( n25861 ) ? ( n4782 ) : ( iram_217 ) ;
assign n25863 = wr_addr[7:7] ;
assign n25864 =  ( n25863 ) == ( bv_1_0_n53 )  ;
assign n25865 =  ( wr_addr ) == ( bv_8_217_n503 )  ;
assign n25866 =  ( n25864 ) & (n25865 )  ;
assign n25867 =  ( n25866 ) & (wr )  ;
assign n25868 =  ( n25867 ) ? ( n4841 ) : ( iram_217 ) ;
assign n25869 = wr_addr[7:7] ;
assign n25870 =  ( n25869 ) == ( bv_1_0_n53 )  ;
assign n25871 =  ( wr_addr ) == ( bv_8_217_n503 )  ;
assign n25872 =  ( n25870 ) & (n25871 )  ;
assign n25873 =  ( n25872 ) & (wr )  ;
assign n25874 =  ( n25873 ) ? ( n5449 ) : ( iram_217 ) ;
assign n25875 = wr_addr[7:7] ;
assign n25876 =  ( n25875 ) == ( bv_1_0_n53 )  ;
assign n25877 =  ( wr_addr ) == ( bv_8_217_n503 )  ;
assign n25878 =  ( n25876 ) & (n25877 )  ;
assign n25879 =  ( n25878 ) & (wr )  ;
assign n25880 =  ( n25879 ) ? ( n4906 ) : ( iram_217 ) ;
assign n25881 = wr_addr[7:7] ;
assign n25882 =  ( n25881 ) == ( bv_1_0_n53 )  ;
assign n25883 =  ( wr_addr ) == ( bv_8_217_n503 )  ;
assign n25884 =  ( n25882 ) & (n25883 )  ;
assign n25885 =  ( n25884 ) & (wr )  ;
assign n25886 =  ( n25885 ) ? ( n5485 ) : ( iram_217 ) ;
assign n25887 = wr_addr[7:7] ;
assign n25888 =  ( n25887 ) == ( bv_1_0_n53 )  ;
assign n25889 =  ( wr_addr ) == ( bv_8_217_n503 )  ;
assign n25890 =  ( n25888 ) & (n25889 )  ;
assign n25891 =  ( n25890 ) & (wr )  ;
assign n25892 =  ( n25891 ) ? ( n5512 ) : ( iram_217 ) ;
assign n25893 = wr_addr[7:7] ;
assign n25894 =  ( n25893 ) == ( bv_1_0_n53 )  ;
assign n25895 =  ( wr_addr ) == ( bv_8_217_n503 )  ;
assign n25896 =  ( n25894 ) & (n25895 )  ;
assign n25897 =  ( n25896 ) & (wr )  ;
assign n25898 =  ( n25897 ) ? ( bv_8_0_n69 ) : ( iram_217 ) ;
assign n25899 = wr_addr[7:7] ;
assign n25900 =  ( n25899 ) == ( bv_1_0_n53 )  ;
assign n25901 =  ( wr_addr ) == ( bv_8_217_n503 )  ;
assign n25902 =  ( n25900 ) & (n25901 )  ;
assign n25903 =  ( n25902 ) & (wr )  ;
assign n25904 =  ( n25903 ) ? ( n5071 ) : ( iram_217 ) ;
assign n25905 = wr_addr[7:7] ;
assign n25906 =  ( n25905 ) == ( bv_1_0_n53 )  ;
assign n25907 =  ( wr_addr ) == ( bv_8_217_n503 )  ;
assign n25908 =  ( n25906 ) & (n25907 )  ;
assign n25909 =  ( n25908 ) & (wr )  ;
assign n25910 =  ( n25909 ) ? ( n5096 ) : ( iram_217 ) ;
assign n25911 = wr_addr[7:7] ;
assign n25912 =  ( n25911 ) == ( bv_1_0_n53 )  ;
assign n25913 =  ( wr_addr ) == ( bv_8_217_n503 )  ;
assign n25914 =  ( n25912 ) & (n25913 )  ;
assign n25915 =  ( n25914 ) & (wr )  ;
assign n25916 =  ( n25915 ) ? ( n5123 ) : ( iram_217 ) ;
assign n25917 = wr_addr[7:7] ;
assign n25918 =  ( n25917 ) == ( bv_1_0_n53 )  ;
assign n25919 =  ( wr_addr ) == ( bv_8_217_n503 )  ;
assign n25920 =  ( n25918 ) & (n25919 )  ;
assign n25921 =  ( n25920 ) & (wr )  ;
assign n25922 =  ( n25921 ) ? ( n5165 ) : ( iram_217 ) ;
assign n25923 = wr_addr[7:7] ;
assign n25924 =  ( n25923 ) == ( bv_1_0_n53 )  ;
assign n25925 =  ( wr_addr ) == ( bv_8_217_n503 )  ;
assign n25926 =  ( n25924 ) & (n25925 )  ;
assign n25927 =  ( n25926 ) & (wr )  ;
assign n25928 =  ( n25927 ) ? ( n5204 ) : ( iram_217 ) ;
assign n25929 = wr_addr[7:7] ;
assign n25930 =  ( n25929 ) == ( bv_1_0_n53 )  ;
assign n25931 =  ( wr_addr ) == ( bv_8_217_n503 )  ;
assign n25932 =  ( n25930 ) & (n25931 )  ;
assign n25933 =  ( n25932 ) & (wr )  ;
assign n25934 =  ( n25933 ) ? ( n5262 ) : ( iram_217 ) ;
assign n25935 = wr_addr[7:7] ;
assign n25936 =  ( n25935 ) == ( bv_1_0_n53 )  ;
assign n25937 =  ( wr_addr ) == ( bv_8_217_n503 )  ;
assign n25938 =  ( n25936 ) & (n25937 )  ;
assign n25939 =  ( n25938 ) & (wr )  ;
assign n25940 =  ( n25939 ) ? ( n5298 ) : ( iram_217 ) ;
assign n25941 = wr_addr[7:7] ;
assign n25942 =  ( n25941 ) == ( bv_1_0_n53 )  ;
assign n25943 =  ( wr_addr ) == ( bv_8_217_n503 )  ;
assign n25944 =  ( n25942 ) & (n25943 )  ;
assign n25945 =  ( n25944 ) & (wr )  ;
assign n25946 =  ( n25945 ) ? ( n5325 ) : ( iram_217 ) ;
assign n25947 = wr_addr[7:7] ;
assign n25948 =  ( n25947 ) == ( bv_1_0_n53 )  ;
assign n25949 =  ( wr_addr ) == ( bv_8_218_n505 )  ;
assign n25950 =  ( n25948 ) & (n25949 )  ;
assign n25951 =  ( n25950 ) & (wr )  ;
assign n25952 =  ( n25951 ) ? ( n4782 ) : ( iram_218 ) ;
assign n25953 = wr_addr[7:7] ;
assign n25954 =  ( n25953 ) == ( bv_1_0_n53 )  ;
assign n25955 =  ( wr_addr ) == ( bv_8_218_n505 )  ;
assign n25956 =  ( n25954 ) & (n25955 )  ;
assign n25957 =  ( n25956 ) & (wr )  ;
assign n25958 =  ( n25957 ) ? ( n4841 ) : ( iram_218 ) ;
assign n25959 = wr_addr[7:7] ;
assign n25960 =  ( n25959 ) == ( bv_1_0_n53 )  ;
assign n25961 =  ( wr_addr ) == ( bv_8_218_n505 )  ;
assign n25962 =  ( n25960 ) & (n25961 )  ;
assign n25963 =  ( n25962 ) & (wr )  ;
assign n25964 =  ( n25963 ) ? ( n5449 ) : ( iram_218 ) ;
assign n25965 = wr_addr[7:7] ;
assign n25966 =  ( n25965 ) == ( bv_1_0_n53 )  ;
assign n25967 =  ( wr_addr ) == ( bv_8_218_n505 )  ;
assign n25968 =  ( n25966 ) & (n25967 )  ;
assign n25969 =  ( n25968 ) & (wr )  ;
assign n25970 =  ( n25969 ) ? ( n4906 ) : ( iram_218 ) ;
assign n25971 = wr_addr[7:7] ;
assign n25972 =  ( n25971 ) == ( bv_1_0_n53 )  ;
assign n25973 =  ( wr_addr ) == ( bv_8_218_n505 )  ;
assign n25974 =  ( n25972 ) & (n25973 )  ;
assign n25975 =  ( n25974 ) & (wr )  ;
assign n25976 =  ( n25975 ) ? ( n5485 ) : ( iram_218 ) ;
assign n25977 = wr_addr[7:7] ;
assign n25978 =  ( n25977 ) == ( bv_1_0_n53 )  ;
assign n25979 =  ( wr_addr ) == ( bv_8_218_n505 )  ;
assign n25980 =  ( n25978 ) & (n25979 )  ;
assign n25981 =  ( n25980 ) & (wr )  ;
assign n25982 =  ( n25981 ) ? ( n5512 ) : ( iram_218 ) ;
assign n25983 = wr_addr[7:7] ;
assign n25984 =  ( n25983 ) == ( bv_1_0_n53 )  ;
assign n25985 =  ( wr_addr ) == ( bv_8_218_n505 )  ;
assign n25986 =  ( n25984 ) & (n25985 )  ;
assign n25987 =  ( n25986 ) & (wr )  ;
assign n25988 =  ( n25987 ) ? ( bv_8_0_n69 ) : ( iram_218 ) ;
assign n25989 = wr_addr[7:7] ;
assign n25990 =  ( n25989 ) == ( bv_1_0_n53 )  ;
assign n25991 =  ( wr_addr ) == ( bv_8_218_n505 )  ;
assign n25992 =  ( n25990 ) & (n25991 )  ;
assign n25993 =  ( n25992 ) & (wr )  ;
assign n25994 =  ( n25993 ) ? ( n5071 ) : ( iram_218 ) ;
assign n25995 = wr_addr[7:7] ;
assign n25996 =  ( n25995 ) == ( bv_1_0_n53 )  ;
assign n25997 =  ( wr_addr ) == ( bv_8_218_n505 )  ;
assign n25998 =  ( n25996 ) & (n25997 )  ;
assign n25999 =  ( n25998 ) & (wr )  ;
assign n26000 =  ( n25999 ) ? ( n5096 ) : ( iram_218 ) ;
assign n26001 = wr_addr[7:7] ;
assign n26002 =  ( n26001 ) == ( bv_1_0_n53 )  ;
assign n26003 =  ( wr_addr ) == ( bv_8_218_n505 )  ;
assign n26004 =  ( n26002 ) & (n26003 )  ;
assign n26005 =  ( n26004 ) & (wr )  ;
assign n26006 =  ( n26005 ) ? ( n5123 ) : ( iram_218 ) ;
assign n26007 = wr_addr[7:7] ;
assign n26008 =  ( n26007 ) == ( bv_1_0_n53 )  ;
assign n26009 =  ( wr_addr ) == ( bv_8_218_n505 )  ;
assign n26010 =  ( n26008 ) & (n26009 )  ;
assign n26011 =  ( n26010 ) & (wr )  ;
assign n26012 =  ( n26011 ) ? ( n5165 ) : ( iram_218 ) ;
assign n26013 = wr_addr[7:7] ;
assign n26014 =  ( n26013 ) == ( bv_1_0_n53 )  ;
assign n26015 =  ( wr_addr ) == ( bv_8_218_n505 )  ;
assign n26016 =  ( n26014 ) & (n26015 )  ;
assign n26017 =  ( n26016 ) & (wr )  ;
assign n26018 =  ( n26017 ) ? ( n5204 ) : ( iram_218 ) ;
assign n26019 = wr_addr[7:7] ;
assign n26020 =  ( n26019 ) == ( bv_1_0_n53 )  ;
assign n26021 =  ( wr_addr ) == ( bv_8_218_n505 )  ;
assign n26022 =  ( n26020 ) & (n26021 )  ;
assign n26023 =  ( n26022 ) & (wr )  ;
assign n26024 =  ( n26023 ) ? ( n5262 ) : ( iram_218 ) ;
assign n26025 = wr_addr[7:7] ;
assign n26026 =  ( n26025 ) == ( bv_1_0_n53 )  ;
assign n26027 =  ( wr_addr ) == ( bv_8_218_n505 )  ;
assign n26028 =  ( n26026 ) & (n26027 )  ;
assign n26029 =  ( n26028 ) & (wr )  ;
assign n26030 =  ( n26029 ) ? ( n5298 ) : ( iram_218 ) ;
assign n26031 = wr_addr[7:7] ;
assign n26032 =  ( n26031 ) == ( bv_1_0_n53 )  ;
assign n26033 =  ( wr_addr ) == ( bv_8_218_n505 )  ;
assign n26034 =  ( n26032 ) & (n26033 )  ;
assign n26035 =  ( n26034 ) & (wr )  ;
assign n26036 =  ( n26035 ) ? ( n5325 ) : ( iram_218 ) ;
assign n26037 = wr_addr[7:7] ;
assign n26038 =  ( n26037 ) == ( bv_1_0_n53 )  ;
assign n26039 =  ( wr_addr ) == ( bv_8_219_n507 )  ;
assign n26040 =  ( n26038 ) & (n26039 )  ;
assign n26041 =  ( n26040 ) & (wr )  ;
assign n26042 =  ( n26041 ) ? ( n4782 ) : ( iram_219 ) ;
assign n26043 = wr_addr[7:7] ;
assign n26044 =  ( n26043 ) == ( bv_1_0_n53 )  ;
assign n26045 =  ( wr_addr ) == ( bv_8_219_n507 )  ;
assign n26046 =  ( n26044 ) & (n26045 )  ;
assign n26047 =  ( n26046 ) & (wr )  ;
assign n26048 =  ( n26047 ) ? ( n4841 ) : ( iram_219 ) ;
assign n26049 = wr_addr[7:7] ;
assign n26050 =  ( n26049 ) == ( bv_1_0_n53 )  ;
assign n26051 =  ( wr_addr ) == ( bv_8_219_n507 )  ;
assign n26052 =  ( n26050 ) & (n26051 )  ;
assign n26053 =  ( n26052 ) & (wr )  ;
assign n26054 =  ( n26053 ) ? ( n5449 ) : ( iram_219 ) ;
assign n26055 = wr_addr[7:7] ;
assign n26056 =  ( n26055 ) == ( bv_1_0_n53 )  ;
assign n26057 =  ( wr_addr ) == ( bv_8_219_n507 )  ;
assign n26058 =  ( n26056 ) & (n26057 )  ;
assign n26059 =  ( n26058 ) & (wr )  ;
assign n26060 =  ( n26059 ) ? ( n4906 ) : ( iram_219 ) ;
assign n26061 = wr_addr[7:7] ;
assign n26062 =  ( n26061 ) == ( bv_1_0_n53 )  ;
assign n26063 =  ( wr_addr ) == ( bv_8_219_n507 )  ;
assign n26064 =  ( n26062 ) & (n26063 )  ;
assign n26065 =  ( n26064 ) & (wr )  ;
assign n26066 =  ( n26065 ) ? ( n5485 ) : ( iram_219 ) ;
assign n26067 = wr_addr[7:7] ;
assign n26068 =  ( n26067 ) == ( bv_1_0_n53 )  ;
assign n26069 =  ( wr_addr ) == ( bv_8_219_n507 )  ;
assign n26070 =  ( n26068 ) & (n26069 )  ;
assign n26071 =  ( n26070 ) & (wr )  ;
assign n26072 =  ( n26071 ) ? ( n5512 ) : ( iram_219 ) ;
assign n26073 = wr_addr[7:7] ;
assign n26074 =  ( n26073 ) == ( bv_1_0_n53 )  ;
assign n26075 =  ( wr_addr ) == ( bv_8_219_n507 )  ;
assign n26076 =  ( n26074 ) & (n26075 )  ;
assign n26077 =  ( n26076 ) & (wr )  ;
assign n26078 =  ( n26077 ) ? ( bv_8_0_n69 ) : ( iram_219 ) ;
assign n26079 = wr_addr[7:7] ;
assign n26080 =  ( n26079 ) == ( bv_1_0_n53 )  ;
assign n26081 =  ( wr_addr ) == ( bv_8_219_n507 )  ;
assign n26082 =  ( n26080 ) & (n26081 )  ;
assign n26083 =  ( n26082 ) & (wr )  ;
assign n26084 =  ( n26083 ) ? ( n5071 ) : ( iram_219 ) ;
assign n26085 = wr_addr[7:7] ;
assign n26086 =  ( n26085 ) == ( bv_1_0_n53 )  ;
assign n26087 =  ( wr_addr ) == ( bv_8_219_n507 )  ;
assign n26088 =  ( n26086 ) & (n26087 )  ;
assign n26089 =  ( n26088 ) & (wr )  ;
assign n26090 =  ( n26089 ) ? ( n5096 ) : ( iram_219 ) ;
assign n26091 = wr_addr[7:7] ;
assign n26092 =  ( n26091 ) == ( bv_1_0_n53 )  ;
assign n26093 =  ( wr_addr ) == ( bv_8_219_n507 )  ;
assign n26094 =  ( n26092 ) & (n26093 )  ;
assign n26095 =  ( n26094 ) & (wr )  ;
assign n26096 =  ( n26095 ) ? ( n5123 ) : ( iram_219 ) ;
assign n26097 = wr_addr[7:7] ;
assign n26098 =  ( n26097 ) == ( bv_1_0_n53 )  ;
assign n26099 =  ( wr_addr ) == ( bv_8_219_n507 )  ;
assign n26100 =  ( n26098 ) & (n26099 )  ;
assign n26101 =  ( n26100 ) & (wr )  ;
assign n26102 =  ( n26101 ) ? ( n5165 ) : ( iram_219 ) ;
assign n26103 = wr_addr[7:7] ;
assign n26104 =  ( n26103 ) == ( bv_1_0_n53 )  ;
assign n26105 =  ( wr_addr ) == ( bv_8_219_n507 )  ;
assign n26106 =  ( n26104 ) & (n26105 )  ;
assign n26107 =  ( n26106 ) & (wr )  ;
assign n26108 =  ( n26107 ) ? ( n5204 ) : ( iram_219 ) ;
assign n26109 = wr_addr[7:7] ;
assign n26110 =  ( n26109 ) == ( bv_1_0_n53 )  ;
assign n26111 =  ( wr_addr ) == ( bv_8_219_n507 )  ;
assign n26112 =  ( n26110 ) & (n26111 )  ;
assign n26113 =  ( n26112 ) & (wr )  ;
assign n26114 =  ( n26113 ) ? ( n5262 ) : ( iram_219 ) ;
assign n26115 = wr_addr[7:7] ;
assign n26116 =  ( n26115 ) == ( bv_1_0_n53 )  ;
assign n26117 =  ( wr_addr ) == ( bv_8_219_n507 )  ;
assign n26118 =  ( n26116 ) & (n26117 )  ;
assign n26119 =  ( n26118 ) & (wr )  ;
assign n26120 =  ( n26119 ) ? ( n5298 ) : ( iram_219 ) ;
assign n26121 = wr_addr[7:7] ;
assign n26122 =  ( n26121 ) == ( bv_1_0_n53 )  ;
assign n26123 =  ( wr_addr ) == ( bv_8_219_n507 )  ;
assign n26124 =  ( n26122 ) & (n26123 )  ;
assign n26125 =  ( n26124 ) & (wr )  ;
assign n26126 =  ( n26125 ) ? ( n5325 ) : ( iram_219 ) ;
assign n26127 = wr_addr[7:7] ;
assign n26128 =  ( n26127 ) == ( bv_1_0_n53 )  ;
assign n26129 =  ( wr_addr ) == ( bv_8_220_n509 )  ;
assign n26130 =  ( n26128 ) & (n26129 )  ;
assign n26131 =  ( n26130 ) & (wr )  ;
assign n26132 =  ( n26131 ) ? ( n4782 ) : ( iram_220 ) ;
assign n26133 = wr_addr[7:7] ;
assign n26134 =  ( n26133 ) == ( bv_1_0_n53 )  ;
assign n26135 =  ( wr_addr ) == ( bv_8_220_n509 )  ;
assign n26136 =  ( n26134 ) & (n26135 )  ;
assign n26137 =  ( n26136 ) & (wr )  ;
assign n26138 =  ( n26137 ) ? ( n4841 ) : ( iram_220 ) ;
assign n26139 = wr_addr[7:7] ;
assign n26140 =  ( n26139 ) == ( bv_1_0_n53 )  ;
assign n26141 =  ( wr_addr ) == ( bv_8_220_n509 )  ;
assign n26142 =  ( n26140 ) & (n26141 )  ;
assign n26143 =  ( n26142 ) & (wr )  ;
assign n26144 =  ( n26143 ) ? ( n5449 ) : ( iram_220 ) ;
assign n26145 = wr_addr[7:7] ;
assign n26146 =  ( n26145 ) == ( bv_1_0_n53 )  ;
assign n26147 =  ( wr_addr ) == ( bv_8_220_n509 )  ;
assign n26148 =  ( n26146 ) & (n26147 )  ;
assign n26149 =  ( n26148 ) & (wr )  ;
assign n26150 =  ( n26149 ) ? ( n4906 ) : ( iram_220 ) ;
assign n26151 = wr_addr[7:7] ;
assign n26152 =  ( n26151 ) == ( bv_1_0_n53 )  ;
assign n26153 =  ( wr_addr ) == ( bv_8_220_n509 )  ;
assign n26154 =  ( n26152 ) & (n26153 )  ;
assign n26155 =  ( n26154 ) & (wr )  ;
assign n26156 =  ( n26155 ) ? ( n5485 ) : ( iram_220 ) ;
assign n26157 = wr_addr[7:7] ;
assign n26158 =  ( n26157 ) == ( bv_1_0_n53 )  ;
assign n26159 =  ( wr_addr ) == ( bv_8_220_n509 )  ;
assign n26160 =  ( n26158 ) & (n26159 )  ;
assign n26161 =  ( n26160 ) & (wr )  ;
assign n26162 =  ( n26161 ) ? ( n5512 ) : ( iram_220 ) ;
assign n26163 = wr_addr[7:7] ;
assign n26164 =  ( n26163 ) == ( bv_1_0_n53 )  ;
assign n26165 =  ( wr_addr ) == ( bv_8_220_n509 )  ;
assign n26166 =  ( n26164 ) & (n26165 )  ;
assign n26167 =  ( n26166 ) & (wr )  ;
assign n26168 =  ( n26167 ) ? ( bv_8_0_n69 ) : ( iram_220 ) ;
assign n26169 = wr_addr[7:7] ;
assign n26170 =  ( n26169 ) == ( bv_1_0_n53 )  ;
assign n26171 =  ( wr_addr ) == ( bv_8_220_n509 )  ;
assign n26172 =  ( n26170 ) & (n26171 )  ;
assign n26173 =  ( n26172 ) & (wr )  ;
assign n26174 =  ( n26173 ) ? ( n5071 ) : ( iram_220 ) ;
assign n26175 = wr_addr[7:7] ;
assign n26176 =  ( n26175 ) == ( bv_1_0_n53 )  ;
assign n26177 =  ( wr_addr ) == ( bv_8_220_n509 )  ;
assign n26178 =  ( n26176 ) & (n26177 )  ;
assign n26179 =  ( n26178 ) & (wr )  ;
assign n26180 =  ( n26179 ) ? ( n5096 ) : ( iram_220 ) ;
assign n26181 = wr_addr[7:7] ;
assign n26182 =  ( n26181 ) == ( bv_1_0_n53 )  ;
assign n26183 =  ( wr_addr ) == ( bv_8_220_n509 )  ;
assign n26184 =  ( n26182 ) & (n26183 )  ;
assign n26185 =  ( n26184 ) & (wr )  ;
assign n26186 =  ( n26185 ) ? ( n5123 ) : ( iram_220 ) ;
assign n26187 = wr_addr[7:7] ;
assign n26188 =  ( n26187 ) == ( bv_1_0_n53 )  ;
assign n26189 =  ( wr_addr ) == ( bv_8_220_n509 )  ;
assign n26190 =  ( n26188 ) & (n26189 )  ;
assign n26191 =  ( n26190 ) & (wr )  ;
assign n26192 =  ( n26191 ) ? ( n5165 ) : ( iram_220 ) ;
assign n26193 = wr_addr[7:7] ;
assign n26194 =  ( n26193 ) == ( bv_1_0_n53 )  ;
assign n26195 =  ( wr_addr ) == ( bv_8_220_n509 )  ;
assign n26196 =  ( n26194 ) & (n26195 )  ;
assign n26197 =  ( n26196 ) & (wr )  ;
assign n26198 =  ( n26197 ) ? ( n5204 ) : ( iram_220 ) ;
assign n26199 = wr_addr[7:7] ;
assign n26200 =  ( n26199 ) == ( bv_1_0_n53 )  ;
assign n26201 =  ( wr_addr ) == ( bv_8_220_n509 )  ;
assign n26202 =  ( n26200 ) & (n26201 )  ;
assign n26203 =  ( n26202 ) & (wr )  ;
assign n26204 =  ( n26203 ) ? ( n5262 ) : ( iram_220 ) ;
assign n26205 = wr_addr[7:7] ;
assign n26206 =  ( n26205 ) == ( bv_1_0_n53 )  ;
assign n26207 =  ( wr_addr ) == ( bv_8_220_n509 )  ;
assign n26208 =  ( n26206 ) & (n26207 )  ;
assign n26209 =  ( n26208 ) & (wr )  ;
assign n26210 =  ( n26209 ) ? ( n5298 ) : ( iram_220 ) ;
assign n26211 = wr_addr[7:7] ;
assign n26212 =  ( n26211 ) == ( bv_1_0_n53 )  ;
assign n26213 =  ( wr_addr ) == ( bv_8_220_n509 )  ;
assign n26214 =  ( n26212 ) & (n26213 )  ;
assign n26215 =  ( n26214 ) & (wr )  ;
assign n26216 =  ( n26215 ) ? ( n5325 ) : ( iram_220 ) ;
assign n26217 = wr_addr[7:7] ;
assign n26218 =  ( n26217 ) == ( bv_1_0_n53 )  ;
assign n26219 =  ( wr_addr ) == ( bv_8_221_n511 )  ;
assign n26220 =  ( n26218 ) & (n26219 )  ;
assign n26221 =  ( n26220 ) & (wr )  ;
assign n26222 =  ( n26221 ) ? ( n4782 ) : ( iram_221 ) ;
assign n26223 = wr_addr[7:7] ;
assign n26224 =  ( n26223 ) == ( bv_1_0_n53 )  ;
assign n26225 =  ( wr_addr ) == ( bv_8_221_n511 )  ;
assign n26226 =  ( n26224 ) & (n26225 )  ;
assign n26227 =  ( n26226 ) & (wr )  ;
assign n26228 =  ( n26227 ) ? ( n4841 ) : ( iram_221 ) ;
assign n26229 = wr_addr[7:7] ;
assign n26230 =  ( n26229 ) == ( bv_1_0_n53 )  ;
assign n26231 =  ( wr_addr ) == ( bv_8_221_n511 )  ;
assign n26232 =  ( n26230 ) & (n26231 )  ;
assign n26233 =  ( n26232 ) & (wr )  ;
assign n26234 =  ( n26233 ) ? ( n5449 ) : ( iram_221 ) ;
assign n26235 = wr_addr[7:7] ;
assign n26236 =  ( n26235 ) == ( bv_1_0_n53 )  ;
assign n26237 =  ( wr_addr ) == ( bv_8_221_n511 )  ;
assign n26238 =  ( n26236 ) & (n26237 )  ;
assign n26239 =  ( n26238 ) & (wr )  ;
assign n26240 =  ( n26239 ) ? ( n4906 ) : ( iram_221 ) ;
assign n26241 = wr_addr[7:7] ;
assign n26242 =  ( n26241 ) == ( bv_1_0_n53 )  ;
assign n26243 =  ( wr_addr ) == ( bv_8_221_n511 )  ;
assign n26244 =  ( n26242 ) & (n26243 )  ;
assign n26245 =  ( n26244 ) & (wr )  ;
assign n26246 =  ( n26245 ) ? ( n5485 ) : ( iram_221 ) ;
assign n26247 = wr_addr[7:7] ;
assign n26248 =  ( n26247 ) == ( bv_1_0_n53 )  ;
assign n26249 =  ( wr_addr ) == ( bv_8_221_n511 )  ;
assign n26250 =  ( n26248 ) & (n26249 )  ;
assign n26251 =  ( n26250 ) & (wr )  ;
assign n26252 =  ( n26251 ) ? ( n5512 ) : ( iram_221 ) ;
assign n26253 = wr_addr[7:7] ;
assign n26254 =  ( n26253 ) == ( bv_1_0_n53 )  ;
assign n26255 =  ( wr_addr ) == ( bv_8_221_n511 )  ;
assign n26256 =  ( n26254 ) & (n26255 )  ;
assign n26257 =  ( n26256 ) & (wr )  ;
assign n26258 =  ( n26257 ) ? ( bv_8_0_n69 ) : ( iram_221 ) ;
assign n26259 = wr_addr[7:7] ;
assign n26260 =  ( n26259 ) == ( bv_1_0_n53 )  ;
assign n26261 =  ( wr_addr ) == ( bv_8_221_n511 )  ;
assign n26262 =  ( n26260 ) & (n26261 )  ;
assign n26263 =  ( n26262 ) & (wr )  ;
assign n26264 =  ( n26263 ) ? ( n5071 ) : ( iram_221 ) ;
assign n26265 = wr_addr[7:7] ;
assign n26266 =  ( n26265 ) == ( bv_1_0_n53 )  ;
assign n26267 =  ( wr_addr ) == ( bv_8_221_n511 )  ;
assign n26268 =  ( n26266 ) & (n26267 )  ;
assign n26269 =  ( n26268 ) & (wr )  ;
assign n26270 =  ( n26269 ) ? ( n5096 ) : ( iram_221 ) ;
assign n26271 = wr_addr[7:7] ;
assign n26272 =  ( n26271 ) == ( bv_1_0_n53 )  ;
assign n26273 =  ( wr_addr ) == ( bv_8_221_n511 )  ;
assign n26274 =  ( n26272 ) & (n26273 )  ;
assign n26275 =  ( n26274 ) & (wr )  ;
assign n26276 =  ( n26275 ) ? ( n5123 ) : ( iram_221 ) ;
assign n26277 = wr_addr[7:7] ;
assign n26278 =  ( n26277 ) == ( bv_1_0_n53 )  ;
assign n26279 =  ( wr_addr ) == ( bv_8_221_n511 )  ;
assign n26280 =  ( n26278 ) & (n26279 )  ;
assign n26281 =  ( n26280 ) & (wr )  ;
assign n26282 =  ( n26281 ) ? ( n5165 ) : ( iram_221 ) ;
assign n26283 = wr_addr[7:7] ;
assign n26284 =  ( n26283 ) == ( bv_1_0_n53 )  ;
assign n26285 =  ( wr_addr ) == ( bv_8_221_n511 )  ;
assign n26286 =  ( n26284 ) & (n26285 )  ;
assign n26287 =  ( n26286 ) & (wr )  ;
assign n26288 =  ( n26287 ) ? ( n5204 ) : ( iram_221 ) ;
assign n26289 = wr_addr[7:7] ;
assign n26290 =  ( n26289 ) == ( bv_1_0_n53 )  ;
assign n26291 =  ( wr_addr ) == ( bv_8_221_n511 )  ;
assign n26292 =  ( n26290 ) & (n26291 )  ;
assign n26293 =  ( n26292 ) & (wr )  ;
assign n26294 =  ( n26293 ) ? ( n5262 ) : ( iram_221 ) ;
assign n26295 = wr_addr[7:7] ;
assign n26296 =  ( n26295 ) == ( bv_1_0_n53 )  ;
assign n26297 =  ( wr_addr ) == ( bv_8_221_n511 )  ;
assign n26298 =  ( n26296 ) & (n26297 )  ;
assign n26299 =  ( n26298 ) & (wr )  ;
assign n26300 =  ( n26299 ) ? ( n5298 ) : ( iram_221 ) ;
assign n26301 = wr_addr[7:7] ;
assign n26302 =  ( n26301 ) == ( bv_1_0_n53 )  ;
assign n26303 =  ( wr_addr ) == ( bv_8_221_n511 )  ;
assign n26304 =  ( n26302 ) & (n26303 )  ;
assign n26305 =  ( n26304 ) & (wr )  ;
assign n26306 =  ( n26305 ) ? ( n5325 ) : ( iram_221 ) ;
assign n26307 = wr_addr[7:7] ;
assign n26308 =  ( n26307 ) == ( bv_1_0_n53 )  ;
assign n26309 =  ( wr_addr ) == ( bv_8_222_n513 )  ;
assign n26310 =  ( n26308 ) & (n26309 )  ;
assign n26311 =  ( n26310 ) & (wr )  ;
assign n26312 =  ( n26311 ) ? ( n4782 ) : ( iram_222 ) ;
assign n26313 = wr_addr[7:7] ;
assign n26314 =  ( n26313 ) == ( bv_1_0_n53 )  ;
assign n26315 =  ( wr_addr ) == ( bv_8_222_n513 )  ;
assign n26316 =  ( n26314 ) & (n26315 )  ;
assign n26317 =  ( n26316 ) & (wr )  ;
assign n26318 =  ( n26317 ) ? ( n4841 ) : ( iram_222 ) ;
assign n26319 = wr_addr[7:7] ;
assign n26320 =  ( n26319 ) == ( bv_1_0_n53 )  ;
assign n26321 =  ( wr_addr ) == ( bv_8_222_n513 )  ;
assign n26322 =  ( n26320 ) & (n26321 )  ;
assign n26323 =  ( n26322 ) & (wr )  ;
assign n26324 =  ( n26323 ) ? ( n5449 ) : ( iram_222 ) ;
assign n26325 = wr_addr[7:7] ;
assign n26326 =  ( n26325 ) == ( bv_1_0_n53 )  ;
assign n26327 =  ( wr_addr ) == ( bv_8_222_n513 )  ;
assign n26328 =  ( n26326 ) & (n26327 )  ;
assign n26329 =  ( n26328 ) & (wr )  ;
assign n26330 =  ( n26329 ) ? ( n4906 ) : ( iram_222 ) ;
assign n26331 = wr_addr[7:7] ;
assign n26332 =  ( n26331 ) == ( bv_1_0_n53 )  ;
assign n26333 =  ( wr_addr ) == ( bv_8_222_n513 )  ;
assign n26334 =  ( n26332 ) & (n26333 )  ;
assign n26335 =  ( n26334 ) & (wr )  ;
assign n26336 =  ( n26335 ) ? ( n5485 ) : ( iram_222 ) ;
assign n26337 = wr_addr[7:7] ;
assign n26338 =  ( n26337 ) == ( bv_1_0_n53 )  ;
assign n26339 =  ( wr_addr ) == ( bv_8_222_n513 )  ;
assign n26340 =  ( n26338 ) & (n26339 )  ;
assign n26341 =  ( n26340 ) & (wr )  ;
assign n26342 =  ( n26341 ) ? ( n5512 ) : ( iram_222 ) ;
assign n26343 = wr_addr[7:7] ;
assign n26344 =  ( n26343 ) == ( bv_1_0_n53 )  ;
assign n26345 =  ( wr_addr ) == ( bv_8_222_n513 )  ;
assign n26346 =  ( n26344 ) & (n26345 )  ;
assign n26347 =  ( n26346 ) & (wr )  ;
assign n26348 =  ( n26347 ) ? ( bv_8_0_n69 ) : ( iram_222 ) ;
assign n26349 = wr_addr[7:7] ;
assign n26350 =  ( n26349 ) == ( bv_1_0_n53 )  ;
assign n26351 =  ( wr_addr ) == ( bv_8_222_n513 )  ;
assign n26352 =  ( n26350 ) & (n26351 )  ;
assign n26353 =  ( n26352 ) & (wr )  ;
assign n26354 =  ( n26353 ) ? ( n5071 ) : ( iram_222 ) ;
assign n26355 = wr_addr[7:7] ;
assign n26356 =  ( n26355 ) == ( bv_1_0_n53 )  ;
assign n26357 =  ( wr_addr ) == ( bv_8_222_n513 )  ;
assign n26358 =  ( n26356 ) & (n26357 )  ;
assign n26359 =  ( n26358 ) & (wr )  ;
assign n26360 =  ( n26359 ) ? ( n5096 ) : ( iram_222 ) ;
assign n26361 = wr_addr[7:7] ;
assign n26362 =  ( n26361 ) == ( bv_1_0_n53 )  ;
assign n26363 =  ( wr_addr ) == ( bv_8_222_n513 )  ;
assign n26364 =  ( n26362 ) & (n26363 )  ;
assign n26365 =  ( n26364 ) & (wr )  ;
assign n26366 =  ( n26365 ) ? ( n5123 ) : ( iram_222 ) ;
assign n26367 = wr_addr[7:7] ;
assign n26368 =  ( n26367 ) == ( bv_1_0_n53 )  ;
assign n26369 =  ( wr_addr ) == ( bv_8_222_n513 )  ;
assign n26370 =  ( n26368 ) & (n26369 )  ;
assign n26371 =  ( n26370 ) & (wr )  ;
assign n26372 =  ( n26371 ) ? ( n5165 ) : ( iram_222 ) ;
assign n26373 = wr_addr[7:7] ;
assign n26374 =  ( n26373 ) == ( bv_1_0_n53 )  ;
assign n26375 =  ( wr_addr ) == ( bv_8_222_n513 )  ;
assign n26376 =  ( n26374 ) & (n26375 )  ;
assign n26377 =  ( n26376 ) & (wr )  ;
assign n26378 =  ( n26377 ) ? ( n5204 ) : ( iram_222 ) ;
assign n26379 = wr_addr[7:7] ;
assign n26380 =  ( n26379 ) == ( bv_1_0_n53 )  ;
assign n26381 =  ( wr_addr ) == ( bv_8_222_n513 )  ;
assign n26382 =  ( n26380 ) & (n26381 )  ;
assign n26383 =  ( n26382 ) & (wr )  ;
assign n26384 =  ( n26383 ) ? ( n5262 ) : ( iram_222 ) ;
assign n26385 = wr_addr[7:7] ;
assign n26386 =  ( n26385 ) == ( bv_1_0_n53 )  ;
assign n26387 =  ( wr_addr ) == ( bv_8_222_n513 )  ;
assign n26388 =  ( n26386 ) & (n26387 )  ;
assign n26389 =  ( n26388 ) & (wr )  ;
assign n26390 =  ( n26389 ) ? ( n5298 ) : ( iram_222 ) ;
assign n26391 = wr_addr[7:7] ;
assign n26392 =  ( n26391 ) == ( bv_1_0_n53 )  ;
assign n26393 =  ( wr_addr ) == ( bv_8_222_n513 )  ;
assign n26394 =  ( n26392 ) & (n26393 )  ;
assign n26395 =  ( n26394 ) & (wr )  ;
assign n26396 =  ( n26395 ) ? ( n5325 ) : ( iram_222 ) ;
assign n26397 = wr_addr[7:7] ;
assign n26398 =  ( n26397 ) == ( bv_1_0_n53 )  ;
assign n26399 =  ( wr_addr ) == ( bv_8_223_n515 )  ;
assign n26400 =  ( n26398 ) & (n26399 )  ;
assign n26401 =  ( n26400 ) & (wr )  ;
assign n26402 =  ( n26401 ) ? ( n4782 ) : ( iram_223 ) ;
assign n26403 = wr_addr[7:7] ;
assign n26404 =  ( n26403 ) == ( bv_1_0_n53 )  ;
assign n26405 =  ( wr_addr ) == ( bv_8_223_n515 )  ;
assign n26406 =  ( n26404 ) & (n26405 )  ;
assign n26407 =  ( n26406 ) & (wr )  ;
assign n26408 =  ( n26407 ) ? ( n4841 ) : ( iram_223 ) ;
assign n26409 = wr_addr[7:7] ;
assign n26410 =  ( n26409 ) == ( bv_1_0_n53 )  ;
assign n26411 =  ( wr_addr ) == ( bv_8_223_n515 )  ;
assign n26412 =  ( n26410 ) & (n26411 )  ;
assign n26413 =  ( n26412 ) & (wr )  ;
assign n26414 =  ( n26413 ) ? ( n5449 ) : ( iram_223 ) ;
assign n26415 = wr_addr[7:7] ;
assign n26416 =  ( n26415 ) == ( bv_1_0_n53 )  ;
assign n26417 =  ( wr_addr ) == ( bv_8_223_n515 )  ;
assign n26418 =  ( n26416 ) & (n26417 )  ;
assign n26419 =  ( n26418 ) & (wr )  ;
assign n26420 =  ( n26419 ) ? ( n4906 ) : ( iram_223 ) ;
assign n26421 = wr_addr[7:7] ;
assign n26422 =  ( n26421 ) == ( bv_1_0_n53 )  ;
assign n26423 =  ( wr_addr ) == ( bv_8_223_n515 )  ;
assign n26424 =  ( n26422 ) & (n26423 )  ;
assign n26425 =  ( n26424 ) & (wr )  ;
assign n26426 =  ( n26425 ) ? ( n5485 ) : ( iram_223 ) ;
assign n26427 = wr_addr[7:7] ;
assign n26428 =  ( n26427 ) == ( bv_1_0_n53 )  ;
assign n26429 =  ( wr_addr ) == ( bv_8_223_n515 )  ;
assign n26430 =  ( n26428 ) & (n26429 )  ;
assign n26431 =  ( n26430 ) & (wr )  ;
assign n26432 =  ( n26431 ) ? ( n5512 ) : ( iram_223 ) ;
assign n26433 = wr_addr[7:7] ;
assign n26434 =  ( n26433 ) == ( bv_1_0_n53 )  ;
assign n26435 =  ( wr_addr ) == ( bv_8_223_n515 )  ;
assign n26436 =  ( n26434 ) & (n26435 )  ;
assign n26437 =  ( n26436 ) & (wr )  ;
assign n26438 =  ( n26437 ) ? ( bv_8_0_n69 ) : ( iram_223 ) ;
assign n26439 = wr_addr[7:7] ;
assign n26440 =  ( n26439 ) == ( bv_1_0_n53 )  ;
assign n26441 =  ( wr_addr ) == ( bv_8_223_n515 )  ;
assign n26442 =  ( n26440 ) & (n26441 )  ;
assign n26443 =  ( n26442 ) & (wr )  ;
assign n26444 =  ( n26443 ) ? ( n5071 ) : ( iram_223 ) ;
assign n26445 = wr_addr[7:7] ;
assign n26446 =  ( n26445 ) == ( bv_1_0_n53 )  ;
assign n26447 =  ( wr_addr ) == ( bv_8_223_n515 )  ;
assign n26448 =  ( n26446 ) & (n26447 )  ;
assign n26449 =  ( n26448 ) & (wr )  ;
assign n26450 =  ( n26449 ) ? ( n5096 ) : ( iram_223 ) ;
assign n26451 = wr_addr[7:7] ;
assign n26452 =  ( n26451 ) == ( bv_1_0_n53 )  ;
assign n26453 =  ( wr_addr ) == ( bv_8_223_n515 )  ;
assign n26454 =  ( n26452 ) & (n26453 )  ;
assign n26455 =  ( n26454 ) & (wr )  ;
assign n26456 =  ( n26455 ) ? ( n5123 ) : ( iram_223 ) ;
assign n26457 = wr_addr[7:7] ;
assign n26458 =  ( n26457 ) == ( bv_1_0_n53 )  ;
assign n26459 =  ( wr_addr ) == ( bv_8_223_n515 )  ;
assign n26460 =  ( n26458 ) & (n26459 )  ;
assign n26461 =  ( n26460 ) & (wr )  ;
assign n26462 =  ( n26461 ) ? ( n5165 ) : ( iram_223 ) ;
assign n26463 = wr_addr[7:7] ;
assign n26464 =  ( n26463 ) == ( bv_1_0_n53 )  ;
assign n26465 =  ( wr_addr ) == ( bv_8_223_n515 )  ;
assign n26466 =  ( n26464 ) & (n26465 )  ;
assign n26467 =  ( n26466 ) & (wr )  ;
assign n26468 =  ( n26467 ) ? ( n5204 ) : ( iram_223 ) ;
assign n26469 = wr_addr[7:7] ;
assign n26470 =  ( n26469 ) == ( bv_1_0_n53 )  ;
assign n26471 =  ( wr_addr ) == ( bv_8_223_n515 )  ;
assign n26472 =  ( n26470 ) & (n26471 )  ;
assign n26473 =  ( n26472 ) & (wr )  ;
assign n26474 =  ( n26473 ) ? ( n5262 ) : ( iram_223 ) ;
assign n26475 = wr_addr[7:7] ;
assign n26476 =  ( n26475 ) == ( bv_1_0_n53 )  ;
assign n26477 =  ( wr_addr ) == ( bv_8_223_n515 )  ;
assign n26478 =  ( n26476 ) & (n26477 )  ;
assign n26479 =  ( n26478 ) & (wr )  ;
assign n26480 =  ( n26479 ) ? ( n5298 ) : ( iram_223 ) ;
assign n26481 = wr_addr[7:7] ;
assign n26482 =  ( n26481 ) == ( bv_1_0_n53 )  ;
assign n26483 =  ( wr_addr ) == ( bv_8_223_n515 )  ;
assign n26484 =  ( n26482 ) & (n26483 )  ;
assign n26485 =  ( n26484 ) & (wr )  ;
assign n26486 =  ( n26485 ) ? ( n5325 ) : ( iram_223 ) ;
assign n26487 = wr_addr[7:7] ;
assign n26488 =  ( n26487 ) == ( bv_1_0_n53 )  ;
assign n26489 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n26490 =  ( n26488 ) & (n26489 )  ;
assign n26491 =  ( n26490 ) & (wr )  ;
assign n26492 =  ( n26491 ) ? ( n4782 ) : ( iram_224 ) ;
assign n26493 = wr_addr[7:7] ;
assign n26494 =  ( n26493 ) == ( bv_1_0_n53 )  ;
assign n26495 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n26496 =  ( n26494 ) & (n26495 )  ;
assign n26497 =  ( n26496 ) & (wr )  ;
assign n26498 =  ( n26497 ) ? ( n4841 ) : ( iram_224 ) ;
assign n26499 = wr_addr[7:7] ;
assign n26500 =  ( n26499 ) == ( bv_1_0_n53 )  ;
assign n26501 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n26502 =  ( n26500 ) & (n26501 )  ;
assign n26503 =  ( n26502 ) & (wr )  ;
assign n26504 =  ( n26503 ) ? ( n5449 ) : ( iram_224 ) ;
assign n26505 = wr_addr[7:7] ;
assign n26506 =  ( n26505 ) == ( bv_1_0_n53 )  ;
assign n26507 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n26508 =  ( n26506 ) & (n26507 )  ;
assign n26509 =  ( n26508 ) & (wr )  ;
assign n26510 =  ( n26509 ) ? ( n4906 ) : ( iram_224 ) ;
assign n26511 = wr_addr[7:7] ;
assign n26512 =  ( n26511 ) == ( bv_1_0_n53 )  ;
assign n26513 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n26514 =  ( n26512 ) & (n26513 )  ;
assign n26515 =  ( n26514 ) & (wr )  ;
assign n26516 =  ( n26515 ) ? ( n5485 ) : ( iram_224 ) ;
assign n26517 = wr_addr[7:7] ;
assign n26518 =  ( n26517 ) == ( bv_1_0_n53 )  ;
assign n26519 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n26520 =  ( n26518 ) & (n26519 )  ;
assign n26521 =  ( n26520 ) & (wr )  ;
assign n26522 =  ( n26521 ) ? ( n5512 ) : ( iram_224 ) ;
assign n26523 = wr_addr[7:7] ;
assign n26524 =  ( n26523 ) == ( bv_1_0_n53 )  ;
assign n26525 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n26526 =  ( n26524 ) & (n26525 )  ;
assign n26527 =  ( n26526 ) & (wr )  ;
assign n26528 =  ( n26527 ) ? ( bv_8_0_n69 ) : ( iram_224 ) ;
assign n26529 = wr_addr[7:7] ;
assign n26530 =  ( n26529 ) == ( bv_1_0_n53 )  ;
assign n26531 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n26532 =  ( n26530 ) & (n26531 )  ;
assign n26533 =  ( n26532 ) & (wr )  ;
assign n26534 =  ( n26533 ) ? ( n5071 ) : ( iram_224 ) ;
assign n26535 = wr_addr[7:7] ;
assign n26536 =  ( n26535 ) == ( bv_1_0_n53 )  ;
assign n26537 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n26538 =  ( n26536 ) & (n26537 )  ;
assign n26539 =  ( n26538 ) & (wr )  ;
assign n26540 =  ( n26539 ) ? ( n5096 ) : ( iram_224 ) ;
assign n26541 = wr_addr[7:7] ;
assign n26542 =  ( n26541 ) == ( bv_1_0_n53 )  ;
assign n26543 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n26544 =  ( n26542 ) & (n26543 )  ;
assign n26545 =  ( n26544 ) & (wr )  ;
assign n26546 =  ( n26545 ) ? ( n5123 ) : ( iram_224 ) ;
assign n26547 = wr_addr[7:7] ;
assign n26548 =  ( n26547 ) == ( bv_1_0_n53 )  ;
assign n26549 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n26550 =  ( n26548 ) & (n26549 )  ;
assign n26551 =  ( n26550 ) & (wr )  ;
assign n26552 =  ( n26551 ) ? ( n5165 ) : ( iram_224 ) ;
assign n26553 = wr_addr[7:7] ;
assign n26554 =  ( n26553 ) == ( bv_1_0_n53 )  ;
assign n26555 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n26556 =  ( n26554 ) & (n26555 )  ;
assign n26557 =  ( n26556 ) & (wr )  ;
assign n26558 =  ( n26557 ) ? ( n5204 ) : ( iram_224 ) ;
assign n26559 = wr_addr[7:7] ;
assign n26560 =  ( n26559 ) == ( bv_1_0_n53 )  ;
assign n26561 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n26562 =  ( n26560 ) & (n26561 )  ;
assign n26563 =  ( n26562 ) & (wr )  ;
assign n26564 =  ( n26563 ) ? ( n5262 ) : ( iram_224 ) ;
assign n26565 = wr_addr[7:7] ;
assign n26566 =  ( n26565 ) == ( bv_1_0_n53 )  ;
assign n26567 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n26568 =  ( n26566 ) & (n26567 )  ;
assign n26569 =  ( n26568 ) & (wr )  ;
assign n26570 =  ( n26569 ) ? ( n5298 ) : ( iram_224 ) ;
assign n26571 = wr_addr[7:7] ;
assign n26572 =  ( n26571 ) == ( bv_1_0_n53 )  ;
assign n26573 =  ( wr_addr ) == ( bv_8_224_n517 )  ;
assign n26574 =  ( n26572 ) & (n26573 )  ;
assign n26575 =  ( n26574 ) & (wr )  ;
assign n26576 =  ( n26575 ) ? ( n5325 ) : ( iram_224 ) ;
assign n26577 = wr_addr[7:7] ;
assign n26578 =  ( n26577 ) == ( bv_1_0_n53 )  ;
assign n26579 =  ( wr_addr ) == ( bv_8_225_n519 )  ;
assign n26580 =  ( n26578 ) & (n26579 )  ;
assign n26581 =  ( n26580 ) & (wr )  ;
assign n26582 =  ( n26581 ) ? ( n4782 ) : ( iram_225 ) ;
assign n26583 = wr_addr[7:7] ;
assign n26584 =  ( n26583 ) == ( bv_1_0_n53 )  ;
assign n26585 =  ( wr_addr ) == ( bv_8_225_n519 )  ;
assign n26586 =  ( n26584 ) & (n26585 )  ;
assign n26587 =  ( n26586 ) & (wr )  ;
assign n26588 =  ( n26587 ) ? ( n4841 ) : ( iram_225 ) ;
assign n26589 = wr_addr[7:7] ;
assign n26590 =  ( n26589 ) == ( bv_1_0_n53 )  ;
assign n26591 =  ( wr_addr ) == ( bv_8_225_n519 )  ;
assign n26592 =  ( n26590 ) & (n26591 )  ;
assign n26593 =  ( n26592 ) & (wr )  ;
assign n26594 =  ( n26593 ) ? ( n5449 ) : ( iram_225 ) ;
assign n26595 = wr_addr[7:7] ;
assign n26596 =  ( n26595 ) == ( bv_1_0_n53 )  ;
assign n26597 =  ( wr_addr ) == ( bv_8_225_n519 )  ;
assign n26598 =  ( n26596 ) & (n26597 )  ;
assign n26599 =  ( n26598 ) & (wr )  ;
assign n26600 =  ( n26599 ) ? ( n4906 ) : ( iram_225 ) ;
assign n26601 = wr_addr[7:7] ;
assign n26602 =  ( n26601 ) == ( bv_1_0_n53 )  ;
assign n26603 =  ( wr_addr ) == ( bv_8_225_n519 )  ;
assign n26604 =  ( n26602 ) & (n26603 )  ;
assign n26605 =  ( n26604 ) & (wr )  ;
assign n26606 =  ( n26605 ) ? ( n5485 ) : ( iram_225 ) ;
assign n26607 = wr_addr[7:7] ;
assign n26608 =  ( n26607 ) == ( bv_1_0_n53 )  ;
assign n26609 =  ( wr_addr ) == ( bv_8_225_n519 )  ;
assign n26610 =  ( n26608 ) & (n26609 )  ;
assign n26611 =  ( n26610 ) & (wr )  ;
assign n26612 =  ( n26611 ) ? ( n5512 ) : ( iram_225 ) ;
assign n26613 = wr_addr[7:7] ;
assign n26614 =  ( n26613 ) == ( bv_1_0_n53 )  ;
assign n26615 =  ( wr_addr ) == ( bv_8_225_n519 )  ;
assign n26616 =  ( n26614 ) & (n26615 )  ;
assign n26617 =  ( n26616 ) & (wr )  ;
assign n26618 =  ( n26617 ) ? ( bv_8_0_n69 ) : ( iram_225 ) ;
assign n26619 = wr_addr[7:7] ;
assign n26620 =  ( n26619 ) == ( bv_1_0_n53 )  ;
assign n26621 =  ( wr_addr ) == ( bv_8_225_n519 )  ;
assign n26622 =  ( n26620 ) & (n26621 )  ;
assign n26623 =  ( n26622 ) & (wr )  ;
assign n26624 =  ( n26623 ) ? ( n5071 ) : ( iram_225 ) ;
assign n26625 = wr_addr[7:7] ;
assign n26626 =  ( n26625 ) == ( bv_1_0_n53 )  ;
assign n26627 =  ( wr_addr ) == ( bv_8_225_n519 )  ;
assign n26628 =  ( n26626 ) & (n26627 )  ;
assign n26629 =  ( n26628 ) & (wr )  ;
assign n26630 =  ( n26629 ) ? ( n5096 ) : ( iram_225 ) ;
assign n26631 = wr_addr[7:7] ;
assign n26632 =  ( n26631 ) == ( bv_1_0_n53 )  ;
assign n26633 =  ( wr_addr ) == ( bv_8_225_n519 )  ;
assign n26634 =  ( n26632 ) & (n26633 )  ;
assign n26635 =  ( n26634 ) & (wr )  ;
assign n26636 =  ( n26635 ) ? ( n5123 ) : ( iram_225 ) ;
assign n26637 = wr_addr[7:7] ;
assign n26638 =  ( n26637 ) == ( bv_1_0_n53 )  ;
assign n26639 =  ( wr_addr ) == ( bv_8_225_n519 )  ;
assign n26640 =  ( n26638 ) & (n26639 )  ;
assign n26641 =  ( n26640 ) & (wr )  ;
assign n26642 =  ( n26641 ) ? ( n5165 ) : ( iram_225 ) ;
assign n26643 = wr_addr[7:7] ;
assign n26644 =  ( n26643 ) == ( bv_1_0_n53 )  ;
assign n26645 =  ( wr_addr ) == ( bv_8_225_n519 )  ;
assign n26646 =  ( n26644 ) & (n26645 )  ;
assign n26647 =  ( n26646 ) & (wr )  ;
assign n26648 =  ( n26647 ) ? ( n5204 ) : ( iram_225 ) ;
assign n26649 = wr_addr[7:7] ;
assign n26650 =  ( n26649 ) == ( bv_1_0_n53 )  ;
assign n26651 =  ( wr_addr ) == ( bv_8_225_n519 )  ;
assign n26652 =  ( n26650 ) & (n26651 )  ;
assign n26653 =  ( n26652 ) & (wr )  ;
assign n26654 =  ( n26653 ) ? ( n5262 ) : ( iram_225 ) ;
assign n26655 = wr_addr[7:7] ;
assign n26656 =  ( n26655 ) == ( bv_1_0_n53 )  ;
assign n26657 =  ( wr_addr ) == ( bv_8_225_n519 )  ;
assign n26658 =  ( n26656 ) & (n26657 )  ;
assign n26659 =  ( n26658 ) & (wr )  ;
assign n26660 =  ( n26659 ) ? ( n5298 ) : ( iram_225 ) ;
assign n26661 = wr_addr[7:7] ;
assign n26662 =  ( n26661 ) == ( bv_1_0_n53 )  ;
assign n26663 =  ( wr_addr ) == ( bv_8_225_n519 )  ;
assign n26664 =  ( n26662 ) & (n26663 )  ;
assign n26665 =  ( n26664 ) & (wr )  ;
assign n26666 =  ( n26665 ) ? ( n5325 ) : ( iram_225 ) ;
assign n26667 = wr_addr[7:7] ;
assign n26668 =  ( n26667 ) == ( bv_1_0_n53 )  ;
assign n26669 =  ( wr_addr ) == ( bv_8_226_n521 )  ;
assign n26670 =  ( n26668 ) & (n26669 )  ;
assign n26671 =  ( n26670 ) & (wr )  ;
assign n26672 =  ( n26671 ) ? ( n4782 ) : ( iram_226 ) ;
assign n26673 = wr_addr[7:7] ;
assign n26674 =  ( n26673 ) == ( bv_1_0_n53 )  ;
assign n26675 =  ( wr_addr ) == ( bv_8_226_n521 )  ;
assign n26676 =  ( n26674 ) & (n26675 )  ;
assign n26677 =  ( n26676 ) & (wr )  ;
assign n26678 =  ( n26677 ) ? ( n4841 ) : ( iram_226 ) ;
assign n26679 = wr_addr[7:7] ;
assign n26680 =  ( n26679 ) == ( bv_1_0_n53 )  ;
assign n26681 =  ( wr_addr ) == ( bv_8_226_n521 )  ;
assign n26682 =  ( n26680 ) & (n26681 )  ;
assign n26683 =  ( n26682 ) & (wr )  ;
assign n26684 =  ( n26683 ) ? ( n5449 ) : ( iram_226 ) ;
assign n26685 = wr_addr[7:7] ;
assign n26686 =  ( n26685 ) == ( bv_1_0_n53 )  ;
assign n26687 =  ( wr_addr ) == ( bv_8_226_n521 )  ;
assign n26688 =  ( n26686 ) & (n26687 )  ;
assign n26689 =  ( n26688 ) & (wr )  ;
assign n26690 =  ( n26689 ) ? ( n4906 ) : ( iram_226 ) ;
assign n26691 = wr_addr[7:7] ;
assign n26692 =  ( n26691 ) == ( bv_1_0_n53 )  ;
assign n26693 =  ( wr_addr ) == ( bv_8_226_n521 )  ;
assign n26694 =  ( n26692 ) & (n26693 )  ;
assign n26695 =  ( n26694 ) & (wr )  ;
assign n26696 =  ( n26695 ) ? ( n5485 ) : ( iram_226 ) ;
assign n26697 = wr_addr[7:7] ;
assign n26698 =  ( n26697 ) == ( bv_1_0_n53 )  ;
assign n26699 =  ( wr_addr ) == ( bv_8_226_n521 )  ;
assign n26700 =  ( n26698 ) & (n26699 )  ;
assign n26701 =  ( n26700 ) & (wr )  ;
assign n26702 =  ( n26701 ) ? ( n5512 ) : ( iram_226 ) ;
assign n26703 = wr_addr[7:7] ;
assign n26704 =  ( n26703 ) == ( bv_1_0_n53 )  ;
assign n26705 =  ( wr_addr ) == ( bv_8_226_n521 )  ;
assign n26706 =  ( n26704 ) & (n26705 )  ;
assign n26707 =  ( n26706 ) & (wr )  ;
assign n26708 =  ( n26707 ) ? ( bv_8_0_n69 ) : ( iram_226 ) ;
assign n26709 = wr_addr[7:7] ;
assign n26710 =  ( n26709 ) == ( bv_1_0_n53 )  ;
assign n26711 =  ( wr_addr ) == ( bv_8_226_n521 )  ;
assign n26712 =  ( n26710 ) & (n26711 )  ;
assign n26713 =  ( n26712 ) & (wr )  ;
assign n26714 =  ( n26713 ) ? ( n5071 ) : ( iram_226 ) ;
assign n26715 = wr_addr[7:7] ;
assign n26716 =  ( n26715 ) == ( bv_1_0_n53 )  ;
assign n26717 =  ( wr_addr ) == ( bv_8_226_n521 )  ;
assign n26718 =  ( n26716 ) & (n26717 )  ;
assign n26719 =  ( n26718 ) & (wr )  ;
assign n26720 =  ( n26719 ) ? ( n5096 ) : ( iram_226 ) ;
assign n26721 = wr_addr[7:7] ;
assign n26722 =  ( n26721 ) == ( bv_1_0_n53 )  ;
assign n26723 =  ( wr_addr ) == ( bv_8_226_n521 )  ;
assign n26724 =  ( n26722 ) & (n26723 )  ;
assign n26725 =  ( n26724 ) & (wr )  ;
assign n26726 =  ( n26725 ) ? ( n5123 ) : ( iram_226 ) ;
assign n26727 = wr_addr[7:7] ;
assign n26728 =  ( n26727 ) == ( bv_1_0_n53 )  ;
assign n26729 =  ( wr_addr ) == ( bv_8_226_n521 )  ;
assign n26730 =  ( n26728 ) & (n26729 )  ;
assign n26731 =  ( n26730 ) & (wr )  ;
assign n26732 =  ( n26731 ) ? ( n5165 ) : ( iram_226 ) ;
assign n26733 = wr_addr[7:7] ;
assign n26734 =  ( n26733 ) == ( bv_1_0_n53 )  ;
assign n26735 =  ( wr_addr ) == ( bv_8_226_n521 )  ;
assign n26736 =  ( n26734 ) & (n26735 )  ;
assign n26737 =  ( n26736 ) & (wr )  ;
assign n26738 =  ( n26737 ) ? ( n5204 ) : ( iram_226 ) ;
assign n26739 = wr_addr[7:7] ;
assign n26740 =  ( n26739 ) == ( bv_1_0_n53 )  ;
assign n26741 =  ( wr_addr ) == ( bv_8_226_n521 )  ;
assign n26742 =  ( n26740 ) & (n26741 )  ;
assign n26743 =  ( n26742 ) & (wr )  ;
assign n26744 =  ( n26743 ) ? ( n5262 ) : ( iram_226 ) ;
assign n26745 = wr_addr[7:7] ;
assign n26746 =  ( n26745 ) == ( bv_1_0_n53 )  ;
assign n26747 =  ( wr_addr ) == ( bv_8_226_n521 )  ;
assign n26748 =  ( n26746 ) & (n26747 )  ;
assign n26749 =  ( n26748 ) & (wr )  ;
assign n26750 =  ( n26749 ) ? ( n5298 ) : ( iram_226 ) ;
assign n26751 = wr_addr[7:7] ;
assign n26752 =  ( n26751 ) == ( bv_1_0_n53 )  ;
assign n26753 =  ( wr_addr ) == ( bv_8_226_n521 )  ;
assign n26754 =  ( n26752 ) & (n26753 )  ;
assign n26755 =  ( n26754 ) & (wr )  ;
assign n26756 =  ( n26755 ) ? ( n5325 ) : ( iram_226 ) ;
assign n26757 = wr_addr[7:7] ;
assign n26758 =  ( n26757 ) == ( bv_1_0_n53 )  ;
assign n26759 =  ( wr_addr ) == ( bv_8_227_n523 )  ;
assign n26760 =  ( n26758 ) & (n26759 )  ;
assign n26761 =  ( n26760 ) & (wr )  ;
assign n26762 =  ( n26761 ) ? ( n4782 ) : ( iram_227 ) ;
assign n26763 = wr_addr[7:7] ;
assign n26764 =  ( n26763 ) == ( bv_1_0_n53 )  ;
assign n26765 =  ( wr_addr ) == ( bv_8_227_n523 )  ;
assign n26766 =  ( n26764 ) & (n26765 )  ;
assign n26767 =  ( n26766 ) & (wr )  ;
assign n26768 =  ( n26767 ) ? ( n4841 ) : ( iram_227 ) ;
assign n26769 = wr_addr[7:7] ;
assign n26770 =  ( n26769 ) == ( bv_1_0_n53 )  ;
assign n26771 =  ( wr_addr ) == ( bv_8_227_n523 )  ;
assign n26772 =  ( n26770 ) & (n26771 )  ;
assign n26773 =  ( n26772 ) & (wr )  ;
assign n26774 =  ( n26773 ) ? ( n5449 ) : ( iram_227 ) ;
assign n26775 = wr_addr[7:7] ;
assign n26776 =  ( n26775 ) == ( bv_1_0_n53 )  ;
assign n26777 =  ( wr_addr ) == ( bv_8_227_n523 )  ;
assign n26778 =  ( n26776 ) & (n26777 )  ;
assign n26779 =  ( n26778 ) & (wr )  ;
assign n26780 =  ( n26779 ) ? ( n4906 ) : ( iram_227 ) ;
assign n26781 = wr_addr[7:7] ;
assign n26782 =  ( n26781 ) == ( bv_1_0_n53 )  ;
assign n26783 =  ( wr_addr ) == ( bv_8_227_n523 )  ;
assign n26784 =  ( n26782 ) & (n26783 )  ;
assign n26785 =  ( n26784 ) & (wr )  ;
assign n26786 =  ( n26785 ) ? ( n5485 ) : ( iram_227 ) ;
assign n26787 = wr_addr[7:7] ;
assign n26788 =  ( n26787 ) == ( bv_1_0_n53 )  ;
assign n26789 =  ( wr_addr ) == ( bv_8_227_n523 )  ;
assign n26790 =  ( n26788 ) & (n26789 )  ;
assign n26791 =  ( n26790 ) & (wr )  ;
assign n26792 =  ( n26791 ) ? ( n5512 ) : ( iram_227 ) ;
assign n26793 = wr_addr[7:7] ;
assign n26794 =  ( n26793 ) == ( bv_1_0_n53 )  ;
assign n26795 =  ( wr_addr ) == ( bv_8_227_n523 )  ;
assign n26796 =  ( n26794 ) & (n26795 )  ;
assign n26797 =  ( n26796 ) & (wr )  ;
assign n26798 =  ( n26797 ) ? ( bv_8_0_n69 ) : ( iram_227 ) ;
assign n26799 = wr_addr[7:7] ;
assign n26800 =  ( n26799 ) == ( bv_1_0_n53 )  ;
assign n26801 =  ( wr_addr ) == ( bv_8_227_n523 )  ;
assign n26802 =  ( n26800 ) & (n26801 )  ;
assign n26803 =  ( n26802 ) & (wr )  ;
assign n26804 =  ( n26803 ) ? ( n5071 ) : ( iram_227 ) ;
assign n26805 = wr_addr[7:7] ;
assign n26806 =  ( n26805 ) == ( bv_1_0_n53 )  ;
assign n26807 =  ( wr_addr ) == ( bv_8_227_n523 )  ;
assign n26808 =  ( n26806 ) & (n26807 )  ;
assign n26809 =  ( n26808 ) & (wr )  ;
assign n26810 =  ( n26809 ) ? ( n5096 ) : ( iram_227 ) ;
assign n26811 = wr_addr[7:7] ;
assign n26812 =  ( n26811 ) == ( bv_1_0_n53 )  ;
assign n26813 =  ( wr_addr ) == ( bv_8_227_n523 )  ;
assign n26814 =  ( n26812 ) & (n26813 )  ;
assign n26815 =  ( n26814 ) & (wr )  ;
assign n26816 =  ( n26815 ) ? ( n5123 ) : ( iram_227 ) ;
assign n26817 = wr_addr[7:7] ;
assign n26818 =  ( n26817 ) == ( bv_1_0_n53 )  ;
assign n26819 =  ( wr_addr ) == ( bv_8_227_n523 )  ;
assign n26820 =  ( n26818 ) & (n26819 )  ;
assign n26821 =  ( n26820 ) & (wr )  ;
assign n26822 =  ( n26821 ) ? ( n5165 ) : ( iram_227 ) ;
assign n26823 = wr_addr[7:7] ;
assign n26824 =  ( n26823 ) == ( bv_1_0_n53 )  ;
assign n26825 =  ( wr_addr ) == ( bv_8_227_n523 )  ;
assign n26826 =  ( n26824 ) & (n26825 )  ;
assign n26827 =  ( n26826 ) & (wr )  ;
assign n26828 =  ( n26827 ) ? ( n5204 ) : ( iram_227 ) ;
assign n26829 = wr_addr[7:7] ;
assign n26830 =  ( n26829 ) == ( bv_1_0_n53 )  ;
assign n26831 =  ( wr_addr ) == ( bv_8_227_n523 )  ;
assign n26832 =  ( n26830 ) & (n26831 )  ;
assign n26833 =  ( n26832 ) & (wr )  ;
assign n26834 =  ( n26833 ) ? ( n5262 ) : ( iram_227 ) ;
assign n26835 = wr_addr[7:7] ;
assign n26836 =  ( n26835 ) == ( bv_1_0_n53 )  ;
assign n26837 =  ( wr_addr ) == ( bv_8_227_n523 )  ;
assign n26838 =  ( n26836 ) & (n26837 )  ;
assign n26839 =  ( n26838 ) & (wr )  ;
assign n26840 =  ( n26839 ) ? ( n5298 ) : ( iram_227 ) ;
assign n26841 = wr_addr[7:7] ;
assign n26842 =  ( n26841 ) == ( bv_1_0_n53 )  ;
assign n26843 =  ( wr_addr ) == ( bv_8_227_n523 )  ;
assign n26844 =  ( n26842 ) & (n26843 )  ;
assign n26845 =  ( n26844 ) & (wr )  ;
assign n26846 =  ( n26845 ) ? ( n5325 ) : ( iram_227 ) ;
assign n26847 = wr_addr[7:7] ;
assign n26848 =  ( n26847 ) == ( bv_1_0_n53 )  ;
assign n26849 =  ( wr_addr ) == ( bv_8_228_n525 )  ;
assign n26850 =  ( n26848 ) & (n26849 )  ;
assign n26851 =  ( n26850 ) & (wr )  ;
assign n26852 =  ( n26851 ) ? ( n4782 ) : ( iram_228 ) ;
assign n26853 = wr_addr[7:7] ;
assign n26854 =  ( n26853 ) == ( bv_1_0_n53 )  ;
assign n26855 =  ( wr_addr ) == ( bv_8_228_n525 )  ;
assign n26856 =  ( n26854 ) & (n26855 )  ;
assign n26857 =  ( n26856 ) & (wr )  ;
assign n26858 =  ( n26857 ) ? ( n4841 ) : ( iram_228 ) ;
assign n26859 = wr_addr[7:7] ;
assign n26860 =  ( n26859 ) == ( bv_1_0_n53 )  ;
assign n26861 =  ( wr_addr ) == ( bv_8_228_n525 )  ;
assign n26862 =  ( n26860 ) & (n26861 )  ;
assign n26863 =  ( n26862 ) & (wr )  ;
assign n26864 =  ( n26863 ) ? ( n5449 ) : ( iram_228 ) ;
assign n26865 = wr_addr[7:7] ;
assign n26866 =  ( n26865 ) == ( bv_1_0_n53 )  ;
assign n26867 =  ( wr_addr ) == ( bv_8_228_n525 )  ;
assign n26868 =  ( n26866 ) & (n26867 )  ;
assign n26869 =  ( n26868 ) & (wr )  ;
assign n26870 =  ( n26869 ) ? ( n4906 ) : ( iram_228 ) ;
assign n26871 = wr_addr[7:7] ;
assign n26872 =  ( n26871 ) == ( bv_1_0_n53 )  ;
assign n26873 =  ( wr_addr ) == ( bv_8_228_n525 )  ;
assign n26874 =  ( n26872 ) & (n26873 )  ;
assign n26875 =  ( n26874 ) & (wr )  ;
assign n26876 =  ( n26875 ) ? ( n5485 ) : ( iram_228 ) ;
assign n26877 = wr_addr[7:7] ;
assign n26878 =  ( n26877 ) == ( bv_1_0_n53 )  ;
assign n26879 =  ( wr_addr ) == ( bv_8_228_n525 )  ;
assign n26880 =  ( n26878 ) & (n26879 )  ;
assign n26881 =  ( n26880 ) & (wr )  ;
assign n26882 =  ( n26881 ) ? ( n5512 ) : ( iram_228 ) ;
assign n26883 = wr_addr[7:7] ;
assign n26884 =  ( n26883 ) == ( bv_1_0_n53 )  ;
assign n26885 =  ( wr_addr ) == ( bv_8_228_n525 )  ;
assign n26886 =  ( n26884 ) & (n26885 )  ;
assign n26887 =  ( n26886 ) & (wr )  ;
assign n26888 =  ( n26887 ) ? ( bv_8_0_n69 ) : ( iram_228 ) ;
assign n26889 = wr_addr[7:7] ;
assign n26890 =  ( n26889 ) == ( bv_1_0_n53 )  ;
assign n26891 =  ( wr_addr ) == ( bv_8_228_n525 )  ;
assign n26892 =  ( n26890 ) & (n26891 )  ;
assign n26893 =  ( n26892 ) & (wr )  ;
assign n26894 =  ( n26893 ) ? ( n5071 ) : ( iram_228 ) ;
assign n26895 = wr_addr[7:7] ;
assign n26896 =  ( n26895 ) == ( bv_1_0_n53 )  ;
assign n26897 =  ( wr_addr ) == ( bv_8_228_n525 )  ;
assign n26898 =  ( n26896 ) & (n26897 )  ;
assign n26899 =  ( n26898 ) & (wr )  ;
assign n26900 =  ( n26899 ) ? ( n5096 ) : ( iram_228 ) ;
assign n26901 = wr_addr[7:7] ;
assign n26902 =  ( n26901 ) == ( bv_1_0_n53 )  ;
assign n26903 =  ( wr_addr ) == ( bv_8_228_n525 )  ;
assign n26904 =  ( n26902 ) & (n26903 )  ;
assign n26905 =  ( n26904 ) & (wr )  ;
assign n26906 =  ( n26905 ) ? ( n5123 ) : ( iram_228 ) ;
assign n26907 = wr_addr[7:7] ;
assign n26908 =  ( n26907 ) == ( bv_1_0_n53 )  ;
assign n26909 =  ( wr_addr ) == ( bv_8_228_n525 )  ;
assign n26910 =  ( n26908 ) & (n26909 )  ;
assign n26911 =  ( n26910 ) & (wr )  ;
assign n26912 =  ( n26911 ) ? ( n5165 ) : ( iram_228 ) ;
assign n26913 = wr_addr[7:7] ;
assign n26914 =  ( n26913 ) == ( bv_1_0_n53 )  ;
assign n26915 =  ( wr_addr ) == ( bv_8_228_n525 )  ;
assign n26916 =  ( n26914 ) & (n26915 )  ;
assign n26917 =  ( n26916 ) & (wr )  ;
assign n26918 =  ( n26917 ) ? ( n5204 ) : ( iram_228 ) ;
assign n26919 = wr_addr[7:7] ;
assign n26920 =  ( n26919 ) == ( bv_1_0_n53 )  ;
assign n26921 =  ( wr_addr ) == ( bv_8_228_n525 )  ;
assign n26922 =  ( n26920 ) & (n26921 )  ;
assign n26923 =  ( n26922 ) & (wr )  ;
assign n26924 =  ( n26923 ) ? ( n5262 ) : ( iram_228 ) ;
assign n26925 = wr_addr[7:7] ;
assign n26926 =  ( n26925 ) == ( bv_1_0_n53 )  ;
assign n26927 =  ( wr_addr ) == ( bv_8_228_n525 )  ;
assign n26928 =  ( n26926 ) & (n26927 )  ;
assign n26929 =  ( n26928 ) & (wr )  ;
assign n26930 =  ( n26929 ) ? ( n5298 ) : ( iram_228 ) ;
assign n26931 = wr_addr[7:7] ;
assign n26932 =  ( n26931 ) == ( bv_1_0_n53 )  ;
assign n26933 =  ( wr_addr ) == ( bv_8_228_n525 )  ;
assign n26934 =  ( n26932 ) & (n26933 )  ;
assign n26935 =  ( n26934 ) & (wr )  ;
assign n26936 =  ( n26935 ) ? ( n5325 ) : ( iram_228 ) ;
assign n26937 = wr_addr[7:7] ;
assign n26938 =  ( n26937 ) == ( bv_1_0_n53 )  ;
assign n26939 =  ( wr_addr ) == ( bv_8_229_n527 )  ;
assign n26940 =  ( n26938 ) & (n26939 )  ;
assign n26941 =  ( n26940 ) & (wr )  ;
assign n26942 =  ( n26941 ) ? ( n4782 ) : ( iram_229 ) ;
assign n26943 = wr_addr[7:7] ;
assign n26944 =  ( n26943 ) == ( bv_1_0_n53 )  ;
assign n26945 =  ( wr_addr ) == ( bv_8_229_n527 )  ;
assign n26946 =  ( n26944 ) & (n26945 )  ;
assign n26947 =  ( n26946 ) & (wr )  ;
assign n26948 =  ( n26947 ) ? ( n4841 ) : ( iram_229 ) ;
assign n26949 = wr_addr[7:7] ;
assign n26950 =  ( n26949 ) == ( bv_1_0_n53 )  ;
assign n26951 =  ( wr_addr ) == ( bv_8_229_n527 )  ;
assign n26952 =  ( n26950 ) & (n26951 )  ;
assign n26953 =  ( n26952 ) & (wr )  ;
assign n26954 =  ( n26953 ) ? ( n5449 ) : ( iram_229 ) ;
assign n26955 = wr_addr[7:7] ;
assign n26956 =  ( n26955 ) == ( bv_1_0_n53 )  ;
assign n26957 =  ( wr_addr ) == ( bv_8_229_n527 )  ;
assign n26958 =  ( n26956 ) & (n26957 )  ;
assign n26959 =  ( n26958 ) & (wr )  ;
assign n26960 =  ( n26959 ) ? ( n4906 ) : ( iram_229 ) ;
assign n26961 = wr_addr[7:7] ;
assign n26962 =  ( n26961 ) == ( bv_1_0_n53 )  ;
assign n26963 =  ( wr_addr ) == ( bv_8_229_n527 )  ;
assign n26964 =  ( n26962 ) & (n26963 )  ;
assign n26965 =  ( n26964 ) & (wr )  ;
assign n26966 =  ( n26965 ) ? ( n5485 ) : ( iram_229 ) ;
assign n26967 = wr_addr[7:7] ;
assign n26968 =  ( n26967 ) == ( bv_1_0_n53 )  ;
assign n26969 =  ( wr_addr ) == ( bv_8_229_n527 )  ;
assign n26970 =  ( n26968 ) & (n26969 )  ;
assign n26971 =  ( n26970 ) & (wr )  ;
assign n26972 =  ( n26971 ) ? ( n5512 ) : ( iram_229 ) ;
assign n26973 = wr_addr[7:7] ;
assign n26974 =  ( n26973 ) == ( bv_1_0_n53 )  ;
assign n26975 =  ( wr_addr ) == ( bv_8_229_n527 )  ;
assign n26976 =  ( n26974 ) & (n26975 )  ;
assign n26977 =  ( n26976 ) & (wr )  ;
assign n26978 =  ( n26977 ) ? ( bv_8_0_n69 ) : ( iram_229 ) ;
assign n26979 = wr_addr[7:7] ;
assign n26980 =  ( n26979 ) == ( bv_1_0_n53 )  ;
assign n26981 =  ( wr_addr ) == ( bv_8_229_n527 )  ;
assign n26982 =  ( n26980 ) & (n26981 )  ;
assign n26983 =  ( n26982 ) & (wr )  ;
assign n26984 =  ( n26983 ) ? ( n5071 ) : ( iram_229 ) ;
assign n26985 = wr_addr[7:7] ;
assign n26986 =  ( n26985 ) == ( bv_1_0_n53 )  ;
assign n26987 =  ( wr_addr ) == ( bv_8_229_n527 )  ;
assign n26988 =  ( n26986 ) & (n26987 )  ;
assign n26989 =  ( n26988 ) & (wr )  ;
assign n26990 =  ( n26989 ) ? ( n5096 ) : ( iram_229 ) ;
assign n26991 = wr_addr[7:7] ;
assign n26992 =  ( n26991 ) == ( bv_1_0_n53 )  ;
assign n26993 =  ( wr_addr ) == ( bv_8_229_n527 )  ;
assign n26994 =  ( n26992 ) & (n26993 )  ;
assign n26995 =  ( n26994 ) & (wr )  ;
assign n26996 =  ( n26995 ) ? ( n5123 ) : ( iram_229 ) ;
assign n26997 = wr_addr[7:7] ;
assign n26998 =  ( n26997 ) == ( bv_1_0_n53 )  ;
assign n26999 =  ( wr_addr ) == ( bv_8_229_n527 )  ;
assign n27000 =  ( n26998 ) & (n26999 )  ;
assign n27001 =  ( n27000 ) & (wr )  ;
assign n27002 =  ( n27001 ) ? ( n5165 ) : ( iram_229 ) ;
assign n27003 = wr_addr[7:7] ;
assign n27004 =  ( n27003 ) == ( bv_1_0_n53 )  ;
assign n27005 =  ( wr_addr ) == ( bv_8_229_n527 )  ;
assign n27006 =  ( n27004 ) & (n27005 )  ;
assign n27007 =  ( n27006 ) & (wr )  ;
assign n27008 =  ( n27007 ) ? ( n5204 ) : ( iram_229 ) ;
assign n27009 = wr_addr[7:7] ;
assign n27010 =  ( n27009 ) == ( bv_1_0_n53 )  ;
assign n27011 =  ( wr_addr ) == ( bv_8_229_n527 )  ;
assign n27012 =  ( n27010 ) & (n27011 )  ;
assign n27013 =  ( n27012 ) & (wr )  ;
assign n27014 =  ( n27013 ) ? ( n5262 ) : ( iram_229 ) ;
assign n27015 = wr_addr[7:7] ;
assign n27016 =  ( n27015 ) == ( bv_1_0_n53 )  ;
assign n27017 =  ( wr_addr ) == ( bv_8_229_n527 )  ;
assign n27018 =  ( n27016 ) & (n27017 )  ;
assign n27019 =  ( n27018 ) & (wr )  ;
assign n27020 =  ( n27019 ) ? ( n5298 ) : ( iram_229 ) ;
assign n27021 = wr_addr[7:7] ;
assign n27022 =  ( n27021 ) == ( bv_1_0_n53 )  ;
assign n27023 =  ( wr_addr ) == ( bv_8_229_n527 )  ;
assign n27024 =  ( n27022 ) & (n27023 )  ;
assign n27025 =  ( n27024 ) & (wr )  ;
assign n27026 =  ( n27025 ) ? ( n5325 ) : ( iram_229 ) ;
assign n27027 = wr_addr[7:7] ;
assign n27028 =  ( n27027 ) == ( bv_1_0_n53 )  ;
assign n27029 =  ( wr_addr ) == ( bv_8_230_n529 )  ;
assign n27030 =  ( n27028 ) & (n27029 )  ;
assign n27031 =  ( n27030 ) & (wr )  ;
assign n27032 =  ( n27031 ) ? ( n4782 ) : ( iram_230 ) ;
assign n27033 = wr_addr[7:7] ;
assign n27034 =  ( n27033 ) == ( bv_1_0_n53 )  ;
assign n27035 =  ( wr_addr ) == ( bv_8_230_n529 )  ;
assign n27036 =  ( n27034 ) & (n27035 )  ;
assign n27037 =  ( n27036 ) & (wr )  ;
assign n27038 =  ( n27037 ) ? ( n4841 ) : ( iram_230 ) ;
assign n27039 = wr_addr[7:7] ;
assign n27040 =  ( n27039 ) == ( bv_1_0_n53 )  ;
assign n27041 =  ( wr_addr ) == ( bv_8_230_n529 )  ;
assign n27042 =  ( n27040 ) & (n27041 )  ;
assign n27043 =  ( n27042 ) & (wr )  ;
assign n27044 =  ( n27043 ) ? ( n5449 ) : ( iram_230 ) ;
assign n27045 = wr_addr[7:7] ;
assign n27046 =  ( n27045 ) == ( bv_1_0_n53 )  ;
assign n27047 =  ( wr_addr ) == ( bv_8_230_n529 )  ;
assign n27048 =  ( n27046 ) & (n27047 )  ;
assign n27049 =  ( n27048 ) & (wr )  ;
assign n27050 =  ( n27049 ) ? ( n4906 ) : ( iram_230 ) ;
assign n27051 = wr_addr[7:7] ;
assign n27052 =  ( n27051 ) == ( bv_1_0_n53 )  ;
assign n27053 =  ( wr_addr ) == ( bv_8_230_n529 )  ;
assign n27054 =  ( n27052 ) & (n27053 )  ;
assign n27055 =  ( n27054 ) & (wr )  ;
assign n27056 =  ( n27055 ) ? ( n5485 ) : ( iram_230 ) ;
assign n27057 = wr_addr[7:7] ;
assign n27058 =  ( n27057 ) == ( bv_1_0_n53 )  ;
assign n27059 =  ( wr_addr ) == ( bv_8_230_n529 )  ;
assign n27060 =  ( n27058 ) & (n27059 )  ;
assign n27061 =  ( n27060 ) & (wr )  ;
assign n27062 =  ( n27061 ) ? ( n5512 ) : ( iram_230 ) ;
assign n27063 = wr_addr[7:7] ;
assign n27064 =  ( n27063 ) == ( bv_1_0_n53 )  ;
assign n27065 =  ( wr_addr ) == ( bv_8_230_n529 )  ;
assign n27066 =  ( n27064 ) & (n27065 )  ;
assign n27067 =  ( n27066 ) & (wr )  ;
assign n27068 =  ( n27067 ) ? ( bv_8_0_n69 ) : ( iram_230 ) ;
assign n27069 = wr_addr[7:7] ;
assign n27070 =  ( n27069 ) == ( bv_1_0_n53 )  ;
assign n27071 =  ( wr_addr ) == ( bv_8_230_n529 )  ;
assign n27072 =  ( n27070 ) & (n27071 )  ;
assign n27073 =  ( n27072 ) & (wr )  ;
assign n27074 =  ( n27073 ) ? ( n5071 ) : ( iram_230 ) ;
assign n27075 = wr_addr[7:7] ;
assign n27076 =  ( n27075 ) == ( bv_1_0_n53 )  ;
assign n27077 =  ( wr_addr ) == ( bv_8_230_n529 )  ;
assign n27078 =  ( n27076 ) & (n27077 )  ;
assign n27079 =  ( n27078 ) & (wr )  ;
assign n27080 =  ( n27079 ) ? ( n5096 ) : ( iram_230 ) ;
assign n27081 = wr_addr[7:7] ;
assign n27082 =  ( n27081 ) == ( bv_1_0_n53 )  ;
assign n27083 =  ( wr_addr ) == ( bv_8_230_n529 )  ;
assign n27084 =  ( n27082 ) & (n27083 )  ;
assign n27085 =  ( n27084 ) & (wr )  ;
assign n27086 =  ( n27085 ) ? ( n5123 ) : ( iram_230 ) ;
assign n27087 = wr_addr[7:7] ;
assign n27088 =  ( n27087 ) == ( bv_1_0_n53 )  ;
assign n27089 =  ( wr_addr ) == ( bv_8_230_n529 )  ;
assign n27090 =  ( n27088 ) & (n27089 )  ;
assign n27091 =  ( n27090 ) & (wr )  ;
assign n27092 =  ( n27091 ) ? ( n5165 ) : ( iram_230 ) ;
assign n27093 = wr_addr[7:7] ;
assign n27094 =  ( n27093 ) == ( bv_1_0_n53 )  ;
assign n27095 =  ( wr_addr ) == ( bv_8_230_n529 )  ;
assign n27096 =  ( n27094 ) & (n27095 )  ;
assign n27097 =  ( n27096 ) & (wr )  ;
assign n27098 =  ( n27097 ) ? ( n5204 ) : ( iram_230 ) ;
assign n27099 = wr_addr[7:7] ;
assign n27100 =  ( n27099 ) == ( bv_1_0_n53 )  ;
assign n27101 =  ( wr_addr ) == ( bv_8_230_n529 )  ;
assign n27102 =  ( n27100 ) & (n27101 )  ;
assign n27103 =  ( n27102 ) & (wr )  ;
assign n27104 =  ( n27103 ) ? ( n5262 ) : ( iram_230 ) ;
assign n27105 = wr_addr[7:7] ;
assign n27106 =  ( n27105 ) == ( bv_1_0_n53 )  ;
assign n27107 =  ( wr_addr ) == ( bv_8_230_n529 )  ;
assign n27108 =  ( n27106 ) & (n27107 )  ;
assign n27109 =  ( n27108 ) & (wr )  ;
assign n27110 =  ( n27109 ) ? ( n5298 ) : ( iram_230 ) ;
assign n27111 = wr_addr[7:7] ;
assign n27112 =  ( n27111 ) == ( bv_1_0_n53 )  ;
assign n27113 =  ( wr_addr ) == ( bv_8_230_n529 )  ;
assign n27114 =  ( n27112 ) & (n27113 )  ;
assign n27115 =  ( n27114 ) & (wr )  ;
assign n27116 =  ( n27115 ) ? ( n5325 ) : ( iram_230 ) ;
assign n27117 = wr_addr[7:7] ;
assign n27118 =  ( n27117 ) == ( bv_1_0_n53 )  ;
assign n27119 =  ( wr_addr ) == ( bv_8_231_n531 )  ;
assign n27120 =  ( n27118 ) & (n27119 )  ;
assign n27121 =  ( n27120 ) & (wr )  ;
assign n27122 =  ( n27121 ) ? ( n4782 ) : ( iram_231 ) ;
assign n27123 = wr_addr[7:7] ;
assign n27124 =  ( n27123 ) == ( bv_1_0_n53 )  ;
assign n27125 =  ( wr_addr ) == ( bv_8_231_n531 )  ;
assign n27126 =  ( n27124 ) & (n27125 )  ;
assign n27127 =  ( n27126 ) & (wr )  ;
assign n27128 =  ( n27127 ) ? ( n4841 ) : ( iram_231 ) ;
assign n27129 = wr_addr[7:7] ;
assign n27130 =  ( n27129 ) == ( bv_1_0_n53 )  ;
assign n27131 =  ( wr_addr ) == ( bv_8_231_n531 )  ;
assign n27132 =  ( n27130 ) & (n27131 )  ;
assign n27133 =  ( n27132 ) & (wr )  ;
assign n27134 =  ( n27133 ) ? ( n5449 ) : ( iram_231 ) ;
assign n27135 = wr_addr[7:7] ;
assign n27136 =  ( n27135 ) == ( bv_1_0_n53 )  ;
assign n27137 =  ( wr_addr ) == ( bv_8_231_n531 )  ;
assign n27138 =  ( n27136 ) & (n27137 )  ;
assign n27139 =  ( n27138 ) & (wr )  ;
assign n27140 =  ( n27139 ) ? ( n4906 ) : ( iram_231 ) ;
assign n27141 = wr_addr[7:7] ;
assign n27142 =  ( n27141 ) == ( bv_1_0_n53 )  ;
assign n27143 =  ( wr_addr ) == ( bv_8_231_n531 )  ;
assign n27144 =  ( n27142 ) & (n27143 )  ;
assign n27145 =  ( n27144 ) & (wr )  ;
assign n27146 =  ( n27145 ) ? ( n5485 ) : ( iram_231 ) ;
assign n27147 = wr_addr[7:7] ;
assign n27148 =  ( n27147 ) == ( bv_1_0_n53 )  ;
assign n27149 =  ( wr_addr ) == ( bv_8_231_n531 )  ;
assign n27150 =  ( n27148 ) & (n27149 )  ;
assign n27151 =  ( n27150 ) & (wr )  ;
assign n27152 =  ( n27151 ) ? ( n5512 ) : ( iram_231 ) ;
assign n27153 = wr_addr[7:7] ;
assign n27154 =  ( n27153 ) == ( bv_1_0_n53 )  ;
assign n27155 =  ( wr_addr ) == ( bv_8_231_n531 )  ;
assign n27156 =  ( n27154 ) & (n27155 )  ;
assign n27157 =  ( n27156 ) & (wr )  ;
assign n27158 =  ( n27157 ) ? ( bv_8_0_n69 ) : ( iram_231 ) ;
assign n27159 = wr_addr[7:7] ;
assign n27160 =  ( n27159 ) == ( bv_1_0_n53 )  ;
assign n27161 =  ( wr_addr ) == ( bv_8_231_n531 )  ;
assign n27162 =  ( n27160 ) & (n27161 )  ;
assign n27163 =  ( n27162 ) & (wr )  ;
assign n27164 =  ( n27163 ) ? ( n5071 ) : ( iram_231 ) ;
assign n27165 = wr_addr[7:7] ;
assign n27166 =  ( n27165 ) == ( bv_1_0_n53 )  ;
assign n27167 =  ( wr_addr ) == ( bv_8_231_n531 )  ;
assign n27168 =  ( n27166 ) & (n27167 )  ;
assign n27169 =  ( n27168 ) & (wr )  ;
assign n27170 =  ( n27169 ) ? ( n5096 ) : ( iram_231 ) ;
assign n27171 = wr_addr[7:7] ;
assign n27172 =  ( n27171 ) == ( bv_1_0_n53 )  ;
assign n27173 =  ( wr_addr ) == ( bv_8_231_n531 )  ;
assign n27174 =  ( n27172 ) & (n27173 )  ;
assign n27175 =  ( n27174 ) & (wr )  ;
assign n27176 =  ( n27175 ) ? ( n5123 ) : ( iram_231 ) ;
assign n27177 = wr_addr[7:7] ;
assign n27178 =  ( n27177 ) == ( bv_1_0_n53 )  ;
assign n27179 =  ( wr_addr ) == ( bv_8_231_n531 )  ;
assign n27180 =  ( n27178 ) & (n27179 )  ;
assign n27181 =  ( n27180 ) & (wr )  ;
assign n27182 =  ( n27181 ) ? ( n5165 ) : ( iram_231 ) ;
assign n27183 = wr_addr[7:7] ;
assign n27184 =  ( n27183 ) == ( bv_1_0_n53 )  ;
assign n27185 =  ( wr_addr ) == ( bv_8_231_n531 )  ;
assign n27186 =  ( n27184 ) & (n27185 )  ;
assign n27187 =  ( n27186 ) & (wr )  ;
assign n27188 =  ( n27187 ) ? ( n5204 ) : ( iram_231 ) ;
assign n27189 = wr_addr[7:7] ;
assign n27190 =  ( n27189 ) == ( bv_1_0_n53 )  ;
assign n27191 =  ( wr_addr ) == ( bv_8_231_n531 )  ;
assign n27192 =  ( n27190 ) & (n27191 )  ;
assign n27193 =  ( n27192 ) & (wr )  ;
assign n27194 =  ( n27193 ) ? ( n5262 ) : ( iram_231 ) ;
assign n27195 = wr_addr[7:7] ;
assign n27196 =  ( n27195 ) == ( bv_1_0_n53 )  ;
assign n27197 =  ( wr_addr ) == ( bv_8_231_n531 )  ;
assign n27198 =  ( n27196 ) & (n27197 )  ;
assign n27199 =  ( n27198 ) & (wr )  ;
assign n27200 =  ( n27199 ) ? ( n5298 ) : ( iram_231 ) ;
assign n27201 = wr_addr[7:7] ;
assign n27202 =  ( n27201 ) == ( bv_1_0_n53 )  ;
assign n27203 =  ( wr_addr ) == ( bv_8_231_n531 )  ;
assign n27204 =  ( n27202 ) & (n27203 )  ;
assign n27205 =  ( n27204 ) & (wr )  ;
assign n27206 =  ( n27205 ) ? ( n5325 ) : ( iram_231 ) ;
assign n27207 = wr_addr[7:7] ;
assign n27208 =  ( n27207 ) == ( bv_1_0_n53 )  ;
assign n27209 =  ( wr_addr ) == ( bv_8_232_n533 )  ;
assign n27210 =  ( n27208 ) & (n27209 )  ;
assign n27211 =  ( n27210 ) & (wr )  ;
assign n27212 =  ( n27211 ) ? ( n4782 ) : ( iram_232 ) ;
assign n27213 = wr_addr[7:7] ;
assign n27214 =  ( n27213 ) == ( bv_1_0_n53 )  ;
assign n27215 =  ( wr_addr ) == ( bv_8_232_n533 )  ;
assign n27216 =  ( n27214 ) & (n27215 )  ;
assign n27217 =  ( n27216 ) & (wr )  ;
assign n27218 =  ( n27217 ) ? ( n4841 ) : ( iram_232 ) ;
assign n27219 = wr_addr[7:7] ;
assign n27220 =  ( n27219 ) == ( bv_1_0_n53 )  ;
assign n27221 =  ( wr_addr ) == ( bv_8_232_n533 )  ;
assign n27222 =  ( n27220 ) & (n27221 )  ;
assign n27223 =  ( n27222 ) & (wr )  ;
assign n27224 =  ( n27223 ) ? ( n5449 ) : ( iram_232 ) ;
assign n27225 = wr_addr[7:7] ;
assign n27226 =  ( n27225 ) == ( bv_1_0_n53 )  ;
assign n27227 =  ( wr_addr ) == ( bv_8_232_n533 )  ;
assign n27228 =  ( n27226 ) & (n27227 )  ;
assign n27229 =  ( n27228 ) & (wr )  ;
assign n27230 =  ( n27229 ) ? ( n4906 ) : ( iram_232 ) ;
assign n27231 = wr_addr[7:7] ;
assign n27232 =  ( n27231 ) == ( bv_1_0_n53 )  ;
assign n27233 =  ( wr_addr ) == ( bv_8_232_n533 )  ;
assign n27234 =  ( n27232 ) & (n27233 )  ;
assign n27235 =  ( n27234 ) & (wr )  ;
assign n27236 =  ( n27235 ) ? ( n5485 ) : ( iram_232 ) ;
assign n27237 = wr_addr[7:7] ;
assign n27238 =  ( n27237 ) == ( bv_1_0_n53 )  ;
assign n27239 =  ( wr_addr ) == ( bv_8_232_n533 )  ;
assign n27240 =  ( n27238 ) & (n27239 )  ;
assign n27241 =  ( n27240 ) & (wr )  ;
assign n27242 =  ( n27241 ) ? ( n5512 ) : ( iram_232 ) ;
assign n27243 = wr_addr[7:7] ;
assign n27244 =  ( n27243 ) == ( bv_1_0_n53 )  ;
assign n27245 =  ( wr_addr ) == ( bv_8_232_n533 )  ;
assign n27246 =  ( n27244 ) & (n27245 )  ;
assign n27247 =  ( n27246 ) & (wr )  ;
assign n27248 =  ( n27247 ) ? ( bv_8_0_n69 ) : ( iram_232 ) ;
assign n27249 = wr_addr[7:7] ;
assign n27250 =  ( n27249 ) == ( bv_1_0_n53 )  ;
assign n27251 =  ( wr_addr ) == ( bv_8_232_n533 )  ;
assign n27252 =  ( n27250 ) & (n27251 )  ;
assign n27253 =  ( n27252 ) & (wr )  ;
assign n27254 =  ( n27253 ) ? ( n5071 ) : ( iram_232 ) ;
assign n27255 = wr_addr[7:7] ;
assign n27256 =  ( n27255 ) == ( bv_1_0_n53 )  ;
assign n27257 =  ( wr_addr ) == ( bv_8_232_n533 )  ;
assign n27258 =  ( n27256 ) & (n27257 )  ;
assign n27259 =  ( n27258 ) & (wr )  ;
assign n27260 =  ( n27259 ) ? ( n5096 ) : ( iram_232 ) ;
assign n27261 = wr_addr[7:7] ;
assign n27262 =  ( n27261 ) == ( bv_1_0_n53 )  ;
assign n27263 =  ( wr_addr ) == ( bv_8_232_n533 )  ;
assign n27264 =  ( n27262 ) & (n27263 )  ;
assign n27265 =  ( n27264 ) & (wr )  ;
assign n27266 =  ( n27265 ) ? ( n5123 ) : ( iram_232 ) ;
assign n27267 = wr_addr[7:7] ;
assign n27268 =  ( n27267 ) == ( bv_1_0_n53 )  ;
assign n27269 =  ( wr_addr ) == ( bv_8_232_n533 )  ;
assign n27270 =  ( n27268 ) & (n27269 )  ;
assign n27271 =  ( n27270 ) & (wr )  ;
assign n27272 =  ( n27271 ) ? ( n5165 ) : ( iram_232 ) ;
assign n27273 = wr_addr[7:7] ;
assign n27274 =  ( n27273 ) == ( bv_1_0_n53 )  ;
assign n27275 =  ( wr_addr ) == ( bv_8_232_n533 )  ;
assign n27276 =  ( n27274 ) & (n27275 )  ;
assign n27277 =  ( n27276 ) & (wr )  ;
assign n27278 =  ( n27277 ) ? ( n5204 ) : ( iram_232 ) ;
assign n27279 = wr_addr[7:7] ;
assign n27280 =  ( n27279 ) == ( bv_1_0_n53 )  ;
assign n27281 =  ( wr_addr ) == ( bv_8_232_n533 )  ;
assign n27282 =  ( n27280 ) & (n27281 )  ;
assign n27283 =  ( n27282 ) & (wr )  ;
assign n27284 =  ( n27283 ) ? ( n5262 ) : ( iram_232 ) ;
assign n27285 = wr_addr[7:7] ;
assign n27286 =  ( n27285 ) == ( bv_1_0_n53 )  ;
assign n27287 =  ( wr_addr ) == ( bv_8_232_n533 )  ;
assign n27288 =  ( n27286 ) & (n27287 )  ;
assign n27289 =  ( n27288 ) & (wr )  ;
assign n27290 =  ( n27289 ) ? ( n5298 ) : ( iram_232 ) ;
assign n27291 = wr_addr[7:7] ;
assign n27292 =  ( n27291 ) == ( bv_1_0_n53 )  ;
assign n27293 =  ( wr_addr ) == ( bv_8_232_n533 )  ;
assign n27294 =  ( n27292 ) & (n27293 )  ;
assign n27295 =  ( n27294 ) & (wr )  ;
assign n27296 =  ( n27295 ) ? ( n5325 ) : ( iram_232 ) ;
assign n27297 = wr_addr[7:7] ;
assign n27298 =  ( n27297 ) == ( bv_1_0_n53 )  ;
assign n27299 =  ( wr_addr ) == ( bv_8_233_n535 )  ;
assign n27300 =  ( n27298 ) & (n27299 )  ;
assign n27301 =  ( n27300 ) & (wr )  ;
assign n27302 =  ( n27301 ) ? ( n4782 ) : ( iram_233 ) ;
assign n27303 = wr_addr[7:7] ;
assign n27304 =  ( n27303 ) == ( bv_1_0_n53 )  ;
assign n27305 =  ( wr_addr ) == ( bv_8_233_n535 )  ;
assign n27306 =  ( n27304 ) & (n27305 )  ;
assign n27307 =  ( n27306 ) & (wr )  ;
assign n27308 =  ( n27307 ) ? ( n4841 ) : ( iram_233 ) ;
assign n27309 = wr_addr[7:7] ;
assign n27310 =  ( n27309 ) == ( bv_1_0_n53 )  ;
assign n27311 =  ( wr_addr ) == ( bv_8_233_n535 )  ;
assign n27312 =  ( n27310 ) & (n27311 )  ;
assign n27313 =  ( n27312 ) & (wr )  ;
assign n27314 =  ( n27313 ) ? ( n5449 ) : ( iram_233 ) ;
assign n27315 = wr_addr[7:7] ;
assign n27316 =  ( n27315 ) == ( bv_1_0_n53 )  ;
assign n27317 =  ( wr_addr ) == ( bv_8_233_n535 )  ;
assign n27318 =  ( n27316 ) & (n27317 )  ;
assign n27319 =  ( n27318 ) & (wr )  ;
assign n27320 =  ( n27319 ) ? ( n4906 ) : ( iram_233 ) ;
assign n27321 = wr_addr[7:7] ;
assign n27322 =  ( n27321 ) == ( bv_1_0_n53 )  ;
assign n27323 =  ( wr_addr ) == ( bv_8_233_n535 )  ;
assign n27324 =  ( n27322 ) & (n27323 )  ;
assign n27325 =  ( n27324 ) & (wr )  ;
assign n27326 =  ( n27325 ) ? ( n5485 ) : ( iram_233 ) ;
assign n27327 = wr_addr[7:7] ;
assign n27328 =  ( n27327 ) == ( bv_1_0_n53 )  ;
assign n27329 =  ( wr_addr ) == ( bv_8_233_n535 )  ;
assign n27330 =  ( n27328 ) & (n27329 )  ;
assign n27331 =  ( n27330 ) & (wr )  ;
assign n27332 =  ( n27331 ) ? ( n5512 ) : ( iram_233 ) ;
assign n27333 = wr_addr[7:7] ;
assign n27334 =  ( n27333 ) == ( bv_1_0_n53 )  ;
assign n27335 =  ( wr_addr ) == ( bv_8_233_n535 )  ;
assign n27336 =  ( n27334 ) & (n27335 )  ;
assign n27337 =  ( n27336 ) & (wr )  ;
assign n27338 =  ( n27337 ) ? ( bv_8_0_n69 ) : ( iram_233 ) ;
assign n27339 = wr_addr[7:7] ;
assign n27340 =  ( n27339 ) == ( bv_1_0_n53 )  ;
assign n27341 =  ( wr_addr ) == ( bv_8_233_n535 )  ;
assign n27342 =  ( n27340 ) & (n27341 )  ;
assign n27343 =  ( n27342 ) & (wr )  ;
assign n27344 =  ( n27343 ) ? ( n5071 ) : ( iram_233 ) ;
assign n27345 = wr_addr[7:7] ;
assign n27346 =  ( n27345 ) == ( bv_1_0_n53 )  ;
assign n27347 =  ( wr_addr ) == ( bv_8_233_n535 )  ;
assign n27348 =  ( n27346 ) & (n27347 )  ;
assign n27349 =  ( n27348 ) & (wr )  ;
assign n27350 =  ( n27349 ) ? ( n5096 ) : ( iram_233 ) ;
assign n27351 = wr_addr[7:7] ;
assign n27352 =  ( n27351 ) == ( bv_1_0_n53 )  ;
assign n27353 =  ( wr_addr ) == ( bv_8_233_n535 )  ;
assign n27354 =  ( n27352 ) & (n27353 )  ;
assign n27355 =  ( n27354 ) & (wr )  ;
assign n27356 =  ( n27355 ) ? ( n5123 ) : ( iram_233 ) ;
assign n27357 = wr_addr[7:7] ;
assign n27358 =  ( n27357 ) == ( bv_1_0_n53 )  ;
assign n27359 =  ( wr_addr ) == ( bv_8_233_n535 )  ;
assign n27360 =  ( n27358 ) & (n27359 )  ;
assign n27361 =  ( n27360 ) & (wr )  ;
assign n27362 =  ( n27361 ) ? ( n5165 ) : ( iram_233 ) ;
assign n27363 = wr_addr[7:7] ;
assign n27364 =  ( n27363 ) == ( bv_1_0_n53 )  ;
assign n27365 =  ( wr_addr ) == ( bv_8_233_n535 )  ;
assign n27366 =  ( n27364 ) & (n27365 )  ;
assign n27367 =  ( n27366 ) & (wr )  ;
assign n27368 =  ( n27367 ) ? ( n5204 ) : ( iram_233 ) ;
assign n27369 = wr_addr[7:7] ;
assign n27370 =  ( n27369 ) == ( bv_1_0_n53 )  ;
assign n27371 =  ( wr_addr ) == ( bv_8_233_n535 )  ;
assign n27372 =  ( n27370 ) & (n27371 )  ;
assign n27373 =  ( n27372 ) & (wr )  ;
assign n27374 =  ( n27373 ) ? ( n5262 ) : ( iram_233 ) ;
assign n27375 = wr_addr[7:7] ;
assign n27376 =  ( n27375 ) == ( bv_1_0_n53 )  ;
assign n27377 =  ( wr_addr ) == ( bv_8_233_n535 )  ;
assign n27378 =  ( n27376 ) & (n27377 )  ;
assign n27379 =  ( n27378 ) & (wr )  ;
assign n27380 =  ( n27379 ) ? ( n5298 ) : ( iram_233 ) ;
assign n27381 = wr_addr[7:7] ;
assign n27382 =  ( n27381 ) == ( bv_1_0_n53 )  ;
assign n27383 =  ( wr_addr ) == ( bv_8_233_n535 )  ;
assign n27384 =  ( n27382 ) & (n27383 )  ;
assign n27385 =  ( n27384 ) & (wr )  ;
assign n27386 =  ( n27385 ) ? ( n5325 ) : ( iram_233 ) ;
assign n27387 = wr_addr[7:7] ;
assign n27388 =  ( n27387 ) == ( bv_1_0_n53 )  ;
assign n27389 =  ( wr_addr ) == ( bv_8_234_n537 )  ;
assign n27390 =  ( n27388 ) & (n27389 )  ;
assign n27391 =  ( n27390 ) & (wr )  ;
assign n27392 =  ( n27391 ) ? ( n4782 ) : ( iram_234 ) ;
assign n27393 = wr_addr[7:7] ;
assign n27394 =  ( n27393 ) == ( bv_1_0_n53 )  ;
assign n27395 =  ( wr_addr ) == ( bv_8_234_n537 )  ;
assign n27396 =  ( n27394 ) & (n27395 )  ;
assign n27397 =  ( n27396 ) & (wr )  ;
assign n27398 =  ( n27397 ) ? ( n4841 ) : ( iram_234 ) ;
assign n27399 = wr_addr[7:7] ;
assign n27400 =  ( n27399 ) == ( bv_1_0_n53 )  ;
assign n27401 =  ( wr_addr ) == ( bv_8_234_n537 )  ;
assign n27402 =  ( n27400 ) & (n27401 )  ;
assign n27403 =  ( n27402 ) & (wr )  ;
assign n27404 =  ( n27403 ) ? ( n5449 ) : ( iram_234 ) ;
assign n27405 = wr_addr[7:7] ;
assign n27406 =  ( n27405 ) == ( bv_1_0_n53 )  ;
assign n27407 =  ( wr_addr ) == ( bv_8_234_n537 )  ;
assign n27408 =  ( n27406 ) & (n27407 )  ;
assign n27409 =  ( n27408 ) & (wr )  ;
assign n27410 =  ( n27409 ) ? ( n4906 ) : ( iram_234 ) ;
assign n27411 = wr_addr[7:7] ;
assign n27412 =  ( n27411 ) == ( bv_1_0_n53 )  ;
assign n27413 =  ( wr_addr ) == ( bv_8_234_n537 )  ;
assign n27414 =  ( n27412 ) & (n27413 )  ;
assign n27415 =  ( n27414 ) & (wr )  ;
assign n27416 =  ( n27415 ) ? ( n5485 ) : ( iram_234 ) ;
assign n27417 = wr_addr[7:7] ;
assign n27418 =  ( n27417 ) == ( bv_1_0_n53 )  ;
assign n27419 =  ( wr_addr ) == ( bv_8_234_n537 )  ;
assign n27420 =  ( n27418 ) & (n27419 )  ;
assign n27421 =  ( n27420 ) & (wr )  ;
assign n27422 =  ( n27421 ) ? ( n5512 ) : ( iram_234 ) ;
assign n27423 = wr_addr[7:7] ;
assign n27424 =  ( n27423 ) == ( bv_1_0_n53 )  ;
assign n27425 =  ( wr_addr ) == ( bv_8_234_n537 )  ;
assign n27426 =  ( n27424 ) & (n27425 )  ;
assign n27427 =  ( n27426 ) & (wr )  ;
assign n27428 =  ( n27427 ) ? ( bv_8_0_n69 ) : ( iram_234 ) ;
assign n27429 = wr_addr[7:7] ;
assign n27430 =  ( n27429 ) == ( bv_1_0_n53 )  ;
assign n27431 =  ( wr_addr ) == ( bv_8_234_n537 )  ;
assign n27432 =  ( n27430 ) & (n27431 )  ;
assign n27433 =  ( n27432 ) & (wr )  ;
assign n27434 =  ( n27433 ) ? ( n5071 ) : ( iram_234 ) ;
assign n27435 = wr_addr[7:7] ;
assign n27436 =  ( n27435 ) == ( bv_1_0_n53 )  ;
assign n27437 =  ( wr_addr ) == ( bv_8_234_n537 )  ;
assign n27438 =  ( n27436 ) & (n27437 )  ;
assign n27439 =  ( n27438 ) & (wr )  ;
assign n27440 =  ( n27439 ) ? ( n5096 ) : ( iram_234 ) ;
assign n27441 = wr_addr[7:7] ;
assign n27442 =  ( n27441 ) == ( bv_1_0_n53 )  ;
assign n27443 =  ( wr_addr ) == ( bv_8_234_n537 )  ;
assign n27444 =  ( n27442 ) & (n27443 )  ;
assign n27445 =  ( n27444 ) & (wr )  ;
assign n27446 =  ( n27445 ) ? ( n5123 ) : ( iram_234 ) ;
assign n27447 = wr_addr[7:7] ;
assign n27448 =  ( n27447 ) == ( bv_1_0_n53 )  ;
assign n27449 =  ( wr_addr ) == ( bv_8_234_n537 )  ;
assign n27450 =  ( n27448 ) & (n27449 )  ;
assign n27451 =  ( n27450 ) & (wr )  ;
assign n27452 =  ( n27451 ) ? ( n5165 ) : ( iram_234 ) ;
assign n27453 = wr_addr[7:7] ;
assign n27454 =  ( n27453 ) == ( bv_1_0_n53 )  ;
assign n27455 =  ( wr_addr ) == ( bv_8_234_n537 )  ;
assign n27456 =  ( n27454 ) & (n27455 )  ;
assign n27457 =  ( n27456 ) & (wr )  ;
assign n27458 =  ( n27457 ) ? ( n5204 ) : ( iram_234 ) ;
assign n27459 = wr_addr[7:7] ;
assign n27460 =  ( n27459 ) == ( bv_1_0_n53 )  ;
assign n27461 =  ( wr_addr ) == ( bv_8_234_n537 )  ;
assign n27462 =  ( n27460 ) & (n27461 )  ;
assign n27463 =  ( n27462 ) & (wr )  ;
assign n27464 =  ( n27463 ) ? ( n5262 ) : ( iram_234 ) ;
assign n27465 = wr_addr[7:7] ;
assign n27466 =  ( n27465 ) == ( bv_1_0_n53 )  ;
assign n27467 =  ( wr_addr ) == ( bv_8_234_n537 )  ;
assign n27468 =  ( n27466 ) & (n27467 )  ;
assign n27469 =  ( n27468 ) & (wr )  ;
assign n27470 =  ( n27469 ) ? ( n5298 ) : ( iram_234 ) ;
assign n27471 = wr_addr[7:7] ;
assign n27472 =  ( n27471 ) == ( bv_1_0_n53 )  ;
assign n27473 =  ( wr_addr ) == ( bv_8_234_n537 )  ;
assign n27474 =  ( n27472 ) & (n27473 )  ;
assign n27475 =  ( n27474 ) & (wr )  ;
assign n27476 =  ( n27475 ) ? ( n5325 ) : ( iram_234 ) ;
assign n27477 = wr_addr[7:7] ;
assign n27478 =  ( n27477 ) == ( bv_1_0_n53 )  ;
assign n27479 =  ( wr_addr ) == ( bv_8_235_n539 )  ;
assign n27480 =  ( n27478 ) & (n27479 )  ;
assign n27481 =  ( n27480 ) & (wr )  ;
assign n27482 =  ( n27481 ) ? ( n4782 ) : ( iram_235 ) ;
assign n27483 = wr_addr[7:7] ;
assign n27484 =  ( n27483 ) == ( bv_1_0_n53 )  ;
assign n27485 =  ( wr_addr ) == ( bv_8_235_n539 )  ;
assign n27486 =  ( n27484 ) & (n27485 )  ;
assign n27487 =  ( n27486 ) & (wr )  ;
assign n27488 =  ( n27487 ) ? ( n4841 ) : ( iram_235 ) ;
assign n27489 = wr_addr[7:7] ;
assign n27490 =  ( n27489 ) == ( bv_1_0_n53 )  ;
assign n27491 =  ( wr_addr ) == ( bv_8_235_n539 )  ;
assign n27492 =  ( n27490 ) & (n27491 )  ;
assign n27493 =  ( n27492 ) & (wr )  ;
assign n27494 =  ( n27493 ) ? ( n5449 ) : ( iram_235 ) ;
assign n27495 = wr_addr[7:7] ;
assign n27496 =  ( n27495 ) == ( bv_1_0_n53 )  ;
assign n27497 =  ( wr_addr ) == ( bv_8_235_n539 )  ;
assign n27498 =  ( n27496 ) & (n27497 )  ;
assign n27499 =  ( n27498 ) & (wr )  ;
assign n27500 =  ( n27499 ) ? ( n4906 ) : ( iram_235 ) ;
assign n27501 = wr_addr[7:7] ;
assign n27502 =  ( n27501 ) == ( bv_1_0_n53 )  ;
assign n27503 =  ( wr_addr ) == ( bv_8_235_n539 )  ;
assign n27504 =  ( n27502 ) & (n27503 )  ;
assign n27505 =  ( n27504 ) & (wr )  ;
assign n27506 =  ( n27505 ) ? ( n5485 ) : ( iram_235 ) ;
assign n27507 = wr_addr[7:7] ;
assign n27508 =  ( n27507 ) == ( bv_1_0_n53 )  ;
assign n27509 =  ( wr_addr ) == ( bv_8_235_n539 )  ;
assign n27510 =  ( n27508 ) & (n27509 )  ;
assign n27511 =  ( n27510 ) & (wr )  ;
assign n27512 =  ( n27511 ) ? ( n5512 ) : ( iram_235 ) ;
assign n27513 = wr_addr[7:7] ;
assign n27514 =  ( n27513 ) == ( bv_1_0_n53 )  ;
assign n27515 =  ( wr_addr ) == ( bv_8_235_n539 )  ;
assign n27516 =  ( n27514 ) & (n27515 )  ;
assign n27517 =  ( n27516 ) & (wr )  ;
assign n27518 =  ( n27517 ) ? ( bv_8_0_n69 ) : ( iram_235 ) ;
assign n27519 = wr_addr[7:7] ;
assign n27520 =  ( n27519 ) == ( bv_1_0_n53 )  ;
assign n27521 =  ( wr_addr ) == ( bv_8_235_n539 )  ;
assign n27522 =  ( n27520 ) & (n27521 )  ;
assign n27523 =  ( n27522 ) & (wr )  ;
assign n27524 =  ( n27523 ) ? ( n5071 ) : ( iram_235 ) ;
assign n27525 = wr_addr[7:7] ;
assign n27526 =  ( n27525 ) == ( bv_1_0_n53 )  ;
assign n27527 =  ( wr_addr ) == ( bv_8_235_n539 )  ;
assign n27528 =  ( n27526 ) & (n27527 )  ;
assign n27529 =  ( n27528 ) & (wr )  ;
assign n27530 =  ( n27529 ) ? ( n5096 ) : ( iram_235 ) ;
assign n27531 = wr_addr[7:7] ;
assign n27532 =  ( n27531 ) == ( bv_1_0_n53 )  ;
assign n27533 =  ( wr_addr ) == ( bv_8_235_n539 )  ;
assign n27534 =  ( n27532 ) & (n27533 )  ;
assign n27535 =  ( n27534 ) & (wr )  ;
assign n27536 =  ( n27535 ) ? ( n5123 ) : ( iram_235 ) ;
assign n27537 = wr_addr[7:7] ;
assign n27538 =  ( n27537 ) == ( bv_1_0_n53 )  ;
assign n27539 =  ( wr_addr ) == ( bv_8_235_n539 )  ;
assign n27540 =  ( n27538 ) & (n27539 )  ;
assign n27541 =  ( n27540 ) & (wr )  ;
assign n27542 =  ( n27541 ) ? ( n5165 ) : ( iram_235 ) ;
assign n27543 = wr_addr[7:7] ;
assign n27544 =  ( n27543 ) == ( bv_1_0_n53 )  ;
assign n27545 =  ( wr_addr ) == ( bv_8_235_n539 )  ;
assign n27546 =  ( n27544 ) & (n27545 )  ;
assign n27547 =  ( n27546 ) & (wr )  ;
assign n27548 =  ( n27547 ) ? ( n5204 ) : ( iram_235 ) ;
assign n27549 = wr_addr[7:7] ;
assign n27550 =  ( n27549 ) == ( bv_1_0_n53 )  ;
assign n27551 =  ( wr_addr ) == ( bv_8_235_n539 )  ;
assign n27552 =  ( n27550 ) & (n27551 )  ;
assign n27553 =  ( n27552 ) & (wr )  ;
assign n27554 =  ( n27553 ) ? ( n5262 ) : ( iram_235 ) ;
assign n27555 = wr_addr[7:7] ;
assign n27556 =  ( n27555 ) == ( bv_1_0_n53 )  ;
assign n27557 =  ( wr_addr ) == ( bv_8_235_n539 )  ;
assign n27558 =  ( n27556 ) & (n27557 )  ;
assign n27559 =  ( n27558 ) & (wr )  ;
assign n27560 =  ( n27559 ) ? ( n5298 ) : ( iram_235 ) ;
assign n27561 = wr_addr[7:7] ;
assign n27562 =  ( n27561 ) == ( bv_1_0_n53 )  ;
assign n27563 =  ( wr_addr ) == ( bv_8_235_n539 )  ;
assign n27564 =  ( n27562 ) & (n27563 )  ;
assign n27565 =  ( n27564 ) & (wr )  ;
assign n27566 =  ( n27565 ) ? ( n5325 ) : ( iram_235 ) ;
assign n27567 = wr_addr[7:7] ;
assign n27568 =  ( n27567 ) == ( bv_1_0_n53 )  ;
assign n27569 =  ( wr_addr ) == ( bv_8_236_n541 )  ;
assign n27570 =  ( n27568 ) & (n27569 )  ;
assign n27571 =  ( n27570 ) & (wr )  ;
assign n27572 =  ( n27571 ) ? ( n4782 ) : ( iram_236 ) ;
assign n27573 = wr_addr[7:7] ;
assign n27574 =  ( n27573 ) == ( bv_1_0_n53 )  ;
assign n27575 =  ( wr_addr ) == ( bv_8_236_n541 )  ;
assign n27576 =  ( n27574 ) & (n27575 )  ;
assign n27577 =  ( n27576 ) & (wr )  ;
assign n27578 =  ( n27577 ) ? ( n4841 ) : ( iram_236 ) ;
assign n27579 = wr_addr[7:7] ;
assign n27580 =  ( n27579 ) == ( bv_1_0_n53 )  ;
assign n27581 =  ( wr_addr ) == ( bv_8_236_n541 )  ;
assign n27582 =  ( n27580 ) & (n27581 )  ;
assign n27583 =  ( n27582 ) & (wr )  ;
assign n27584 =  ( n27583 ) ? ( n5449 ) : ( iram_236 ) ;
assign n27585 = wr_addr[7:7] ;
assign n27586 =  ( n27585 ) == ( bv_1_0_n53 )  ;
assign n27587 =  ( wr_addr ) == ( bv_8_236_n541 )  ;
assign n27588 =  ( n27586 ) & (n27587 )  ;
assign n27589 =  ( n27588 ) & (wr )  ;
assign n27590 =  ( n27589 ) ? ( n4906 ) : ( iram_236 ) ;
assign n27591 = wr_addr[7:7] ;
assign n27592 =  ( n27591 ) == ( bv_1_0_n53 )  ;
assign n27593 =  ( wr_addr ) == ( bv_8_236_n541 )  ;
assign n27594 =  ( n27592 ) & (n27593 )  ;
assign n27595 =  ( n27594 ) & (wr )  ;
assign n27596 =  ( n27595 ) ? ( n5485 ) : ( iram_236 ) ;
assign n27597 = wr_addr[7:7] ;
assign n27598 =  ( n27597 ) == ( bv_1_0_n53 )  ;
assign n27599 =  ( wr_addr ) == ( bv_8_236_n541 )  ;
assign n27600 =  ( n27598 ) & (n27599 )  ;
assign n27601 =  ( n27600 ) & (wr )  ;
assign n27602 =  ( n27601 ) ? ( n5512 ) : ( iram_236 ) ;
assign n27603 = wr_addr[7:7] ;
assign n27604 =  ( n27603 ) == ( bv_1_0_n53 )  ;
assign n27605 =  ( wr_addr ) == ( bv_8_236_n541 )  ;
assign n27606 =  ( n27604 ) & (n27605 )  ;
assign n27607 =  ( n27606 ) & (wr )  ;
assign n27608 =  ( n27607 ) ? ( bv_8_0_n69 ) : ( iram_236 ) ;
assign n27609 = wr_addr[7:7] ;
assign n27610 =  ( n27609 ) == ( bv_1_0_n53 )  ;
assign n27611 =  ( wr_addr ) == ( bv_8_236_n541 )  ;
assign n27612 =  ( n27610 ) & (n27611 )  ;
assign n27613 =  ( n27612 ) & (wr )  ;
assign n27614 =  ( n27613 ) ? ( n5071 ) : ( iram_236 ) ;
assign n27615 = wr_addr[7:7] ;
assign n27616 =  ( n27615 ) == ( bv_1_0_n53 )  ;
assign n27617 =  ( wr_addr ) == ( bv_8_236_n541 )  ;
assign n27618 =  ( n27616 ) & (n27617 )  ;
assign n27619 =  ( n27618 ) & (wr )  ;
assign n27620 =  ( n27619 ) ? ( n5096 ) : ( iram_236 ) ;
assign n27621 = wr_addr[7:7] ;
assign n27622 =  ( n27621 ) == ( bv_1_0_n53 )  ;
assign n27623 =  ( wr_addr ) == ( bv_8_236_n541 )  ;
assign n27624 =  ( n27622 ) & (n27623 )  ;
assign n27625 =  ( n27624 ) & (wr )  ;
assign n27626 =  ( n27625 ) ? ( n5123 ) : ( iram_236 ) ;
assign n27627 = wr_addr[7:7] ;
assign n27628 =  ( n27627 ) == ( bv_1_0_n53 )  ;
assign n27629 =  ( wr_addr ) == ( bv_8_236_n541 )  ;
assign n27630 =  ( n27628 ) & (n27629 )  ;
assign n27631 =  ( n27630 ) & (wr )  ;
assign n27632 =  ( n27631 ) ? ( n5165 ) : ( iram_236 ) ;
assign n27633 = wr_addr[7:7] ;
assign n27634 =  ( n27633 ) == ( bv_1_0_n53 )  ;
assign n27635 =  ( wr_addr ) == ( bv_8_236_n541 )  ;
assign n27636 =  ( n27634 ) & (n27635 )  ;
assign n27637 =  ( n27636 ) & (wr )  ;
assign n27638 =  ( n27637 ) ? ( n5204 ) : ( iram_236 ) ;
assign n27639 = wr_addr[7:7] ;
assign n27640 =  ( n27639 ) == ( bv_1_0_n53 )  ;
assign n27641 =  ( wr_addr ) == ( bv_8_236_n541 )  ;
assign n27642 =  ( n27640 ) & (n27641 )  ;
assign n27643 =  ( n27642 ) & (wr )  ;
assign n27644 =  ( n27643 ) ? ( n5262 ) : ( iram_236 ) ;
assign n27645 = wr_addr[7:7] ;
assign n27646 =  ( n27645 ) == ( bv_1_0_n53 )  ;
assign n27647 =  ( wr_addr ) == ( bv_8_236_n541 )  ;
assign n27648 =  ( n27646 ) & (n27647 )  ;
assign n27649 =  ( n27648 ) & (wr )  ;
assign n27650 =  ( n27649 ) ? ( n5298 ) : ( iram_236 ) ;
assign n27651 = wr_addr[7:7] ;
assign n27652 =  ( n27651 ) == ( bv_1_0_n53 )  ;
assign n27653 =  ( wr_addr ) == ( bv_8_236_n541 )  ;
assign n27654 =  ( n27652 ) & (n27653 )  ;
assign n27655 =  ( n27654 ) & (wr )  ;
assign n27656 =  ( n27655 ) ? ( n5325 ) : ( iram_236 ) ;
assign n27657 = wr_addr[7:7] ;
assign n27658 =  ( n27657 ) == ( bv_1_0_n53 )  ;
assign n27659 =  ( wr_addr ) == ( bv_8_237_n543 )  ;
assign n27660 =  ( n27658 ) & (n27659 )  ;
assign n27661 =  ( n27660 ) & (wr )  ;
assign n27662 =  ( n27661 ) ? ( n4782 ) : ( iram_237 ) ;
assign n27663 = wr_addr[7:7] ;
assign n27664 =  ( n27663 ) == ( bv_1_0_n53 )  ;
assign n27665 =  ( wr_addr ) == ( bv_8_237_n543 )  ;
assign n27666 =  ( n27664 ) & (n27665 )  ;
assign n27667 =  ( n27666 ) & (wr )  ;
assign n27668 =  ( n27667 ) ? ( n4841 ) : ( iram_237 ) ;
assign n27669 = wr_addr[7:7] ;
assign n27670 =  ( n27669 ) == ( bv_1_0_n53 )  ;
assign n27671 =  ( wr_addr ) == ( bv_8_237_n543 )  ;
assign n27672 =  ( n27670 ) & (n27671 )  ;
assign n27673 =  ( n27672 ) & (wr )  ;
assign n27674 =  ( n27673 ) ? ( n5449 ) : ( iram_237 ) ;
assign n27675 = wr_addr[7:7] ;
assign n27676 =  ( n27675 ) == ( bv_1_0_n53 )  ;
assign n27677 =  ( wr_addr ) == ( bv_8_237_n543 )  ;
assign n27678 =  ( n27676 ) & (n27677 )  ;
assign n27679 =  ( n27678 ) & (wr )  ;
assign n27680 =  ( n27679 ) ? ( n4906 ) : ( iram_237 ) ;
assign n27681 = wr_addr[7:7] ;
assign n27682 =  ( n27681 ) == ( bv_1_0_n53 )  ;
assign n27683 =  ( wr_addr ) == ( bv_8_237_n543 )  ;
assign n27684 =  ( n27682 ) & (n27683 )  ;
assign n27685 =  ( n27684 ) & (wr )  ;
assign n27686 =  ( n27685 ) ? ( n5485 ) : ( iram_237 ) ;
assign n27687 = wr_addr[7:7] ;
assign n27688 =  ( n27687 ) == ( bv_1_0_n53 )  ;
assign n27689 =  ( wr_addr ) == ( bv_8_237_n543 )  ;
assign n27690 =  ( n27688 ) & (n27689 )  ;
assign n27691 =  ( n27690 ) & (wr )  ;
assign n27692 =  ( n27691 ) ? ( n5512 ) : ( iram_237 ) ;
assign n27693 = wr_addr[7:7] ;
assign n27694 =  ( n27693 ) == ( bv_1_0_n53 )  ;
assign n27695 =  ( wr_addr ) == ( bv_8_237_n543 )  ;
assign n27696 =  ( n27694 ) & (n27695 )  ;
assign n27697 =  ( n27696 ) & (wr )  ;
assign n27698 =  ( n27697 ) ? ( bv_8_0_n69 ) : ( iram_237 ) ;
assign n27699 = wr_addr[7:7] ;
assign n27700 =  ( n27699 ) == ( bv_1_0_n53 )  ;
assign n27701 =  ( wr_addr ) == ( bv_8_237_n543 )  ;
assign n27702 =  ( n27700 ) & (n27701 )  ;
assign n27703 =  ( n27702 ) & (wr )  ;
assign n27704 =  ( n27703 ) ? ( n5071 ) : ( iram_237 ) ;
assign n27705 = wr_addr[7:7] ;
assign n27706 =  ( n27705 ) == ( bv_1_0_n53 )  ;
assign n27707 =  ( wr_addr ) == ( bv_8_237_n543 )  ;
assign n27708 =  ( n27706 ) & (n27707 )  ;
assign n27709 =  ( n27708 ) & (wr )  ;
assign n27710 =  ( n27709 ) ? ( n5096 ) : ( iram_237 ) ;
assign n27711 = wr_addr[7:7] ;
assign n27712 =  ( n27711 ) == ( bv_1_0_n53 )  ;
assign n27713 =  ( wr_addr ) == ( bv_8_237_n543 )  ;
assign n27714 =  ( n27712 ) & (n27713 )  ;
assign n27715 =  ( n27714 ) & (wr )  ;
assign n27716 =  ( n27715 ) ? ( n5123 ) : ( iram_237 ) ;
assign n27717 = wr_addr[7:7] ;
assign n27718 =  ( n27717 ) == ( bv_1_0_n53 )  ;
assign n27719 =  ( wr_addr ) == ( bv_8_237_n543 )  ;
assign n27720 =  ( n27718 ) & (n27719 )  ;
assign n27721 =  ( n27720 ) & (wr )  ;
assign n27722 =  ( n27721 ) ? ( n5165 ) : ( iram_237 ) ;
assign n27723 = wr_addr[7:7] ;
assign n27724 =  ( n27723 ) == ( bv_1_0_n53 )  ;
assign n27725 =  ( wr_addr ) == ( bv_8_237_n543 )  ;
assign n27726 =  ( n27724 ) & (n27725 )  ;
assign n27727 =  ( n27726 ) & (wr )  ;
assign n27728 =  ( n27727 ) ? ( n5204 ) : ( iram_237 ) ;
assign n27729 = wr_addr[7:7] ;
assign n27730 =  ( n27729 ) == ( bv_1_0_n53 )  ;
assign n27731 =  ( wr_addr ) == ( bv_8_237_n543 )  ;
assign n27732 =  ( n27730 ) & (n27731 )  ;
assign n27733 =  ( n27732 ) & (wr )  ;
assign n27734 =  ( n27733 ) ? ( n5262 ) : ( iram_237 ) ;
assign n27735 = wr_addr[7:7] ;
assign n27736 =  ( n27735 ) == ( bv_1_0_n53 )  ;
assign n27737 =  ( wr_addr ) == ( bv_8_237_n543 )  ;
assign n27738 =  ( n27736 ) & (n27737 )  ;
assign n27739 =  ( n27738 ) & (wr )  ;
assign n27740 =  ( n27739 ) ? ( n5298 ) : ( iram_237 ) ;
assign n27741 = wr_addr[7:7] ;
assign n27742 =  ( n27741 ) == ( bv_1_0_n53 )  ;
assign n27743 =  ( wr_addr ) == ( bv_8_237_n543 )  ;
assign n27744 =  ( n27742 ) & (n27743 )  ;
assign n27745 =  ( n27744 ) & (wr )  ;
assign n27746 =  ( n27745 ) ? ( n5325 ) : ( iram_237 ) ;
assign n27747 = wr_addr[7:7] ;
assign n27748 =  ( n27747 ) == ( bv_1_0_n53 )  ;
assign n27749 =  ( wr_addr ) == ( bv_8_238_n545 )  ;
assign n27750 =  ( n27748 ) & (n27749 )  ;
assign n27751 =  ( n27750 ) & (wr )  ;
assign n27752 =  ( n27751 ) ? ( n4782 ) : ( iram_238 ) ;
assign n27753 = wr_addr[7:7] ;
assign n27754 =  ( n27753 ) == ( bv_1_0_n53 )  ;
assign n27755 =  ( wr_addr ) == ( bv_8_238_n545 )  ;
assign n27756 =  ( n27754 ) & (n27755 )  ;
assign n27757 =  ( n27756 ) & (wr )  ;
assign n27758 =  ( n27757 ) ? ( n4841 ) : ( iram_238 ) ;
assign n27759 = wr_addr[7:7] ;
assign n27760 =  ( n27759 ) == ( bv_1_0_n53 )  ;
assign n27761 =  ( wr_addr ) == ( bv_8_238_n545 )  ;
assign n27762 =  ( n27760 ) & (n27761 )  ;
assign n27763 =  ( n27762 ) & (wr )  ;
assign n27764 =  ( n27763 ) ? ( n5449 ) : ( iram_238 ) ;
assign n27765 = wr_addr[7:7] ;
assign n27766 =  ( n27765 ) == ( bv_1_0_n53 )  ;
assign n27767 =  ( wr_addr ) == ( bv_8_238_n545 )  ;
assign n27768 =  ( n27766 ) & (n27767 )  ;
assign n27769 =  ( n27768 ) & (wr )  ;
assign n27770 =  ( n27769 ) ? ( n4906 ) : ( iram_238 ) ;
assign n27771 = wr_addr[7:7] ;
assign n27772 =  ( n27771 ) == ( bv_1_0_n53 )  ;
assign n27773 =  ( wr_addr ) == ( bv_8_238_n545 )  ;
assign n27774 =  ( n27772 ) & (n27773 )  ;
assign n27775 =  ( n27774 ) & (wr )  ;
assign n27776 =  ( n27775 ) ? ( n5485 ) : ( iram_238 ) ;
assign n27777 = wr_addr[7:7] ;
assign n27778 =  ( n27777 ) == ( bv_1_0_n53 )  ;
assign n27779 =  ( wr_addr ) == ( bv_8_238_n545 )  ;
assign n27780 =  ( n27778 ) & (n27779 )  ;
assign n27781 =  ( n27780 ) & (wr )  ;
assign n27782 =  ( n27781 ) ? ( n5512 ) : ( iram_238 ) ;
assign n27783 = wr_addr[7:7] ;
assign n27784 =  ( n27783 ) == ( bv_1_0_n53 )  ;
assign n27785 =  ( wr_addr ) == ( bv_8_238_n545 )  ;
assign n27786 =  ( n27784 ) & (n27785 )  ;
assign n27787 =  ( n27786 ) & (wr )  ;
assign n27788 =  ( n27787 ) ? ( bv_8_0_n69 ) : ( iram_238 ) ;
assign n27789 = wr_addr[7:7] ;
assign n27790 =  ( n27789 ) == ( bv_1_0_n53 )  ;
assign n27791 =  ( wr_addr ) == ( bv_8_238_n545 )  ;
assign n27792 =  ( n27790 ) & (n27791 )  ;
assign n27793 =  ( n27792 ) & (wr )  ;
assign n27794 =  ( n27793 ) ? ( n5071 ) : ( iram_238 ) ;
assign n27795 = wr_addr[7:7] ;
assign n27796 =  ( n27795 ) == ( bv_1_0_n53 )  ;
assign n27797 =  ( wr_addr ) == ( bv_8_238_n545 )  ;
assign n27798 =  ( n27796 ) & (n27797 )  ;
assign n27799 =  ( n27798 ) & (wr )  ;
assign n27800 =  ( n27799 ) ? ( n5096 ) : ( iram_238 ) ;
assign n27801 = wr_addr[7:7] ;
assign n27802 =  ( n27801 ) == ( bv_1_0_n53 )  ;
assign n27803 =  ( wr_addr ) == ( bv_8_238_n545 )  ;
assign n27804 =  ( n27802 ) & (n27803 )  ;
assign n27805 =  ( n27804 ) & (wr )  ;
assign n27806 =  ( n27805 ) ? ( n5123 ) : ( iram_238 ) ;
assign n27807 = wr_addr[7:7] ;
assign n27808 =  ( n27807 ) == ( bv_1_0_n53 )  ;
assign n27809 =  ( wr_addr ) == ( bv_8_238_n545 )  ;
assign n27810 =  ( n27808 ) & (n27809 )  ;
assign n27811 =  ( n27810 ) & (wr )  ;
assign n27812 =  ( n27811 ) ? ( n5165 ) : ( iram_238 ) ;
assign n27813 = wr_addr[7:7] ;
assign n27814 =  ( n27813 ) == ( bv_1_0_n53 )  ;
assign n27815 =  ( wr_addr ) == ( bv_8_238_n545 )  ;
assign n27816 =  ( n27814 ) & (n27815 )  ;
assign n27817 =  ( n27816 ) & (wr )  ;
assign n27818 =  ( n27817 ) ? ( n5204 ) : ( iram_238 ) ;
assign n27819 = wr_addr[7:7] ;
assign n27820 =  ( n27819 ) == ( bv_1_0_n53 )  ;
assign n27821 =  ( wr_addr ) == ( bv_8_238_n545 )  ;
assign n27822 =  ( n27820 ) & (n27821 )  ;
assign n27823 =  ( n27822 ) & (wr )  ;
assign n27824 =  ( n27823 ) ? ( n5262 ) : ( iram_238 ) ;
assign n27825 = wr_addr[7:7] ;
assign n27826 =  ( n27825 ) == ( bv_1_0_n53 )  ;
assign n27827 =  ( wr_addr ) == ( bv_8_238_n545 )  ;
assign n27828 =  ( n27826 ) & (n27827 )  ;
assign n27829 =  ( n27828 ) & (wr )  ;
assign n27830 =  ( n27829 ) ? ( n5298 ) : ( iram_238 ) ;
assign n27831 = wr_addr[7:7] ;
assign n27832 =  ( n27831 ) == ( bv_1_0_n53 )  ;
assign n27833 =  ( wr_addr ) == ( bv_8_238_n545 )  ;
assign n27834 =  ( n27832 ) & (n27833 )  ;
assign n27835 =  ( n27834 ) & (wr )  ;
assign n27836 =  ( n27835 ) ? ( n5325 ) : ( iram_238 ) ;
assign n27837 = wr_addr[7:7] ;
assign n27838 =  ( n27837 ) == ( bv_1_0_n53 )  ;
assign n27839 =  ( wr_addr ) == ( bv_8_239_n547 )  ;
assign n27840 =  ( n27838 ) & (n27839 )  ;
assign n27841 =  ( n27840 ) & (wr )  ;
assign n27842 =  ( n27841 ) ? ( n4782 ) : ( iram_239 ) ;
assign n27843 = wr_addr[7:7] ;
assign n27844 =  ( n27843 ) == ( bv_1_0_n53 )  ;
assign n27845 =  ( wr_addr ) == ( bv_8_239_n547 )  ;
assign n27846 =  ( n27844 ) & (n27845 )  ;
assign n27847 =  ( n27846 ) & (wr )  ;
assign n27848 =  ( n27847 ) ? ( n4841 ) : ( iram_239 ) ;
assign n27849 = wr_addr[7:7] ;
assign n27850 =  ( n27849 ) == ( bv_1_0_n53 )  ;
assign n27851 =  ( wr_addr ) == ( bv_8_239_n547 )  ;
assign n27852 =  ( n27850 ) & (n27851 )  ;
assign n27853 =  ( n27852 ) & (wr )  ;
assign n27854 =  ( n27853 ) ? ( n5449 ) : ( iram_239 ) ;
assign n27855 = wr_addr[7:7] ;
assign n27856 =  ( n27855 ) == ( bv_1_0_n53 )  ;
assign n27857 =  ( wr_addr ) == ( bv_8_239_n547 )  ;
assign n27858 =  ( n27856 ) & (n27857 )  ;
assign n27859 =  ( n27858 ) & (wr )  ;
assign n27860 =  ( n27859 ) ? ( n4906 ) : ( iram_239 ) ;
assign n27861 = wr_addr[7:7] ;
assign n27862 =  ( n27861 ) == ( bv_1_0_n53 )  ;
assign n27863 =  ( wr_addr ) == ( bv_8_239_n547 )  ;
assign n27864 =  ( n27862 ) & (n27863 )  ;
assign n27865 =  ( n27864 ) & (wr )  ;
assign n27866 =  ( n27865 ) ? ( n5485 ) : ( iram_239 ) ;
assign n27867 = wr_addr[7:7] ;
assign n27868 =  ( n27867 ) == ( bv_1_0_n53 )  ;
assign n27869 =  ( wr_addr ) == ( bv_8_239_n547 )  ;
assign n27870 =  ( n27868 ) & (n27869 )  ;
assign n27871 =  ( n27870 ) & (wr )  ;
assign n27872 =  ( n27871 ) ? ( n5512 ) : ( iram_239 ) ;
assign n27873 = wr_addr[7:7] ;
assign n27874 =  ( n27873 ) == ( bv_1_0_n53 )  ;
assign n27875 =  ( wr_addr ) == ( bv_8_239_n547 )  ;
assign n27876 =  ( n27874 ) & (n27875 )  ;
assign n27877 =  ( n27876 ) & (wr )  ;
assign n27878 =  ( n27877 ) ? ( bv_8_0_n69 ) : ( iram_239 ) ;
assign n27879 = wr_addr[7:7] ;
assign n27880 =  ( n27879 ) == ( bv_1_0_n53 )  ;
assign n27881 =  ( wr_addr ) == ( bv_8_239_n547 )  ;
assign n27882 =  ( n27880 ) & (n27881 )  ;
assign n27883 =  ( n27882 ) & (wr )  ;
assign n27884 =  ( n27883 ) ? ( n5071 ) : ( iram_239 ) ;
assign n27885 = wr_addr[7:7] ;
assign n27886 =  ( n27885 ) == ( bv_1_0_n53 )  ;
assign n27887 =  ( wr_addr ) == ( bv_8_239_n547 )  ;
assign n27888 =  ( n27886 ) & (n27887 )  ;
assign n27889 =  ( n27888 ) & (wr )  ;
assign n27890 =  ( n27889 ) ? ( n5096 ) : ( iram_239 ) ;
assign n27891 = wr_addr[7:7] ;
assign n27892 =  ( n27891 ) == ( bv_1_0_n53 )  ;
assign n27893 =  ( wr_addr ) == ( bv_8_239_n547 )  ;
assign n27894 =  ( n27892 ) & (n27893 )  ;
assign n27895 =  ( n27894 ) & (wr )  ;
assign n27896 =  ( n27895 ) ? ( n5123 ) : ( iram_239 ) ;
assign n27897 = wr_addr[7:7] ;
assign n27898 =  ( n27897 ) == ( bv_1_0_n53 )  ;
assign n27899 =  ( wr_addr ) == ( bv_8_239_n547 )  ;
assign n27900 =  ( n27898 ) & (n27899 )  ;
assign n27901 =  ( n27900 ) & (wr )  ;
assign n27902 =  ( n27901 ) ? ( n5165 ) : ( iram_239 ) ;
assign n27903 = wr_addr[7:7] ;
assign n27904 =  ( n27903 ) == ( bv_1_0_n53 )  ;
assign n27905 =  ( wr_addr ) == ( bv_8_239_n547 )  ;
assign n27906 =  ( n27904 ) & (n27905 )  ;
assign n27907 =  ( n27906 ) & (wr )  ;
assign n27908 =  ( n27907 ) ? ( n5204 ) : ( iram_239 ) ;
assign n27909 = wr_addr[7:7] ;
assign n27910 =  ( n27909 ) == ( bv_1_0_n53 )  ;
assign n27911 =  ( wr_addr ) == ( bv_8_239_n547 )  ;
assign n27912 =  ( n27910 ) & (n27911 )  ;
assign n27913 =  ( n27912 ) & (wr )  ;
assign n27914 =  ( n27913 ) ? ( n5262 ) : ( iram_239 ) ;
assign n27915 = wr_addr[7:7] ;
assign n27916 =  ( n27915 ) == ( bv_1_0_n53 )  ;
assign n27917 =  ( wr_addr ) == ( bv_8_239_n547 )  ;
assign n27918 =  ( n27916 ) & (n27917 )  ;
assign n27919 =  ( n27918 ) & (wr )  ;
assign n27920 =  ( n27919 ) ? ( n5298 ) : ( iram_239 ) ;
assign n27921 = wr_addr[7:7] ;
assign n27922 =  ( n27921 ) == ( bv_1_0_n53 )  ;
assign n27923 =  ( wr_addr ) == ( bv_8_239_n547 )  ;
assign n27924 =  ( n27922 ) & (n27923 )  ;
assign n27925 =  ( n27924 ) & (wr )  ;
assign n27926 =  ( n27925 ) ? ( n5325 ) : ( iram_239 ) ;
assign n27927 = wr_addr[7:7] ;
assign n27928 =  ( n27927 ) == ( bv_1_0_n53 )  ;
assign n27929 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n27930 =  ( n27928 ) & (n27929 )  ;
assign n27931 =  ( n27930 ) & (wr )  ;
assign n27932 =  ( n27931 ) ? ( n4782 ) : ( iram_240 ) ;
assign n27933 = wr_addr[7:7] ;
assign n27934 =  ( n27933 ) == ( bv_1_0_n53 )  ;
assign n27935 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n27936 =  ( n27934 ) & (n27935 )  ;
assign n27937 =  ( n27936 ) & (wr )  ;
assign n27938 =  ( n27937 ) ? ( n4841 ) : ( iram_240 ) ;
assign n27939 = wr_addr[7:7] ;
assign n27940 =  ( n27939 ) == ( bv_1_0_n53 )  ;
assign n27941 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n27942 =  ( n27940 ) & (n27941 )  ;
assign n27943 =  ( n27942 ) & (wr )  ;
assign n27944 =  ( n27943 ) ? ( n5449 ) : ( iram_240 ) ;
assign n27945 = wr_addr[7:7] ;
assign n27946 =  ( n27945 ) == ( bv_1_0_n53 )  ;
assign n27947 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n27948 =  ( n27946 ) & (n27947 )  ;
assign n27949 =  ( n27948 ) & (wr )  ;
assign n27950 =  ( n27949 ) ? ( n4906 ) : ( iram_240 ) ;
assign n27951 = wr_addr[7:7] ;
assign n27952 =  ( n27951 ) == ( bv_1_0_n53 )  ;
assign n27953 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n27954 =  ( n27952 ) & (n27953 )  ;
assign n27955 =  ( n27954 ) & (wr )  ;
assign n27956 =  ( n27955 ) ? ( n5485 ) : ( iram_240 ) ;
assign n27957 = wr_addr[7:7] ;
assign n27958 =  ( n27957 ) == ( bv_1_0_n53 )  ;
assign n27959 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n27960 =  ( n27958 ) & (n27959 )  ;
assign n27961 =  ( n27960 ) & (wr )  ;
assign n27962 =  ( n27961 ) ? ( n5512 ) : ( iram_240 ) ;
assign n27963 = wr_addr[7:7] ;
assign n27964 =  ( n27963 ) == ( bv_1_0_n53 )  ;
assign n27965 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n27966 =  ( n27964 ) & (n27965 )  ;
assign n27967 =  ( n27966 ) & (wr )  ;
assign n27968 =  ( n27967 ) ? ( bv_8_0_n69 ) : ( iram_240 ) ;
assign n27969 = wr_addr[7:7] ;
assign n27970 =  ( n27969 ) == ( bv_1_0_n53 )  ;
assign n27971 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n27972 =  ( n27970 ) & (n27971 )  ;
assign n27973 =  ( n27972 ) & (wr )  ;
assign n27974 =  ( n27973 ) ? ( n5071 ) : ( iram_240 ) ;
assign n27975 = wr_addr[7:7] ;
assign n27976 =  ( n27975 ) == ( bv_1_0_n53 )  ;
assign n27977 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n27978 =  ( n27976 ) & (n27977 )  ;
assign n27979 =  ( n27978 ) & (wr )  ;
assign n27980 =  ( n27979 ) ? ( n5096 ) : ( iram_240 ) ;
assign n27981 = wr_addr[7:7] ;
assign n27982 =  ( n27981 ) == ( bv_1_0_n53 )  ;
assign n27983 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n27984 =  ( n27982 ) & (n27983 )  ;
assign n27985 =  ( n27984 ) & (wr )  ;
assign n27986 =  ( n27985 ) ? ( n5123 ) : ( iram_240 ) ;
assign n27987 = wr_addr[7:7] ;
assign n27988 =  ( n27987 ) == ( bv_1_0_n53 )  ;
assign n27989 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n27990 =  ( n27988 ) & (n27989 )  ;
assign n27991 =  ( n27990 ) & (wr )  ;
assign n27992 =  ( n27991 ) ? ( n5165 ) : ( iram_240 ) ;
assign n27993 = wr_addr[7:7] ;
assign n27994 =  ( n27993 ) == ( bv_1_0_n53 )  ;
assign n27995 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n27996 =  ( n27994 ) & (n27995 )  ;
assign n27997 =  ( n27996 ) & (wr )  ;
assign n27998 =  ( n27997 ) ? ( n5204 ) : ( iram_240 ) ;
assign n27999 = wr_addr[7:7] ;
assign n28000 =  ( n27999 ) == ( bv_1_0_n53 )  ;
assign n28001 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n28002 =  ( n28000 ) & (n28001 )  ;
assign n28003 =  ( n28002 ) & (wr )  ;
assign n28004 =  ( n28003 ) ? ( n5262 ) : ( iram_240 ) ;
assign n28005 = wr_addr[7:7] ;
assign n28006 =  ( n28005 ) == ( bv_1_0_n53 )  ;
assign n28007 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n28008 =  ( n28006 ) & (n28007 )  ;
assign n28009 =  ( n28008 ) & (wr )  ;
assign n28010 =  ( n28009 ) ? ( n5298 ) : ( iram_240 ) ;
assign n28011 = wr_addr[7:7] ;
assign n28012 =  ( n28011 ) == ( bv_1_0_n53 )  ;
assign n28013 =  ( wr_addr ) == ( bv_8_240_n549 )  ;
assign n28014 =  ( n28012 ) & (n28013 )  ;
assign n28015 =  ( n28014 ) & (wr )  ;
assign n28016 =  ( n28015 ) ? ( n5325 ) : ( iram_240 ) ;
assign n28017 = wr_addr[7:7] ;
assign n28018 =  ( n28017 ) == ( bv_1_0_n53 )  ;
assign n28019 =  ( wr_addr ) == ( bv_8_241_n551 )  ;
assign n28020 =  ( n28018 ) & (n28019 )  ;
assign n28021 =  ( n28020 ) & (wr )  ;
assign n28022 =  ( n28021 ) ? ( n4782 ) : ( iram_241 ) ;
assign n28023 = wr_addr[7:7] ;
assign n28024 =  ( n28023 ) == ( bv_1_0_n53 )  ;
assign n28025 =  ( wr_addr ) == ( bv_8_241_n551 )  ;
assign n28026 =  ( n28024 ) & (n28025 )  ;
assign n28027 =  ( n28026 ) & (wr )  ;
assign n28028 =  ( n28027 ) ? ( n4841 ) : ( iram_241 ) ;
assign n28029 = wr_addr[7:7] ;
assign n28030 =  ( n28029 ) == ( bv_1_0_n53 )  ;
assign n28031 =  ( wr_addr ) == ( bv_8_241_n551 )  ;
assign n28032 =  ( n28030 ) & (n28031 )  ;
assign n28033 =  ( n28032 ) & (wr )  ;
assign n28034 =  ( n28033 ) ? ( n5449 ) : ( iram_241 ) ;
assign n28035 = wr_addr[7:7] ;
assign n28036 =  ( n28035 ) == ( bv_1_0_n53 )  ;
assign n28037 =  ( wr_addr ) == ( bv_8_241_n551 )  ;
assign n28038 =  ( n28036 ) & (n28037 )  ;
assign n28039 =  ( n28038 ) & (wr )  ;
assign n28040 =  ( n28039 ) ? ( n4906 ) : ( iram_241 ) ;
assign n28041 = wr_addr[7:7] ;
assign n28042 =  ( n28041 ) == ( bv_1_0_n53 )  ;
assign n28043 =  ( wr_addr ) == ( bv_8_241_n551 )  ;
assign n28044 =  ( n28042 ) & (n28043 )  ;
assign n28045 =  ( n28044 ) & (wr )  ;
assign n28046 =  ( n28045 ) ? ( n5485 ) : ( iram_241 ) ;
assign n28047 = wr_addr[7:7] ;
assign n28048 =  ( n28047 ) == ( bv_1_0_n53 )  ;
assign n28049 =  ( wr_addr ) == ( bv_8_241_n551 )  ;
assign n28050 =  ( n28048 ) & (n28049 )  ;
assign n28051 =  ( n28050 ) & (wr )  ;
assign n28052 =  ( n28051 ) ? ( n5512 ) : ( iram_241 ) ;
assign n28053 = wr_addr[7:7] ;
assign n28054 =  ( n28053 ) == ( bv_1_0_n53 )  ;
assign n28055 =  ( wr_addr ) == ( bv_8_241_n551 )  ;
assign n28056 =  ( n28054 ) & (n28055 )  ;
assign n28057 =  ( n28056 ) & (wr )  ;
assign n28058 =  ( n28057 ) ? ( bv_8_0_n69 ) : ( iram_241 ) ;
assign n28059 = wr_addr[7:7] ;
assign n28060 =  ( n28059 ) == ( bv_1_0_n53 )  ;
assign n28061 =  ( wr_addr ) == ( bv_8_241_n551 )  ;
assign n28062 =  ( n28060 ) & (n28061 )  ;
assign n28063 =  ( n28062 ) & (wr )  ;
assign n28064 =  ( n28063 ) ? ( n5071 ) : ( iram_241 ) ;
assign n28065 = wr_addr[7:7] ;
assign n28066 =  ( n28065 ) == ( bv_1_0_n53 )  ;
assign n28067 =  ( wr_addr ) == ( bv_8_241_n551 )  ;
assign n28068 =  ( n28066 ) & (n28067 )  ;
assign n28069 =  ( n28068 ) & (wr )  ;
assign n28070 =  ( n28069 ) ? ( n5096 ) : ( iram_241 ) ;
assign n28071 = wr_addr[7:7] ;
assign n28072 =  ( n28071 ) == ( bv_1_0_n53 )  ;
assign n28073 =  ( wr_addr ) == ( bv_8_241_n551 )  ;
assign n28074 =  ( n28072 ) & (n28073 )  ;
assign n28075 =  ( n28074 ) & (wr )  ;
assign n28076 =  ( n28075 ) ? ( n5123 ) : ( iram_241 ) ;
assign n28077 = wr_addr[7:7] ;
assign n28078 =  ( n28077 ) == ( bv_1_0_n53 )  ;
assign n28079 =  ( wr_addr ) == ( bv_8_241_n551 )  ;
assign n28080 =  ( n28078 ) & (n28079 )  ;
assign n28081 =  ( n28080 ) & (wr )  ;
assign n28082 =  ( n28081 ) ? ( n5165 ) : ( iram_241 ) ;
assign n28083 = wr_addr[7:7] ;
assign n28084 =  ( n28083 ) == ( bv_1_0_n53 )  ;
assign n28085 =  ( wr_addr ) == ( bv_8_241_n551 )  ;
assign n28086 =  ( n28084 ) & (n28085 )  ;
assign n28087 =  ( n28086 ) & (wr )  ;
assign n28088 =  ( n28087 ) ? ( n5204 ) : ( iram_241 ) ;
assign n28089 = wr_addr[7:7] ;
assign n28090 =  ( n28089 ) == ( bv_1_0_n53 )  ;
assign n28091 =  ( wr_addr ) == ( bv_8_241_n551 )  ;
assign n28092 =  ( n28090 ) & (n28091 )  ;
assign n28093 =  ( n28092 ) & (wr )  ;
assign n28094 =  ( n28093 ) ? ( n5262 ) : ( iram_241 ) ;
assign n28095 = wr_addr[7:7] ;
assign n28096 =  ( n28095 ) == ( bv_1_0_n53 )  ;
assign n28097 =  ( wr_addr ) == ( bv_8_241_n551 )  ;
assign n28098 =  ( n28096 ) & (n28097 )  ;
assign n28099 =  ( n28098 ) & (wr )  ;
assign n28100 =  ( n28099 ) ? ( n5298 ) : ( iram_241 ) ;
assign n28101 = wr_addr[7:7] ;
assign n28102 =  ( n28101 ) == ( bv_1_0_n53 )  ;
assign n28103 =  ( wr_addr ) == ( bv_8_241_n551 )  ;
assign n28104 =  ( n28102 ) & (n28103 )  ;
assign n28105 =  ( n28104 ) & (wr )  ;
assign n28106 =  ( n28105 ) ? ( n5325 ) : ( iram_241 ) ;
assign n28107 = wr_addr[7:7] ;
assign n28108 =  ( n28107 ) == ( bv_1_0_n53 )  ;
assign n28109 =  ( wr_addr ) == ( bv_8_242_n553 )  ;
assign n28110 =  ( n28108 ) & (n28109 )  ;
assign n28111 =  ( n28110 ) & (wr )  ;
assign n28112 =  ( n28111 ) ? ( n4782 ) : ( iram_242 ) ;
assign n28113 = wr_addr[7:7] ;
assign n28114 =  ( n28113 ) == ( bv_1_0_n53 )  ;
assign n28115 =  ( wr_addr ) == ( bv_8_242_n553 )  ;
assign n28116 =  ( n28114 ) & (n28115 )  ;
assign n28117 =  ( n28116 ) & (wr )  ;
assign n28118 =  ( n28117 ) ? ( n4841 ) : ( iram_242 ) ;
assign n28119 = wr_addr[7:7] ;
assign n28120 =  ( n28119 ) == ( bv_1_0_n53 )  ;
assign n28121 =  ( wr_addr ) == ( bv_8_242_n553 )  ;
assign n28122 =  ( n28120 ) & (n28121 )  ;
assign n28123 =  ( n28122 ) & (wr )  ;
assign n28124 =  ( n28123 ) ? ( n5449 ) : ( iram_242 ) ;
assign n28125 = wr_addr[7:7] ;
assign n28126 =  ( n28125 ) == ( bv_1_0_n53 )  ;
assign n28127 =  ( wr_addr ) == ( bv_8_242_n553 )  ;
assign n28128 =  ( n28126 ) & (n28127 )  ;
assign n28129 =  ( n28128 ) & (wr )  ;
assign n28130 =  ( n28129 ) ? ( n4906 ) : ( iram_242 ) ;
assign n28131 = wr_addr[7:7] ;
assign n28132 =  ( n28131 ) == ( bv_1_0_n53 )  ;
assign n28133 =  ( wr_addr ) == ( bv_8_242_n553 )  ;
assign n28134 =  ( n28132 ) & (n28133 )  ;
assign n28135 =  ( n28134 ) & (wr )  ;
assign n28136 =  ( n28135 ) ? ( n5485 ) : ( iram_242 ) ;
assign n28137 = wr_addr[7:7] ;
assign n28138 =  ( n28137 ) == ( bv_1_0_n53 )  ;
assign n28139 =  ( wr_addr ) == ( bv_8_242_n553 )  ;
assign n28140 =  ( n28138 ) & (n28139 )  ;
assign n28141 =  ( n28140 ) & (wr )  ;
assign n28142 =  ( n28141 ) ? ( n5512 ) : ( iram_242 ) ;
assign n28143 = wr_addr[7:7] ;
assign n28144 =  ( n28143 ) == ( bv_1_0_n53 )  ;
assign n28145 =  ( wr_addr ) == ( bv_8_242_n553 )  ;
assign n28146 =  ( n28144 ) & (n28145 )  ;
assign n28147 =  ( n28146 ) & (wr )  ;
assign n28148 =  ( n28147 ) ? ( bv_8_0_n69 ) : ( iram_242 ) ;
assign n28149 = wr_addr[7:7] ;
assign n28150 =  ( n28149 ) == ( bv_1_0_n53 )  ;
assign n28151 =  ( wr_addr ) == ( bv_8_242_n553 )  ;
assign n28152 =  ( n28150 ) & (n28151 )  ;
assign n28153 =  ( n28152 ) & (wr )  ;
assign n28154 =  ( n28153 ) ? ( n5071 ) : ( iram_242 ) ;
assign n28155 = wr_addr[7:7] ;
assign n28156 =  ( n28155 ) == ( bv_1_0_n53 )  ;
assign n28157 =  ( wr_addr ) == ( bv_8_242_n553 )  ;
assign n28158 =  ( n28156 ) & (n28157 )  ;
assign n28159 =  ( n28158 ) & (wr )  ;
assign n28160 =  ( n28159 ) ? ( n5096 ) : ( iram_242 ) ;
assign n28161 = wr_addr[7:7] ;
assign n28162 =  ( n28161 ) == ( bv_1_0_n53 )  ;
assign n28163 =  ( wr_addr ) == ( bv_8_242_n553 )  ;
assign n28164 =  ( n28162 ) & (n28163 )  ;
assign n28165 =  ( n28164 ) & (wr )  ;
assign n28166 =  ( n28165 ) ? ( n5123 ) : ( iram_242 ) ;
assign n28167 = wr_addr[7:7] ;
assign n28168 =  ( n28167 ) == ( bv_1_0_n53 )  ;
assign n28169 =  ( wr_addr ) == ( bv_8_242_n553 )  ;
assign n28170 =  ( n28168 ) & (n28169 )  ;
assign n28171 =  ( n28170 ) & (wr )  ;
assign n28172 =  ( n28171 ) ? ( n5165 ) : ( iram_242 ) ;
assign n28173 = wr_addr[7:7] ;
assign n28174 =  ( n28173 ) == ( bv_1_0_n53 )  ;
assign n28175 =  ( wr_addr ) == ( bv_8_242_n553 )  ;
assign n28176 =  ( n28174 ) & (n28175 )  ;
assign n28177 =  ( n28176 ) & (wr )  ;
assign n28178 =  ( n28177 ) ? ( n5204 ) : ( iram_242 ) ;
assign n28179 = wr_addr[7:7] ;
assign n28180 =  ( n28179 ) == ( bv_1_0_n53 )  ;
assign n28181 =  ( wr_addr ) == ( bv_8_242_n553 )  ;
assign n28182 =  ( n28180 ) & (n28181 )  ;
assign n28183 =  ( n28182 ) & (wr )  ;
assign n28184 =  ( n28183 ) ? ( n5262 ) : ( iram_242 ) ;
assign n28185 = wr_addr[7:7] ;
assign n28186 =  ( n28185 ) == ( bv_1_0_n53 )  ;
assign n28187 =  ( wr_addr ) == ( bv_8_242_n553 )  ;
assign n28188 =  ( n28186 ) & (n28187 )  ;
assign n28189 =  ( n28188 ) & (wr )  ;
assign n28190 =  ( n28189 ) ? ( n5298 ) : ( iram_242 ) ;
assign n28191 = wr_addr[7:7] ;
assign n28192 =  ( n28191 ) == ( bv_1_0_n53 )  ;
assign n28193 =  ( wr_addr ) == ( bv_8_242_n553 )  ;
assign n28194 =  ( n28192 ) & (n28193 )  ;
assign n28195 =  ( n28194 ) & (wr )  ;
assign n28196 =  ( n28195 ) ? ( n5325 ) : ( iram_242 ) ;
assign n28197 = wr_addr[7:7] ;
assign n28198 =  ( n28197 ) == ( bv_1_0_n53 )  ;
assign n28199 =  ( wr_addr ) == ( bv_8_243_n555 )  ;
assign n28200 =  ( n28198 ) & (n28199 )  ;
assign n28201 =  ( n28200 ) & (wr )  ;
assign n28202 =  ( n28201 ) ? ( n4782 ) : ( iram_243 ) ;
assign n28203 = wr_addr[7:7] ;
assign n28204 =  ( n28203 ) == ( bv_1_0_n53 )  ;
assign n28205 =  ( wr_addr ) == ( bv_8_243_n555 )  ;
assign n28206 =  ( n28204 ) & (n28205 )  ;
assign n28207 =  ( n28206 ) & (wr )  ;
assign n28208 =  ( n28207 ) ? ( n4841 ) : ( iram_243 ) ;
assign n28209 = wr_addr[7:7] ;
assign n28210 =  ( n28209 ) == ( bv_1_0_n53 )  ;
assign n28211 =  ( wr_addr ) == ( bv_8_243_n555 )  ;
assign n28212 =  ( n28210 ) & (n28211 )  ;
assign n28213 =  ( n28212 ) & (wr )  ;
assign n28214 =  ( n28213 ) ? ( n5449 ) : ( iram_243 ) ;
assign n28215 = wr_addr[7:7] ;
assign n28216 =  ( n28215 ) == ( bv_1_0_n53 )  ;
assign n28217 =  ( wr_addr ) == ( bv_8_243_n555 )  ;
assign n28218 =  ( n28216 ) & (n28217 )  ;
assign n28219 =  ( n28218 ) & (wr )  ;
assign n28220 =  ( n28219 ) ? ( n4906 ) : ( iram_243 ) ;
assign n28221 = wr_addr[7:7] ;
assign n28222 =  ( n28221 ) == ( bv_1_0_n53 )  ;
assign n28223 =  ( wr_addr ) == ( bv_8_243_n555 )  ;
assign n28224 =  ( n28222 ) & (n28223 )  ;
assign n28225 =  ( n28224 ) & (wr )  ;
assign n28226 =  ( n28225 ) ? ( n5485 ) : ( iram_243 ) ;
assign n28227 = wr_addr[7:7] ;
assign n28228 =  ( n28227 ) == ( bv_1_0_n53 )  ;
assign n28229 =  ( wr_addr ) == ( bv_8_243_n555 )  ;
assign n28230 =  ( n28228 ) & (n28229 )  ;
assign n28231 =  ( n28230 ) & (wr )  ;
assign n28232 =  ( n28231 ) ? ( n5512 ) : ( iram_243 ) ;
assign n28233 = wr_addr[7:7] ;
assign n28234 =  ( n28233 ) == ( bv_1_0_n53 )  ;
assign n28235 =  ( wr_addr ) == ( bv_8_243_n555 )  ;
assign n28236 =  ( n28234 ) & (n28235 )  ;
assign n28237 =  ( n28236 ) & (wr )  ;
assign n28238 =  ( n28237 ) ? ( bv_8_0_n69 ) : ( iram_243 ) ;
assign n28239 = wr_addr[7:7] ;
assign n28240 =  ( n28239 ) == ( bv_1_0_n53 )  ;
assign n28241 =  ( wr_addr ) == ( bv_8_243_n555 )  ;
assign n28242 =  ( n28240 ) & (n28241 )  ;
assign n28243 =  ( n28242 ) & (wr )  ;
assign n28244 =  ( n28243 ) ? ( n5071 ) : ( iram_243 ) ;
assign n28245 = wr_addr[7:7] ;
assign n28246 =  ( n28245 ) == ( bv_1_0_n53 )  ;
assign n28247 =  ( wr_addr ) == ( bv_8_243_n555 )  ;
assign n28248 =  ( n28246 ) & (n28247 )  ;
assign n28249 =  ( n28248 ) & (wr )  ;
assign n28250 =  ( n28249 ) ? ( n5096 ) : ( iram_243 ) ;
assign n28251 = wr_addr[7:7] ;
assign n28252 =  ( n28251 ) == ( bv_1_0_n53 )  ;
assign n28253 =  ( wr_addr ) == ( bv_8_243_n555 )  ;
assign n28254 =  ( n28252 ) & (n28253 )  ;
assign n28255 =  ( n28254 ) & (wr )  ;
assign n28256 =  ( n28255 ) ? ( n5123 ) : ( iram_243 ) ;
assign n28257 = wr_addr[7:7] ;
assign n28258 =  ( n28257 ) == ( bv_1_0_n53 )  ;
assign n28259 =  ( wr_addr ) == ( bv_8_243_n555 )  ;
assign n28260 =  ( n28258 ) & (n28259 )  ;
assign n28261 =  ( n28260 ) & (wr )  ;
assign n28262 =  ( n28261 ) ? ( n5165 ) : ( iram_243 ) ;
assign n28263 = wr_addr[7:7] ;
assign n28264 =  ( n28263 ) == ( bv_1_0_n53 )  ;
assign n28265 =  ( wr_addr ) == ( bv_8_243_n555 )  ;
assign n28266 =  ( n28264 ) & (n28265 )  ;
assign n28267 =  ( n28266 ) & (wr )  ;
assign n28268 =  ( n28267 ) ? ( n5204 ) : ( iram_243 ) ;
assign n28269 = wr_addr[7:7] ;
assign n28270 =  ( n28269 ) == ( bv_1_0_n53 )  ;
assign n28271 =  ( wr_addr ) == ( bv_8_243_n555 )  ;
assign n28272 =  ( n28270 ) & (n28271 )  ;
assign n28273 =  ( n28272 ) & (wr )  ;
assign n28274 =  ( n28273 ) ? ( n5262 ) : ( iram_243 ) ;
assign n28275 = wr_addr[7:7] ;
assign n28276 =  ( n28275 ) == ( bv_1_0_n53 )  ;
assign n28277 =  ( wr_addr ) == ( bv_8_243_n555 )  ;
assign n28278 =  ( n28276 ) & (n28277 )  ;
assign n28279 =  ( n28278 ) & (wr )  ;
assign n28280 =  ( n28279 ) ? ( n5298 ) : ( iram_243 ) ;
assign n28281 = wr_addr[7:7] ;
assign n28282 =  ( n28281 ) == ( bv_1_0_n53 )  ;
assign n28283 =  ( wr_addr ) == ( bv_8_243_n555 )  ;
assign n28284 =  ( n28282 ) & (n28283 )  ;
assign n28285 =  ( n28284 ) & (wr )  ;
assign n28286 =  ( n28285 ) ? ( n5325 ) : ( iram_243 ) ;
assign n28287 = wr_addr[7:7] ;
assign n28288 =  ( n28287 ) == ( bv_1_0_n53 )  ;
assign n28289 =  ( wr_addr ) == ( bv_8_244_n557 )  ;
assign n28290 =  ( n28288 ) & (n28289 )  ;
assign n28291 =  ( n28290 ) & (wr )  ;
assign n28292 =  ( n28291 ) ? ( n4782 ) : ( iram_244 ) ;
assign n28293 = wr_addr[7:7] ;
assign n28294 =  ( n28293 ) == ( bv_1_0_n53 )  ;
assign n28295 =  ( wr_addr ) == ( bv_8_244_n557 )  ;
assign n28296 =  ( n28294 ) & (n28295 )  ;
assign n28297 =  ( n28296 ) & (wr )  ;
assign n28298 =  ( n28297 ) ? ( n4841 ) : ( iram_244 ) ;
assign n28299 = wr_addr[7:7] ;
assign n28300 =  ( n28299 ) == ( bv_1_0_n53 )  ;
assign n28301 =  ( wr_addr ) == ( bv_8_244_n557 )  ;
assign n28302 =  ( n28300 ) & (n28301 )  ;
assign n28303 =  ( n28302 ) & (wr )  ;
assign n28304 =  ( n28303 ) ? ( n5449 ) : ( iram_244 ) ;
assign n28305 = wr_addr[7:7] ;
assign n28306 =  ( n28305 ) == ( bv_1_0_n53 )  ;
assign n28307 =  ( wr_addr ) == ( bv_8_244_n557 )  ;
assign n28308 =  ( n28306 ) & (n28307 )  ;
assign n28309 =  ( n28308 ) & (wr )  ;
assign n28310 =  ( n28309 ) ? ( n4906 ) : ( iram_244 ) ;
assign n28311 = wr_addr[7:7] ;
assign n28312 =  ( n28311 ) == ( bv_1_0_n53 )  ;
assign n28313 =  ( wr_addr ) == ( bv_8_244_n557 )  ;
assign n28314 =  ( n28312 ) & (n28313 )  ;
assign n28315 =  ( n28314 ) & (wr )  ;
assign n28316 =  ( n28315 ) ? ( n5485 ) : ( iram_244 ) ;
assign n28317 = wr_addr[7:7] ;
assign n28318 =  ( n28317 ) == ( bv_1_0_n53 )  ;
assign n28319 =  ( wr_addr ) == ( bv_8_244_n557 )  ;
assign n28320 =  ( n28318 ) & (n28319 )  ;
assign n28321 =  ( n28320 ) & (wr )  ;
assign n28322 =  ( n28321 ) ? ( n5512 ) : ( iram_244 ) ;
assign n28323 = wr_addr[7:7] ;
assign n28324 =  ( n28323 ) == ( bv_1_0_n53 )  ;
assign n28325 =  ( wr_addr ) == ( bv_8_244_n557 )  ;
assign n28326 =  ( n28324 ) & (n28325 )  ;
assign n28327 =  ( n28326 ) & (wr )  ;
assign n28328 =  ( n28327 ) ? ( bv_8_0_n69 ) : ( iram_244 ) ;
assign n28329 = wr_addr[7:7] ;
assign n28330 =  ( n28329 ) == ( bv_1_0_n53 )  ;
assign n28331 =  ( wr_addr ) == ( bv_8_244_n557 )  ;
assign n28332 =  ( n28330 ) & (n28331 )  ;
assign n28333 =  ( n28332 ) & (wr )  ;
assign n28334 =  ( n28333 ) ? ( n5071 ) : ( iram_244 ) ;
assign n28335 = wr_addr[7:7] ;
assign n28336 =  ( n28335 ) == ( bv_1_0_n53 )  ;
assign n28337 =  ( wr_addr ) == ( bv_8_244_n557 )  ;
assign n28338 =  ( n28336 ) & (n28337 )  ;
assign n28339 =  ( n28338 ) & (wr )  ;
assign n28340 =  ( n28339 ) ? ( n5096 ) : ( iram_244 ) ;
assign n28341 = wr_addr[7:7] ;
assign n28342 =  ( n28341 ) == ( bv_1_0_n53 )  ;
assign n28343 =  ( wr_addr ) == ( bv_8_244_n557 )  ;
assign n28344 =  ( n28342 ) & (n28343 )  ;
assign n28345 =  ( n28344 ) & (wr )  ;
assign n28346 =  ( n28345 ) ? ( n5123 ) : ( iram_244 ) ;
assign n28347 = wr_addr[7:7] ;
assign n28348 =  ( n28347 ) == ( bv_1_0_n53 )  ;
assign n28349 =  ( wr_addr ) == ( bv_8_244_n557 )  ;
assign n28350 =  ( n28348 ) & (n28349 )  ;
assign n28351 =  ( n28350 ) & (wr )  ;
assign n28352 =  ( n28351 ) ? ( n5165 ) : ( iram_244 ) ;
assign n28353 = wr_addr[7:7] ;
assign n28354 =  ( n28353 ) == ( bv_1_0_n53 )  ;
assign n28355 =  ( wr_addr ) == ( bv_8_244_n557 )  ;
assign n28356 =  ( n28354 ) & (n28355 )  ;
assign n28357 =  ( n28356 ) & (wr )  ;
assign n28358 =  ( n28357 ) ? ( n5204 ) : ( iram_244 ) ;
assign n28359 = wr_addr[7:7] ;
assign n28360 =  ( n28359 ) == ( bv_1_0_n53 )  ;
assign n28361 =  ( wr_addr ) == ( bv_8_244_n557 )  ;
assign n28362 =  ( n28360 ) & (n28361 )  ;
assign n28363 =  ( n28362 ) & (wr )  ;
assign n28364 =  ( n28363 ) ? ( n5262 ) : ( iram_244 ) ;
assign n28365 = wr_addr[7:7] ;
assign n28366 =  ( n28365 ) == ( bv_1_0_n53 )  ;
assign n28367 =  ( wr_addr ) == ( bv_8_244_n557 )  ;
assign n28368 =  ( n28366 ) & (n28367 )  ;
assign n28369 =  ( n28368 ) & (wr )  ;
assign n28370 =  ( n28369 ) ? ( n5298 ) : ( iram_244 ) ;
assign n28371 = wr_addr[7:7] ;
assign n28372 =  ( n28371 ) == ( bv_1_0_n53 )  ;
assign n28373 =  ( wr_addr ) == ( bv_8_244_n557 )  ;
assign n28374 =  ( n28372 ) & (n28373 )  ;
assign n28375 =  ( n28374 ) & (wr )  ;
assign n28376 =  ( n28375 ) ? ( n5325 ) : ( iram_244 ) ;
assign n28377 = wr_addr[7:7] ;
assign n28378 =  ( n28377 ) == ( bv_1_0_n53 )  ;
assign n28379 =  ( wr_addr ) == ( bv_8_245_n559 )  ;
assign n28380 =  ( n28378 ) & (n28379 )  ;
assign n28381 =  ( n28380 ) & (wr )  ;
assign n28382 =  ( n28381 ) ? ( n4782 ) : ( iram_245 ) ;
assign n28383 = wr_addr[7:7] ;
assign n28384 =  ( n28383 ) == ( bv_1_0_n53 )  ;
assign n28385 =  ( wr_addr ) == ( bv_8_245_n559 )  ;
assign n28386 =  ( n28384 ) & (n28385 )  ;
assign n28387 =  ( n28386 ) & (wr )  ;
assign n28388 =  ( n28387 ) ? ( n4841 ) : ( iram_245 ) ;
assign n28389 = wr_addr[7:7] ;
assign n28390 =  ( n28389 ) == ( bv_1_0_n53 )  ;
assign n28391 =  ( wr_addr ) == ( bv_8_245_n559 )  ;
assign n28392 =  ( n28390 ) & (n28391 )  ;
assign n28393 =  ( n28392 ) & (wr )  ;
assign n28394 =  ( n28393 ) ? ( n5449 ) : ( iram_245 ) ;
assign n28395 = wr_addr[7:7] ;
assign n28396 =  ( n28395 ) == ( bv_1_0_n53 )  ;
assign n28397 =  ( wr_addr ) == ( bv_8_245_n559 )  ;
assign n28398 =  ( n28396 ) & (n28397 )  ;
assign n28399 =  ( n28398 ) & (wr )  ;
assign n28400 =  ( n28399 ) ? ( n4906 ) : ( iram_245 ) ;
assign n28401 = wr_addr[7:7] ;
assign n28402 =  ( n28401 ) == ( bv_1_0_n53 )  ;
assign n28403 =  ( wr_addr ) == ( bv_8_245_n559 )  ;
assign n28404 =  ( n28402 ) & (n28403 )  ;
assign n28405 =  ( n28404 ) & (wr )  ;
assign n28406 =  ( n28405 ) ? ( n5485 ) : ( iram_245 ) ;
assign n28407 = wr_addr[7:7] ;
assign n28408 =  ( n28407 ) == ( bv_1_0_n53 )  ;
assign n28409 =  ( wr_addr ) == ( bv_8_245_n559 )  ;
assign n28410 =  ( n28408 ) & (n28409 )  ;
assign n28411 =  ( n28410 ) & (wr )  ;
assign n28412 =  ( n28411 ) ? ( n5512 ) : ( iram_245 ) ;
assign n28413 = wr_addr[7:7] ;
assign n28414 =  ( n28413 ) == ( bv_1_0_n53 )  ;
assign n28415 =  ( wr_addr ) == ( bv_8_245_n559 )  ;
assign n28416 =  ( n28414 ) & (n28415 )  ;
assign n28417 =  ( n28416 ) & (wr )  ;
assign n28418 =  ( n28417 ) ? ( bv_8_0_n69 ) : ( iram_245 ) ;
assign n28419 = wr_addr[7:7] ;
assign n28420 =  ( n28419 ) == ( bv_1_0_n53 )  ;
assign n28421 =  ( wr_addr ) == ( bv_8_245_n559 )  ;
assign n28422 =  ( n28420 ) & (n28421 )  ;
assign n28423 =  ( n28422 ) & (wr )  ;
assign n28424 =  ( n28423 ) ? ( n5071 ) : ( iram_245 ) ;
assign n28425 = wr_addr[7:7] ;
assign n28426 =  ( n28425 ) == ( bv_1_0_n53 )  ;
assign n28427 =  ( wr_addr ) == ( bv_8_245_n559 )  ;
assign n28428 =  ( n28426 ) & (n28427 )  ;
assign n28429 =  ( n28428 ) & (wr )  ;
assign n28430 =  ( n28429 ) ? ( n5096 ) : ( iram_245 ) ;
assign n28431 = wr_addr[7:7] ;
assign n28432 =  ( n28431 ) == ( bv_1_0_n53 )  ;
assign n28433 =  ( wr_addr ) == ( bv_8_245_n559 )  ;
assign n28434 =  ( n28432 ) & (n28433 )  ;
assign n28435 =  ( n28434 ) & (wr )  ;
assign n28436 =  ( n28435 ) ? ( n5123 ) : ( iram_245 ) ;
assign n28437 = wr_addr[7:7] ;
assign n28438 =  ( n28437 ) == ( bv_1_0_n53 )  ;
assign n28439 =  ( wr_addr ) == ( bv_8_245_n559 )  ;
assign n28440 =  ( n28438 ) & (n28439 )  ;
assign n28441 =  ( n28440 ) & (wr )  ;
assign n28442 =  ( n28441 ) ? ( n5165 ) : ( iram_245 ) ;
assign n28443 = wr_addr[7:7] ;
assign n28444 =  ( n28443 ) == ( bv_1_0_n53 )  ;
assign n28445 =  ( wr_addr ) == ( bv_8_245_n559 )  ;
assign n28446 =  ( n28444 ) & (n28445 )  ;
assign n28447 =  ( n28446 ) & (wr )  ;
assign n28448 =  ( n28447 ) ? ( n5204 ) : ( iram_245 ) ;
assign n28449 = wr_addr[7:7] ;
assign n28450 =  ( n28449 ) == ( bv_1_0_n53 )  ;
assign n28451 =  ( wr_addr ) == ( bv_8_245_n559 )  ;
assign n28452 =  ( n28450 ) & (n28451 )  ;
assign n28453 =  ( n28452 ) & (wr )  ;
assign n28454 =  ( n28453 ) ? ( n5262 ) : ( iram_245 ) ;
assign n28455 = wr_addr[7:7] ;
assign n28456 =  ( n28455 ) == ( bv_1_0_n53 )  ;
assign n28457 =  ( wr_addr ) == ( bv_8_245_n559 )  ;
assign n28458 =  ( n28456 ) & (n28457 )  ;
assign n28459 =  ( n28458 ) & (wr )  ;
assign n28460 =  ( n28459 ) ? ( n5298 ) : ( iram_245 ) ;
assign n28461 = wr_addr[7:7] ;
assign n28462 =  ( n28461 ) == ( bv_1_0_n53 )  ;
assign n28463 =  ( wr_addr ) == ( bv_8_245_n559 )  ;
assign n28464 =  ( n28462 ) & (n28463 )  ;
assign n28465 =  ( n28464 ) & (wr )  ;
assign n28466 =  ( n28465 ) ? ( n5325 ) : ( iram_245 ) ;
assign n28467 = wr_addr[7:7] ;
assign n28468 =  ( n28467 ) == ( bv_1_0_n53 )  ;
assign n28469 =  ( wr_addr ) == ( bv_8_246_n561 )  ;
assign n28470 =  ( n28468 ) & (n28469 )  ;
assign n28471 =  ( n28470 ) & (wr )  ;
assign n28472 =  ( n28471 ) ? ( n4782 ) : ( iram_246 ) ;
assign n28473 = wr_addr[7:7] ;
assign n28474 =  ( n28473 ) == ( bv_1_0_n53 )  ;
assign n28475 =  ( wr_addr ) == ( bv_8_246_n561 )  ;
assign n28476 =  ( n28474 ) & (n28475 )  ;
assign n28477 =  ( n28476 ) & (wr )  ;
assign n28478 =  ( n28477 ) ? ( n4841 ) : ( iram_246 ) ;
assign n28479 = wr_addr[7:7] ;
assign n28480 =  ( n28479 ) == ( bv_1_0_n53 )  ;
assign n28481 =  ( wr_addr ) == ( bv_8_246_n561 )  ;
assign n28482 =  ( n28480 ) & (n28481 )  ;
assign n28483 =  ( n28482 ) & (wr )  ;
assign n28484 =  ( n28483 ) ? ( n5449 ) : ( iram_246 ) ;
assign n28485 = wr_addr[7:7] ;
assign n28486 =  ( n28485 ) == ( bv_1_0_n53 )  ;
assign n28487 =  ( wr_addr ) == ( bv_8_246_n561 )  ;
assign n28488 =  ( n28486 ) & (n28487 )  ;
assign n28489 =  ( n28488 ) & (wr )  ;
assign n28490 =  ( n28489 ) ? ( n4906 ) : ( iram_246 ) ;
assign n28491 = wr_addr[7:7] ;
assign n28492 =  ( n28491 ) == ( bv_1_0_n53 )  ;
assign n28493 =  ( wr_addr ) == ( bv_8_246_n561 )  ;
assign n28494 =  ( n28492 ) & (n28493 )  ;
assign n28495 =  ( n28494 ) & (wr )  ;
assign n28496 =  ( n28495 ) ? ( n5485 ) : ( iram_246 ) ;
assign n28497 = wr_addr[7:7] ;
assign n28498 =  ( n28497 ) == ( bv_1_0_n53 )  ;
assign n28499 =  ( wr_addr ) == ( bv_8_246_n561 )  ;
assign n28500 =  ( n28498 ) & (n28499 )  ;
assign n28501 =  ( n28500 ) & (wr )  ;
assign n28502 =  ( n28501 ) ? ( n5512 ) : ( iram_246 ) ;
assign n28503 = wr_addr[7:7] ;
assign n28504 =  ( n28503 ) == ( bv_1_0_n53 )  ;
assign n28505 =  ( wr_addr ) == ( bv_8_246_n561 )  ;
assign n28506 =  ( n28504 ) & (n28505 )  ;
assign n28507 =  ( n28506 ) & (wr )  ;
assign n28508 =  ( n28507 ) ? ( bv_8_0_n69 ) : ( iram_246 ) ;
assign n28509 = wr_addr[7:7] ;
assign n28510 =  ( n28509 ) == ( bv_1_0_n53 )  ;
assign n28511 =  ( wr_addr ) == ( bv_8_246_n561 )  ;
assign n28512 =  ( n28510 ) & (n28511 )  ;
assign n28513 =  ( n28512 ) & (wr )  ;
assign n28514 =  ( n28513 ) ? ( n5071 ) : ( iram_246 ) ;
assign n28515 = wr_addr[7:7] ;
assign n28516 =  ( n28515 ) == ( bv_1_0_n53 )  ;
assign n28517 =  ( wr_addr ) == ( bv_8_246_n561 )  ;
assign n28518 =  ( n28516 ) & (n28517 )  ;
assign n28519 =  ( n28518 ) & (wr )  ;
assign n28520 =  ( n28519 ) ? ( n5096 ) : ( iram_246 ) ;
assign n28521 = wr_addr[7:7] ;
assign n28522 =  ( n28521 ) == ( bv_1_0_n53 )  ;
assign n28523 =  ( wr_addr ) == ( bv_8_246_n561 )  ;
assign n28524 =  ( n28522 ) & (n28523 )  ;
assign n28525 =  ( n28524 ) & (wr )  ;
assign n28526 =  ( n28525 ) ? ( n5123 ) : ( iram_246 ) ;
assign n28527 = wr_addr[7:7] ;
assign n28528 =  ( n28527 ) == ( bv_1_0_n53 )  ;
assign n28529 =  ( wr_addr ) == ( bv_8_246_n561 )  ;
assign n28530 =  ( n28528 ) & (n28529 )  ;
assign n28531 =  ( n28530 ) & (wr )  ;
assign n28532 =  ( n28531 ) ? ( n5165 ) : ( iram_246 ) ;
assign n28533 = wr_addr[7:7] ;
assign n28534 =  ( n28533 ) == ( bv_1_0_n53 )  ;
assign n28535 =  ( wr_addr ) == ( bv_8_246_n561 )  ;
assign n28536 =  ( n28534 ) & (n28535 )  ;
assign n28537 =  ( n28536 ) & (wr )  ;
assign n28538 =  ( n28537 ) ? ( n5204 ) : ( iram_246 ) ;
assign n28539 = wr_addr[7:7] ;
assign n28540 =  ( n28539 ) == ( bv_1_0_n53 )  ;
assign n28541 =  ( wr_addr ) == ( bv_8_246_n561 )  ;
assign n28542 =  ( n28540 ) & (n28541 )  ;
assign n28543 =  ( n28542 ) & (wr )  ;
assign n28544 =  ( n28543 ) ? ( n5262 ) : ( iram_246 ) ;
assign n28545 = wr_addr[7:7] ;
assign n28546 =  ( n28545 ) == ( bv_1_0_n53 )  ;
assign n28547 =  ( wr_addr ) == ( bv_8_246_n561 )  ;
assign n28548 =  ( n28546 ) & (n28547 )  ;
assign n28549 =  ( n28548 ) & (wr )  ;
assign n28550 =  ( n28549 ) ? ( n5298 ) : ( iram_246 ) ;
assign n28551 = wr_addr[7:7] ;
assign n28552 =  ( n28551 ) == ( bv_1_0_n53 )  ;
assign n28553 =  ( wr_addr ) == ( bv_8_246_n561 )  ;
assign n28554 =  ( n28552 ) & (n28553 )  ;
assign n28555 =  ( n28554 ) & (wr )  ;
assign n28556 =  ( n28555 ) ? ( n5325 ) : ( iram_246 ) ;
assign n28557 = wr_addr[7:7] ;
assign n28558 =  ( n28557 ) == ( bv_1_0_n53 )  ;
assign n28559 =  ( wr_addr ) == ( bv_8_247_n563 )  ;
assign n28560 =  ( n28558 ) & (n28559 )  ;
assign n28561 =  ( n28560 ) & (wr )  ;
assign n28562 =  ( n28561 ) ? ( n4782 ) : ( iram_247 ) ;
assign n28563 = wr_addr[7:7] ;
assign n28564 =  ( n28563 ) == ( bv_1_0_n53 )  ;
assign n28565 =  ( wr_addr ) == ( bv_8_247_n563 )  ;
assign n28566 =  ( n28564 ) & (n28565 )  ;
assign n28567 =  ( n28566 ) & (wr )  ;
assign n28568 =  ( n28567 ) ? ( n4841 ) : ( iram_247 ) ;
assign n28569 = wr_addr[7:7] ;
assign n28570 =  ( n28569 ) == ( bv_1_0_n53 )  ;
assign n28571 =  ( wr_addr ) == ( bv_8_247_n563 )  ;
assign n28572 =  ( n28570 ) & (n28571 )  ;
assign n28573 =  ( n28572 ) & (wr )  ;
assign n28574 =  ( n28573 ) ? ( n5449 ) : ( iram_247 ) ;
assign n28575 = wr_addr[7:7] ;
assign n28576 =  ( n28575 ) == ( bv_1_0_n53 )  ;
assign n28577 =  ( wr_addr ) == ( bv_8_247_n563 )  ;
assign n28578 =  ( n28576 ) & (n28577 )  ;
assign n28579 =  ( n28578 ) & (wr )  ;
assign n28580 =  ( n28579 ) ? ( n4906 ) : ( iram_247 ) ;
assign n28581 = wr_addr[7:7] ;
assign n28582 =  ( n28581 ) == ( bv_1_0_n53 )  ;
assign n28583 =  ( wr_addr ) == ( bv_8_247_n563 )  ;
assign n28584 =  ( n28582 ) & (n28583 )  ;
assign n28585 =  ( n28584 ) & (wr )  ;
assign n28586 =  ( n28585 ) ? ( n5485 ) : ( iram_247 ) ;
assign n28587 = wr_addr[7:7] ;
assign n28588 =  ( n28587 ) == ( bv_1_0_n53 )  ;
assign n28589 =  ( wr_addr ) == ( bv_8_247_n563 )  ;
assign n28590 =  ( n28588 ) & (n28589 )  ;
assign n28591 =  ( n28590 ) & (wr )  ;
assign n28592 =  ( n28591 ) ? ( n5512 ) : ( iram_247 ) ;
assign n28593 = wr_addr[7:7] ;
assign n28594 =  ( n28593 ) == ( bv_1_0_n53 )  ;
assign n28595 =  ( wr_addr ) == ( bv_8_247_n563 )  ;
assign n28596 =  ( n28594 ) & (n28595 )  ;
assign n28597 =  ( n28596 ) & (wr )  ;
assign n28598 =  ( n28597 ) ? ( bv_8_0_n69 ) : ( iram_247 ) ;
assign n28599 = wr_addr[7:7] ;
assign n28600 =  ( n28599 ) == ( bv_1_0_n53 )  ;
assign n28601 =  ( wr_addr ) == ( bv_8_247_n563 )  ;
assign n28602 =  ( n28600 ) & (n28601 )  ;
assign n28603 =  ( n28602 ) & (wr )  ;
assign n28604 =  ( n28603 ) ? ( n5071 ) : ( iram_247 ) ;
assign n28605 = wr_addr[7:7] ;
assign n28606 =  ( n28605 ) == ( bv_1_0_n53 )  ;
assign n28607 =  ( wr_addr ) == ( bv_8_247_n563 )  ;
assign n28608 =  ( n28606 ) & (n28607 )  ;
assign n28609 =  ( n28608 ) & (wr )  ;
assign n28610 =  ( n28609 ) ? ( n5096 ) : ( iram_247 ) ;
assign n28611 = wr_addr[7:7] ;
assign n28612 =  ( n28611 ) == ( bv_1_0_n53 )  ;
assign n28613 =  ( wr_addr ) == ( bv_8_247_n563 )  ;
assign n28614 =  ( n28612 ) & (n28613 )  ;
assign n28615 =  ( n28614 ) & (wr )  ;
assign n28616 =  ( n28615 ) ? ( n5123 ) : ( iram_247 ) ;
assign n28617 = wr_addr[7:7] ;
assign n28618 =  ( n28617 ) == ( bv_1_0_n53 )  ;
assign n28619 =  ( wr_addr ) == ( bv_8_247_n563 )  ;
assign n28620 =  ( n28618 ) & (n28619 )  ;
assign n28621 =  ( n28620 ) & (wr )  ;
assign n28622 =  ( n28621 ) ? ( n5165 ) : ( iram_247 ) ;
assign n28623 = wr_addr[7:7] ;
assign n28624 =  ( n28623 ) == ( bv_1_0_n53 )  ;
assign n28625 =  ( wr_addr ) == ( bv_8_247_n563 )  ;
assign n28626 =  ( n28624 ) & (n28625 )  ;
assign n28627 =  ( n28626 ) & (wr )  ;
assign n28628 =  ( n28627 ) ? ( n5204 ) : ( iram_247 ) ;
assign n28629 = wr_addr[7:7] ;
assign n28630 =  ( n28629 ) == ( bv_1_0_n53 )  ;
assign n28631 =  ( wr_addr ) == ( bv_8_247_n563 )  ;
assign n28632 =  ( n28630 ) & (n28631 )  ;
assign n28633 =  ( n28632 ) & (wr )  ;
assign n28634 =  ( n28633 ) ? ( n5262 ) : ( iram_247 ) ;
assign n28635 = wr_addr[7:7] ;
assign n28636 =  ( n28635 ) == ( bv_1_0_n53 )  ;
assign n28637 =  ( wr_addr ) == ( bv_8_247_n563 )  ;
assign n28638 =  ( n28636 ) & (n28637 )  ;
assign n28639 =  ( n28638 ) & (wr )  ;
assign n28640 =  ( n28639 ) ? ( n5298 ) : ( iram_247 ) ;
assign n28641 = wr_addr[7:7] ;
assign n28642 =  ( n28641 ) == ( bv_1_0_n53 )  ;
assign n28643 =  ( wr_addr ) == ( bv_8_247_n563 )  ;
assign n28644 =  ( n28642 ) & (n28643 )  ;
assign n28645 =  ( n28644 ) & (wr )  ;
assign n28646 =  ( n28645 ) ? ( n5325 ) : ( iram_247 ) ;
assign n28647 = wr_addr[7:7] ;
assign n28648 =  ( n28647 ) == ( bv_1_0_n53 )  ;
assign n28649 =  ( wr_addr ) == ( bv_8_248_n565 )  ;
assign n28650 =  ( n28648 ) & (n28649 )  ;
assign n28651 =  ( n28650 ) & (wr )  ;
assign n28652 =  ( n28651 ) ? ( n4782 ) : ( iram_248 ) ;
assign n28653 = wr_addr[7:7] ;
assign n28654 =  ( n28653 ) == ( bv_1_0_n53 )  ;
assign n28655 =  ( wr_addr ) == ( bv_8_248_n565 )  ;
assign n28656 =  ( n28654 ) & (n28655 )  ;
assign n28657 =  ( n28656 ) & (wr )  ;
assign n28658 =  ( n28657 ) ? ( n4841 ) : ( iram_248 ) ;
assign n28659 = wr_addr[7:7] ;
assign n28660 =  ( n28659 ) == ( bv_1_0_n53 )  ;
assign n28661 =  ( wr_addr ) == ( bv_8_248_n565 )  ;
assign n28662 =  ( n28660 ) & (n28661 )  ;
assign n28663 =  ( n28662 ) & (wr )  ;
assign n28664 =  ( n28663 ) ? ( n5449 ) : ( iram_248 ) ;
assign n28665 = wr_addr[7:7] ;
assign n28666 =  ( n28665 ) == ( bv_1_0_n53 )  ;
assign n28667 =  ( wr_addr ) == ( bv_8_248_n565 )  ;
assign n28668 =  ( n28666 ) & (n28667 )  ;
assign n28669 =  ( n28668 ) & (wr )  ;
assign n28670 =  ( n28669 ) ? ( n4906 ) : ( iram_248 ) ;
assign n28671 = wr_addr[7:7] ;
assign n28672 =  ( n28671 ) == ( bv_1_0_n53 )  ;
assign n28673 =  ( wr_addr ) == ( bv_8_248_n565 )  ;
assign n28674 =  ( n28672 ) & (n28673 )  ;
assign n28675 =  ( n28674 ) & (wr )  ;
assign n28676 =  ( n28675 ) ? ( n5485 ) : ( iram_248 ) ;
assign n28677 = wr_addr[7:7] ;
assign n28678 =  ( n28677 ) == ( bv_1_0_n53 )  ;
assign n28679 =  ( wr_addr ) == ( bv_8_248_n565 )  ;
assign n28680 =  ( n28678 ) & (n28679 )  ;
assign n28681 =  ( n28680 ) & (wr )  ;
assign n28682 =  ( n28681 ) ? ( n5512 ) : ( iram_248 ) ;
assign n28683 = wr_addr[7:7] ;
assign n28684 =  ( n28683 ) == ( bv_1_0_n53 )  ;
assign n28685 =  ( wr_addr ) == ( bv_8_248_n565 )  ;
assign n28686 =  ( n28684 ) & (n28685 )  ;
assign n28687 =  ( n28686 ) & (wr )  ;
assign n28688 =  ( n28687 ) ? ( bv_8_0_n69 ) : ( iram_248 ) ;
assign n28689 = wr_addr[7:7] ;
assign n28690 =  ( n28689 ) == ( bv_1_0_n53 )  ;
assign n28691 =  ( wr_addr ) == ( bv_8_248_n565 )  ;
assign n28692 =  ( n28690 ) & (n28691 )  ;
assign n28693 =  ( n28692 ) & (wr )  ;
assign n28694 =  ( n28693 ) ? ( n5071 ) : ( iram_248 ) ;
assign n28695 = wr_addr[7:7] ;
assign n28696 =  ( n28695 ) == ( bv_1_0_n53 )  ;
assign n28697 =  ( wr_addr ) == ( bv_8_248_n565 )  ;
assign n28698 =  ( n28696 ) & (n28697 )  ;
assign n28699 =  ( n28698 ) & (wr )  ;
assign n28700 =  ( n28699 ) ? ( n5096 ) : ( iram_248 ) ;
assign n28701 = wr_addr[7:7] ;
assign n28702 =  ( n28701 ) == ( bv_1_0_n53 )  ;
assign n28703 =  ( wr_addr ) == ( bv_8_248_n565 )  ;
assign n28704 =  ( n28702 ) & (n28703 )  ;
assign n28705 =  ( n28704 ) & (wr )  ;
assign n28706 =  ( n28705 ) ? ( n5123 ) : ( iram_248 ) ;
assign n28707 = wr_addr[7:7] ;
assign n28708 =  ( n28707 ) == ( bv_1_0_n53 )  ;
assign n28709 =  ( wr_addr ) == ( bv_8_248_n565 )  ;
assign n28710 =  ( n28708 ) & (n28709 )  ;
assign n28711 =  ( n28710 ) & (wr )  ;
assign n28712 =  ( n28711 ) ? ( n5165 ) : ( iram_248 ) ;
assign n28713 = wr_addr[7:7] ;
assign n28714 =  ( n28713 ) == ( bv_1_0_n53 )  ;
assign n28715 =  ( wr_addr ) == ( bv_8_248_n565 )  ;
assign n28716 =  ( n28714 ) & (n28715 )  ;
assign n28717 =  ( n28716 ) & (wr )  ;
assign n28718 =  ( n28717 ) ? ( n5204 ) : ( iram_248 ) ;
assign n28719 = wr_addr[7:7] ;
assign n28720 =  ( n28719 ) == ( bv_1_0_n53 )  ;
assign n28721 =  ( wr_addr ) == ( bv_8_248_n565 )  ;
assign n28722 =  ( n28720 ) & (n28721 )  ;
assign n28723 =  ( n28722 ) & (wr )  ;
assign n28724 =  ( n28723 ) ? ( n5262 ) : ( iram_248 ) ;
assign n28725 = wr_addr[7:7] ;
assign n28726 =  ( n28725 ) == ( bv_1_0_n53 )  ;
assign n28727 =  ( wr_addr ) == ( bv_8_248_n565 )  ;
assign n28728 =  ( n28726 ) & (n28727 )  ;
assign n28729 =  ( n28728 ) & (wr )  ;
assign n28730 =  ( n28729 ) ? ( n5298 ) : ( iram_248 ) ;
assign n28731 = wr_addr[7:7] ;
assign n28732 =  ( n28731 ) == ( bv_1_0_n53 )  ;
assign n28733 =  ( wr_addr ) == ( bv_8_248_n565 )  ;
assign n28734 =  ( n28732 ) & (n28733 )  ;
assign n28735 =  ( n28734 ) & (wr )  ;
assign n28736 =  ( n28735 ) ? ( n5325 ) : ( iram_248 ) ;
assign n28737 = wr_addr[7:7] ;
assign n28738 =  ( n28737 ) == ( bv_1_0_n53 )  ;
assign n28739 =  ( wr_addr ) == ( bv_8_249_n567 )  ;
assign n28740 =  ( n28738 ) & (n28739 )  ;
assign n28741 =  ( n28740 ) & (wr )  ;
assign n28742 =  ( n28741 ) ? ( n4782 ) : ( iram_249 ) ;
assign n28743 = wr_addr[7:7] ;
assign n28744 =  ( n28743 ) == ( bv_1_0_n53 )  ;
assign n28745 =  ( wr_addr ) == ( bv_8_249_n567 )  ;
assign n28746 =  ( n28744 ) & (n28745 )  ;
assign n28747 =  ( n28746 ) & (wr )  ;
assign n28748 =  ( n28747 ) ? ( n4841 ) : ( iram_249 ) ;
assign n28749 = wr_addr[7:7] ;
assign n28750 =  ( n28749 ) == ( bv_1_0_n53 )  ;
assign n28751 =  ( wr_addr ) == ( bv_8_249_n567 )  ;
assign n28752 =  ( n28750 ) & (n28751 )  ;
assign n28753 =  ( n28752 ) & (wr )  ;
assign n28754 =  ( n28753 ) ? ( n5449 ) : ( iram_249 ) ;
assign n28755 = wr_addr[7:7] ;
assign n28756 =  ( n28755 ) == ( bv_1_0_n53 )  ;
assign n28757 =  ( wr_addr ) == ( bv_8_249_n567 )  ;
assign n28758 =  ( n28756 ) & (n28757 )  ;
assign n28759 =  ( n28758 ) & (wr )  ;
assign n28760 =  ( n28759 ) ? ( n4906 ) : ( iram_249 ) ;
assign n28761 = wr_addr[7:7] ;
assign n28762 =  ( n28761 ) == ( bv_1_0_n53 )  ;
assign n28763 =  ( wr_addr ) == ( bv_8_249_n567 )  ;
assign n28764 =  ( n28762 ) & (n28763 )  ;
assign n28765 =  ( n28764 ) & (wr )  ;
assign n28766 =  ( n28765 ) ? ( n5485 ) : ( iram_249 ) ;
assign n28767 = wr_addr[7:7] ;
assign n28768 =  ( n28767 ) == ( bv_1_0_n53 )  ;
assign n28769 =  ( wr_addr ) == ( bv_8_249_n567 )  ;
assign n28770 =  ( n28768 ) & (n28769 )  ;
assign n28771 =  ( n28770 ) & (wr )  ;
assign n28772 =  ( n28771 ) ? ( n5512 ) : ( iram_249 ) ;
assign n28773 = wr_addr[7:7] ;
assign n28774 =  ( n28773 ) == ( bv_1_0_n53 )  ;
assign n28775 =  ( wr_addr ) == ( bv_8_249_n567 )  ;
assign n28776 =  ( n28774 ) & (n28775 )  ;
assign n28777 =  ( n28776 ) & (wr )  ;
assign n28778 =  ( n28777 ) ? ( bv_8_0_n69 ) : ( iram_249 ) ;
assign n28779 = wr_addr[7:7] ;
assign n28780 =  ( n28779 ) == ( bv_1_0_n53 )  ;
assign n28781 =  ( wr_addr ) == ( bv_8_249_n567 )  ;
assign n28782 =  ( n28780 ) & (n28781 )  ;
assign n28783 =  ( n28782 ) & (wr )  ;
assign n28784 =  ( n28783 ) ? ( n5071 ) : ( iram_249 ) ;
assign n28785 = wr_addr[7:7] ;
assign n28786 =  ( n28785 ) == ( bv_1_0_n53 )  ;
assign n28787 =  ( wr_addr ) == ( bv_8_249_n567 )  ;
assign n28788 =  ( n28786 ) & (n28787 )  ;
assign n28789 =  ( n28788 ) & (wr )  ;
assign n28790 =  ( n28789 ) ? ( n5096 ) : ( iram_249 ) ;
assign n28791 = wr_addr[7:7] ;
assign n28792 =  ( n28791 ) == ( bv_1_0_n53 )  ;
assign n28793 =  ( wr_addr ) == ( bv_8_249_n567 )  ;
assign n28794 =  ( n28792 ) & (n28793 )  ;
assign n28795 =  ( n28794 ) & (wr )  ;
assign n28796 =  ( n28795 ) ? ( n5123 ) : ( iram_249 ) ;
assign n28797 = wr_addr[7:7] ;
assign n28798 =  ( n28797 ) == ( bv_1_0_n53 )  ;
assign n28799 =  ( wr_addr ) == ( bv_8_249_n567 )  ;
assign n28800 =  ( n28798 ) & (n28799 )  ;
assign n28801 =  ( n28800 ) & (wr )  ;
assign n28802 =  ( n28801 ) ? ( n5165 ) : ( iram_249 ) ;
assign n28803 = wr_addr[7:7] ;
assign n28804 =  ( n28803 ) == ( bv_1_0_n53 )  ;
assign n28805 =  ( wr_addr ) == ( bv_8_249_n567 )  ;
assign n28806 =  ( n28804 ) & (n28805 )  ;
assign n28807 =  ( n28806 ) & (wr )  ;
assign n28808 =  ( n28807 ) ? ( n5204 ) : ( iram_249 ) ;
assign n28809 = wr_addr[7:7] ;
assign n28810 =  ( n28809 ) == ( bv_1_0_n53 )  ;
assign n28811 =  ( wr_addr ) == ( bv_8_249_n567 )  ;
assign n28812 =  ( n28810 ) & (n28811 )  ;
assign n28813 =  ( n28812 ) & (wr )  ;
assign n28814 =  ( n28813 ) ? ( n5262 ) : ( iram_249 ) ;
assign n28815 = wr_addr[7:7] ;
assign n28816 =  ( n28815 ) == ( bv_1_0_n53 )  ;
assign n28817 =  ( wr_addr ) == ( bv_8_249_n567 )  ;
assign n28818 =  ( n28816 ) & (n28817 )  ;
assign n28819 =  ( n28818 ) & (wr )  ;
assign n28820 =  ( n28819 ) ? ( n5298 ) : ( iram_249 ) ;
assign n28821 = wr_addr[7:7] ;
assign n28822 =  ( n28821 ) == ( bv_1_0_n53 )  ;
assign n28823 =  ( wr_addr ) == ( bv_8_249_n567 )  ;
assign n28824 =  ( n28822 ) & (n28823 )  ;
assign n28825 =  ( n28824 ) & (wr )  ;
assign n28826 =  ( n28825 ) ? ( n5325 ) : ( iram_249 ) ;
assign n28827 = wr_addr[7:7] ;
assign n28828 =  ( n28827 ) == ( bv_1_0_n53 )  ;
assign n28829 =  ( wr_addr ) == ( bv_8_250_n569 )  ;
assign n28830 =  ( n28828 ) & (n28829 )  ;
assign n28831 =  ( n28830 ) & (wr )  ;
assign n28832 =  ( n28831 ) ? ( n4782 ) : ( iram_250 ) ;
assign n28833 = wr_addr[7:7] ;
assign n28834 =  ( n28833 ) == ( bv_1_0_n53 )  ;
assign n28835 =  ( wr_addr ) == ( bv_8_250_n569 )  ;
assign n28836 =  ( n28834 ) & (n28835 )  ;
assign n28837 =  ( n28836 ) & (wr )  ;
assign n28838 =  ( n28837 ) ? ( n4841 ) : ( iram_250 ) ;
assign n28839 = wr_addr[7:7] ;
assign n28840 =  ( n28839 ) == ( bv_1_0_n53 )  ;
assign n28841 =  ( wr_addr ) == ( bv_8_250_n569 )  ;
assign n28842 =  ( n28840 ) & (n28841 )  ;
assign n28843 =  ( n28842 ) & (wr )  ;
assign n28844 =  ( n28843 ) ? ( n5449 ) : ( iram_250 ) ;
assign n28845 = wr_addr[7:7] ;
assign n28846 =  ( n28845 ) == ( bv_1_0_n53 )  ;
assign n28847 =  ( wr_addr ) == ( bv_8_250_n569 )  ;
assign n28848 =  ( n28846 ) & (n28847 )  ;
assign n28849 =  ( n28848 ) & (wr )  ;
assign n28850 =  ( n28849 ) ? ( n4906 ) : ( iram_250 ) ;
assign n28851 = wr_addr[7:7] ;
assign n28852 =  ( n28851 ) == ( bv_1_0_n53 )  ;
assign n28853 =  ( wr_addr ) == ( bv_8_250_n569 )  ;
assign n28854 =  ( n28852 ) & (n28853 )  ;
assign n28855 =  ( n28854 ) & (wr )  ;
assign n28856 =  ( n28855 ) ? ( n5485 ) : ( iram_250 ) ;
assign n28857 = wr_addr[7:7] ;
assign n28858 =  ( n28857 ) == ( bv_1_0_n53 )  ;
assign n28859 =  ( wr_addr ) == ( bv_8_250_n569 )  ;
assign n28860 =  ( n28858 ) & (n28859 )  ;
assign n28861 =  ( n28860 ) & (wr )  ;
assign n28862 =  ( n28861 ) ? ( n5512 ) : ( iram_250 ) ;
assign n28863 = wr_addr[7:7] ;
assign n28864 =  ( n28863 ) == ( bv_1_0_n53 )  ;
assign n28865 =  ( wr_addr ) == ( bv_8_250_n569 )  ;
assign n28866 =  ( n28864 ) & (n28865 )  ;
assign n28867 =  ( n28866 ) & (wr )  ;
assign n28868 =  ( n28867 ) ? ( bv_8_0_n69 ) : ( iram_250 ) ;
assign n28869 = wr_addr[7:7] ;
assign n28870 =  ( n28869 ) == ( bv_1_0_n53 )  ;
assign n28871 =  ( wr_addr ) == ( bv_8_250_n569 )  ;
assign n28872 =  ( n28870 ) & (n28871 )  ;
assign n28873 =  ( n28872 ) & (wr )  ;
assign n28874 =  ( n28873 ) ? ( n5071 ) : ( iram_250 ) ;
assign n28875 = wr_addr[7:7] ;
assign n28876 =  ( n28875 ) == ( bv_1_0_n53 )  ;
assign n28877 =  ( wr_addr ) == ( bv_8_250_n569 )  ;
assign n28878 =  ( n28876 ) & (n28877 )  ;
assign n28879 =  ( n28878 ) & (wr )  ;
assign n28880 =  ( n28879 ) ? ( n5096 ) : ( iram_250 ) ;
assign n28881 = wr_addr[7:7] ;
assign n28882 =  ( n28881 ) == ( bv_1_0_n53 )  ;
assign n28883 =  ( wr_addr ) == ( bv_8_250_n569 )  ;
assign n28884 =  ( n28882 ) & (n28883 )  ;
assign n28885 =  ( n28884 ) & (wr )  ;
assign n28886 =  ( n28885 ) ? ( n5123 ) : ( iram_250 ) ;
assign n28887 = wr_addr[7:7] ;
assign n28888 =  ( n28887 ) == ( bv_1_0_n53 )  ;
assign n28889 =  ( wr_addr ) == ( bv_8_250_n569 )  ;
assign n28890 =  ( n28888 ) & (n28889 )  ;
assign n28891 =  ( n28890 ) & (wr )  ;
assign n28892 =  ( n28891 ) ? ( n5165 ) : ( iram_250 ) ;
assign n28893 = wr_addr[7:7] ;
assign n28894 =  ( n28893 ) == ( bv_1_0_n53 )  ;
assign n28895 =  ( wr_addr ) == ( bv_8_250_n569 )  ;
assign n28896 =  ( n28894 ) & (n28895 )  ;
assign n28897 =  ( n28896 ) & (wr )  ;
assign n28898 =  ( n28897 ) ? ( n5204 ) : ( iram_250 ) ;
assign n28899 = wr_addr[7:7] ;
assign n28900 =  ( n28899 ) == ( bv_1_0_n53 )  ;
assign n28901 =  ( wr_addr ) == ( bv_8_250_n569 )  ;
assign n28902 =  ( n28900 ) & (n28901 )  ;
assign n28903 =  ( n28902 ) & (wr )  ;
assign n28904 =  ( n28903 ) ? ( n5262 ) : ( iram_250 ) ;
assign n28905 = wr_addr[7:7] ;
assign n28906 =  ( n28905 ) == ( bv_1_0_n53 )  ;
assign n28907 =  ( wr_addr ) == ( bv_8_250_n569 )  ;
assign n28908 =  ( n28906 ) & (n28907 )  ;
assign n28909 =  ( n28908 ) & (wr )  ;
assign n28910 =  ( n28909 ) ? ( n5298 ) : ( iram_250 ) ;
assign n28911 = wr_addr[7:7] ;
assign n28912 =  ( n28911 ) == ( bv_1_0_n53 )  ;
assign n28913 =  ( wr_addr ) == ( bv_8_250_n569 )  ;
assign n28914 =  ( n28912 ) & (n28913 )  ;
assign n28915 =  ( n28914 ) & (wr )  ;
assign n28916 =  ( n28915 ) ? ( n5325 ) : ( iram_250 ) ;
assign n28917 = wr_addr[7:7] ;
assign n28918 =  ( n28917 ) == ( bv_1_0_n53 )  ;
assign n28919 =  ( wr_addr ) == ( bv_8_251_n571 )  ;
assign n28920 =  ( n28918 ) & (n28919 )  ;
assign n28921 =  ( n28920 ) & (wr )  ;
assign n28922 =  ( n28921 ) ? ( n4782 ) : ( iram_251 ) ;
assign n28923 = wr_addr[7:7] ;
assign n28924 =  ( n28923 ) == ( bv_1_0_n53 )  ;
assign n28925 =  ( wr_addr ) == ( bv_8_251_n571 )  ;
assign n28926 =  ( n28924 ) & (n28925 )  ;
assign n28927 =  ( n28926 ) & (wr )  ;
assign n28928 =  ( n28927 ) ? ( n4841 ) : ( iram_251 ) ;
assign n28929 = wr_addr[7:7] ;
assign n28930 =  ( n28929 ) == ( bv_1_0_n53 )  ;
assign n28931 =  ( wr_addr ) == ( bv_8_251_n571 )  ;
assign n28932 =  ( n28930 ) & (n28931 )  ;
assign n28933 =  ( n28932 ) & (wr )  ;
assign n28934 =  ( n28933 ) ? ( n5449 ) : ( iram_251 ) ;
assign n28935 = wr_addr[7:7] ;
assign n28936 =  ( n28935 ) == ( bv_1_0_n53 )  ;
assign n28937 =  ( wr_addr ) == ( bv_8_251_n571 )  ;
assign n28938 =  ( n28936 ) & (n28937 )  ;
assign n28939 =  ( n28938 ) & (wr )  ;
assign n28940 =  ( n28939 ) ? ( n4906 ) : ( iram_251 ) ;
assign n28941 = wr_addr[7:7] ;
assign n28942 =  ( n28941 ) == ( bv_1_0_n53 )  ;
assign n28943 =  ( wr_addr ) == ( bv_8_251_n571 )  ;
assign n28944 =  ( n28942 ) & (n28943 )  ;
assign n28945 =  ( n28944 ) & (wr )  ;
assign n28946 =  ( n28945 ) ? ( n5485 ) : ( iram_251 ) ;
assign n28947 = wr_addr[7:7] ;
assign n28948 =  ( n28947 ) == ( bv_1_0_n53 )  ;
assign n28949 =  ( wr_addr ) == ( bv_8_251_n571 )  ;
assign n28950 =  ( n28948 ) & (n28949 )  ;
assign n28951 =  ( n28950 ) & (wr )  ;
assign n28952 =  ( n28951 ) ? ( n5512 ) : ( iram_251 ) ;
assign n28953 = wr_addr[7:7] ;
assign n28954 =  ( n28953 ) == ( bv_1_0_n53 )  ;
assign n28955 =  ( wr_addr ) == ( bv_8_251_n571 )  ;
assign n28956 =  ( n28954 ) & (n28955 )  ;
assign n28957 =  ( n28956 ) & (wr )  ;
assign n28958 =  ( n28957 ) ? ( bv_8_0_n69 ) : ( iram_251 ) ;
assign n28959 = wr_addr[7:7] ;
assign n28960 =  ( n28959 ) == ( bv_1_0_n53 )  ;
assign n28961 =  ( wr_addr ) == ( bv_8_251_n571 )  ;
assign n28962 =  ( n28960 ) & (n28961 )  ;
assign n28963 =  ( n28962 ) & (wr )  ;
assign n28964 =  ( n28963 ) ? ( n5071 ) : ( iram_251 ) ;
assign n28965 = wr_addr[7:7] ;
assign n28966 =  ( n28965 ) == ( bv_1_0_n53 )  ;
assign n28967 =  ( wr_addr ) == ( bv_8_251_n571 )  ;
assign n28968 =  ( n28966 ) & (n28967 )  ;
assign n28969 =  ( n28968 ) & (wr )  ;
assign n28970 =  ( n28969 ) ? ( n5096 ) : ( iram_251 ) ;
assign n28971 = wr_addr[7:7] ;
assign n28972 =  ( n28971 ) == ( bv_1_0_n53 )  ;
assign n28973 =  ( wr_addr ) == ( bv_8_251_n571 )  ;
assign n28974 =  ( n28972 ) & (n28973 )  ;
assign n28975 =  ( n28974 ) & (wr )  ;
assign n28976 =  ( n28975 ) ? ( n5123 ) : ( iram_251 ) ;
assign n28977 = wr_addr[7:7] ;
assign n28978 =  ( n28977 ) == ( bv_1_0_n53 )  ;
assign n28979 =  ( wr_addr ) == ( bv_8_251_n571 )  ;
assign n28980 =  ( n28978 ) & (n28979 )  ;
assign n28981 =  ( n28980 ) & (wr )  ;
assign n28982 =  ( n28981 ) ? ( n5165 ) : ( iram_251 ) ;
assign n28983 = wr_addr[7:7] ;
assign n28984 =  ( n28983 ) == ( bv_1_0_n53 )  ;
assign n28985 =  ( wr_addr ) == ( bv_8_251_n571 )  ;
assign n28986 =  ( n28984 ) & (n28985 )  ;
assign n28987 =  ( n28986 ) & (wr )  ;
assign n28988 =  ( n28987 ) ? ( n5204 ) : ( iram_251 ) ;
assign n28989 = wr_addr[7:7] ;
assign n28990 =  ( n28989 ) == ( bv_1_0_n53 )  ;
assign n28991 =  ( wr_addr ) == ( bv_8_251_n571 )  ;
assign n28992 =  ( n28990 ) & (n28991 )  ;
assign n28993 =  ( n28992 ) & (wr )  ;
assign n28994 =  ( n28993 ) ? ( n5262 ) : ( iram_251 ) ;
assign n28995 = wr_addr[7:7] ;
assign n28996 =  ( n28995 ) == ( bv_1_0_n53 )  ;
assign n28997 =  ( wr_addr ) == ( bv_8_251_n571 )  ;
assign n28998 =  ( n28996 ) & (n28997 )  ;
assign n28999 =  ( n28998 ) & (wr )  ;
assign n29000 =  ( n28999 ) ? ( n5298 ) : ( iram_251 ) ;
assign n29001 = wr_addr[7:7] ;
assign n29002 =  ( n29001 ) == ( bv_1_0_n53 )  ;
assign n29003 =  ( wr_addr ) == ( bv_8_251_n571 )  ;
assign n29004 =  ( n29002 ) & (n29003 )  ;
assign n29005 =  ( n29004 ) & (wr )  ;
assign n29006 =  ( n29005 ) ? ( n5325 ) : ( iram_251 ) ;
assign n29007 = wr_addr[7:7] ;
assign n29008 =  ( n29007 ) == ( bv_1_0_n53 )  ;
assign n29009 =  ( wr_addr ) == ( bv_8_252_n573 )  ;
assign n29010 =  ( n29008 ) & (n29009 )  ;
assign n29011 =  ( n29010 ) & (wr )  ;
assign n29012 =  ( n29011 ) ? ( n4782 ) : ( iram_252 ) ;
assign n29013 = wr_addr[7:7] ;
assign n29014 =  ( n29013 ) == ( bv_1_0_n53 )  ;
assign n29015 =  ( wr_addr ) == ( bv_8_252_n573 )  ;
assign n29016 =  ( n29014 ) & (n29015 )  ;
assign n29017 =  ( n29016 ) & (wr )  ;
assign n29018 =  ( n29017 ) ? ( n4841 ) : ( iram_252 ) ;
assign n29019 = wr_addr[7:7] ;
assign n29020 =  ( n29019 ) == ( bv_1_0_n53 )  ;
assign n29021 =  ( wr_addr ) == ( bv_8_252_n573 )  ;
assign n29022 =  ( n29020 ) & (n29021 )  ;
assign n29023 =  ( n29022 ) & (wr )  ;
assign n29024 =  ( n29023 ) ? ( n5449 ) : ( iram_252 ) ;
assign n29025 = wr_addr[7:7] ;
assign n29026 =  ( n29025 ) == ( bv_1_0_n53 )  ;
assign n29027 =  ( wr_addr ) == ( bv_8_252_n573 )  ;
assign n29028 =  ( n29026 ) & (n29027 )  ;
assign n29029 =  ( n29028 ) & (wr )  ;
assign n29030 =  ( n29029 ) ? ( n4906 ) : ( iram_252 ) ;
assign n29031 = wr_addr[7:7] ;
assign n29032 =  ( n29031 ) == ( bv_1_0_n53 )  ;
assign n29033 =  ( wr_addr ) == ( bv_8_252_n573 )  ;
assign n29034 =  ( n29032 ) & (n29033 )  ;
assign n29035 =  ( n29034 ) & (wr )  ;
assign n29036 =  ( n29035 ) ? ( n5485 ) : ( iram_252 ) ;
assign n29037 = wr_addr[7:7] ;
assign n29038 =  ( n29037 ) == ( bv_1_0_n53 )  ;
assign n29039 =  ( wr_addr ) == ( bv_8_252_n573 )  ;
assign n29040 =  ( n29038 ) & (n29039 )  ;
assign n29041 =  ( n29040 ) & (wr )  ;
assign n29042 =  ( n29041 ) ? ( n5512 ) : ( iram_252 ) ;
assign n29043 = wr_addr[7:7] ;
assign n29044 =  ( n29043 ) == ( bv_1_0_n53 )  ;
assign n29045 =  ( wr_addr ) == ( bv_8_252_n573 )  ;
assign n29046 =  ( n29044 ) & (n29045 )  ;
assign n29047 =  ( n29046 ) & (wr )  ;
assign n29048 =  ( n29047 ) ? ( bv_8_0_n69 ) : ( iram_252 ) ;
assign n29049 = wr_addr[7:7] ;
assign n29050 =  ( n29049 ) == ( bv_1_0_n53 )  ;
assign n29051 =  ( wr_addr ) == ( bv_8_252_n573 )  ;
assign n29052 =  ( n29050 ) & (n29051 )  ;
assign n29053 =  ( n29052 ) & (wr )  ;
assign n29054 =  ( n29053 ) ? ( n5071 ) : ( iram_252 ) ;
assign n29055 = wr_addr[7:7] ;
assign n29056 =  ( n29055 ) == ( bv_1_0_n53 )  ;
assign n29057 =  ( wr_addr ) == ( bv_8_252_n573 )  ;
assign n29058 =  ( n29056 ) & (n29057 )  ;
assign n29059 =  ( n29058 ) & (wr )  ;
assign n29060 =  ( n29059 ) ? ( n5096 ) : ( iram_252 ) ;
assign n29061 = wr_addr[7:7] ;
assign n29062 =  ( n29061 ) == ( bv_1_0_n53 )  ;
assign n29063 =  ( wr_addr ) == ( bv_8_252_n573 )  ;
assign n29064 =  ( n29062 ) & (n29063 )  ;
assign n29065 =  ( n29064 ) & (wr )  ;
assign n29066 =  ( n29065 ) ? ( n5123 ) : ( iram_252 ) ;
assign n29067 = wr_addr[7:7] ;
assign n29068 =  ( n29067 ) == ( bv_1_0_n53 )  ;
assign n29069 =  ( wr_addr ) == ( bv_8_252_n573 )  ;
assign n29070 =  ( n29068 ) & (n29069 )  ;
assign n29071 =  ( n29070 ) & (wr )  ;
assign n29072 =  ( n29071 ) ? ( n5165 ) : ( iram_252 ) ;
assign n29073 = wr_addr[7:7] ;
assign n29074 =  ( n29073 ) == ( bv_1_0_n53 )  ;
assign n29075 =  ( wr_addr ) == ( bv_8_252_n573 )  ;
assign n29076 =  ( n29074 ) & (n29075 )  ;
assign n29077 =  ( n29076 ) & (wr )  ;
assign n29078 =  ( n29077 ) ? ( n5204 ) : ( iram_252 ) ;
assign n29079 = wr_addr[7:7] ;
assign n29080 =  ( n29079 ) == ( bv_1_0_n53 )  ;
assign n29081 =  ( wr_addr ) == ( bv_8_252_n573 )  ;
assign n29082 =  ( n29080 ) & (n29081 )  ;
assign n29083 =  ( n29082 ) & (wr )  ;
assign n29084 =  ( n29083 ) ? ( n5262 ) : ( iram_252 ) ;
assign n29085 = wr_addr[7:7] ;
assign n29086 =  ( n29085 ) == ( bv_1_0_n53 )  ;
assign n29087 =  ( wr_addr ) == ( bv_8_252_n573 )  ;
assign n29088 =  ( n29086 ) & (n29087 )  ;
assign n29089 =  ( n29088 ) & (wr )  ;
assign n29090 =  ( n29089 ) ? ( n5298 ) : ( iram_252 ) ;
assign n29091 = wr_addr[7:7] ;
assign n29092 =  ( n29091 ) == ( bv_1_0_n53 )  ;
assign n29093 =  ( wr_addr ) == ( bv_8_252_n573 )  ;
assign n29094 =  ( n29092 ) & (n29093 )  ;
assign n29095 =  ( n29094 ) & (wr )  ;
assign n29096 =  ( n29095 ) ? ( n5325 ) : ( iram_252 ) ;
assign n29097 = wr_addr[7:7] ;
assign n29098 =  ( n29097 ) == ( bv_1_0_n53 )  ;
assign n29099 =  ( wr_addr ) == ( bv_8_253_n575 )  ;
assign n29100 =  ( n29098 ) & (n29099 )  ;
assign n29101 =  ( n29100 ) & (wr )  ;
assign n29102 =  ( n29101 ) ? ( n4782 ) : ( iram_253 ) ;
assign n29103 = wr_addr[7:7] ;
assign n29104 =  ( n29103 ) == ( bv_1_0_n53 )  ;
assign n29105 =  ( wr_addr ) == ( bv_8_253_n575 )  ;
assign n29106 =  ( n29104 ) & (n29105 )  ;
assign n29107 =  ( n29106 ) & (wr )  ;
assign n29108 =  ( n29107 ) ? ( n4841 ) : ( iram_253 ) ;
assign n29109 = wr_addr[7:7] ;
assign n29110 =  ( n29109 ) == ( bv_1_0_n53 )  ;
assign n29111 =  ( wr_addr ) == ( bv_8_253_n575 )  ;
assign n29112 =  ( n29110 ) & (n29111 )  ;
assign n29113 =  ( n29112 ) & (wr )  ;
assign n29114 =  ( n29113 ) ? ( n5449 ) : ( iram_253 ) ;
assign n29115 = wr_addr[7:7] ;
assign n29116 =  ( n29115 ) == ( bv_1_0_n53 )  ;
assign n29117 =  ( wr_addr ) == ( bv_8_253_n575 )  ;
assign n29118 =  ( n29116 ) & (n29117 )  ;
assign n29119 =  ( n29118 ) & (wr )  ;
assign n29120 =  ( n29119 ) ? ( n4906 ) : ( iram_253 ) ;
assign n29121 = wr_addr[7:7] ;
assign n29122 =  ( n29121 ) == ( bv_1_0_n53 )  ;
assign n29123 =  ( wr_addr ) == ( bv_8_253_n575 )  ;
assign n29124 =  ( n29122 ) & (n29123 )  ;
assign n29125 =  ( n29124 ) & (wr )  ;
assign n29126 =  ( n29125 ) ? ( n5485 ) : ( iram_253 ) ;
assign n29127 = wr_addr[7:7] ;
assign n29128 =  ( n29127 ) == ( bv_1_0_n53 )  ;
assign n29129 =  ( wr_addr ) == ( bv_8_253_n575 )  ;
assign n29130 =  ( n29128 ) & (n29129 )  ;
assign n29131 =  ( n29130 ) & (wr )  ;
assign n29132 =  ( n29131 ) ? ( n5512 ) : ( iram_253 ) ;
assign n29133 = wr_addr[7:7] ;
assign n29134 =  ( n29133 ) == ( bv_1_0_n53 )  ;
assign n29135 =  ( wr_addr ) == ( bv_8_253_n575 )  ;
assign n29136 =  ( n29134 ) & (n29135 )  ;
assign n29137 =  ( n29136 ) & (wr )  ;
assign n29138 =  ( n29137 ) ? ( bv_8_0_n69 ) : ( iram_253 ) ;
assign n29139 = wr_addr[7:7] ;
assign n29140 =  ( n29139 ) == ( bv_1_0_n53 )  ;
assign n29141 =  ( wr_addr ) == ( bv_8_253_n575 )  ;
assign n29142 =  ( n29140 ) & (n29141 )  ;
assign n29143 =  ( n29142 ) & (wr )  ;
assign n29144 =  ( n29143 ) ? ( n5071 ) : ( iram_253 ) ;
assign n29145 = wr_addr[7:7] ;
assign n29146 =  ( n29145 ) == ( bv_1_0_n53 )  ;
assign n29147 =  ( wr_addr ) == ( bv_8_253_n575 )  ;
assign n29148 =  ( n29146 ) & (n29147 )  ;
assign n29149 =  ( n29148 ) & (wr )  ;
assign n29150 =  ( n29149 ) ? ( n5096 ) : ( iram_253 ) ;
assign n29151 = wr_addr[7:7] ;
assign n29152 =  ( n29151 ) == ( bv_1_0_n53 )  ;
assign n29153 =  ( wr_addr ) == ( bv_8_253_n575 )  ;
assign n29154 =  ( n29152 ) & (n29153 )  ;
assign n29155 =  ( n29154 ) & (wr )  ;
assign n29156 =  ( n29155 ) ? ( n5123 ) : ( iram_253 ) ;
assign n29157 = wr_addr[7:7] ;
assign n29158 =  ( n29157 ) == ( bv_1_0_n53 )  ;
assign n29159 =  ( wr_addr ) == ( bv_8_253_n575 )  ;
assign n29160 =  ( n29158 ) & (n29159 )  ;
assign n29161 =  ( n29160 ) & (wr )  ;
assign n29162 =  ( n29161 ) ? ( n5165 ) : ( iram_253 ) ;
assign n29163 = wr_addr[7:7] ;
assign n29164 =  ( n29163 ) == ( bv_1_0_n53 )  ;
assign n29165 =  ( wr_addr ) == ( bv_8_253_n575 )  ;
assign n29166 =  ( n29164 ) & (n29165 )  ;
assign n29167 =  ( n29166 ) & (wr )  ;
assign n29168 =  ( n29167 ) ? ( n5204 ) : ( iram_253 ) ;
assign n29169 = wr_addr[7:7] ;
assign n29170 =  ( n29169 ) == ( bv_1_0_n53 )  ;
assign n29171 =  ( wr_addr ) == ( bv_8_253_n575 )  ;
assign n29172 =  ( n29170 ) & (n29171 )  ;
assign n29173 =  ( n29172 ) & (wr )  ;
assign n29174 =  ( n29173 ) ? ( n5262 ) : ( iram_253 ) ;
assign n29175 = wr_addr[7:7] ;
assign n29176 =  ( n29175 ) == ( bv_1_0_n53 )  ;
assign n29177 =  ( wr_addr ) == ( bv_8_253_n575 )  ;
assign n29178 =  ( n29176 ) & (n29177 )  ;
assign n29179 =  ( n29178 ) & (wr )  ;
assign n29180 =  ( n29179 ) ? ( n5298 ) : ( iram_253 ) ;
assign n29181 = wr_addr[7:7] ;
assign n29182 =  ( n29181 ) == ( bv_1_0_n53 )  ;
assign n29183 =  ( wr_addr ) == ( bv_8_253_n575 )  ;
assign n29184 =  ( n29182 ) & (n29183 )  ;
assign n29185 =  ( n29184 ) & (wr )  ;
assign n29186 =  ( n29185 ) ? ( n5325 ) : ( iram_253 ) ;
assign n29187 = wr_addr[7:7] ;
assign n29188 =  ( n29187 ) == ( bv_1_0_n53 )  ;
assign n29189 =  ( wr_addr ) == ( bv_8_254_n577 )  ;
assign n29190 =  ( n29188 ) & (n29189 )  ;
assign n29191 =  ( n29190 ) & (wr )  ;
assign n29192 =  ( n29191 ) ? ( n4782 ) : ( iram_254 ) ;
assign n29193 = wr_addr[7:7] ;
assign n29194 =  ( n29193 ) == ( bv_1_0_n53 )  ;
assign n29195 =  ( wr_addr ) == ( bv_8_254_n577 )  ;
assign n29196 =  ( n29194 ) & (n29195 )  ;
assign n29197 =  ( n29196 ) & (wr )  ;
assign n29198 =  ( n29197 ) ? ( n4841 ) : ( iram_254 ) ;
assign n29199 = wr_addr[7:7] ;
assign n29200 =  ( n29199 ) == ( bv_1_0_n53 )  ;
assign n29201 =  ( wr_addr ) == ( bv_8_254_n577 )  ;
assign n29202 =  ( n29200 ) & (n29201 )  ;
assign n29203 =  ( n29202 ) & (wr )  ;
assign n29204 =  ( n29203 ) ? ( n5449 ) : ( iram_254 ) ;
assign n29205 = wr_addr[7:7] ;
assign n29206 =  ( n29205 ) == ( bv_1_0_n53 )  ;
assign n29207 =  ( wr_addr ) == ( bv_8_254_n577 )  ;
assign n29208 =  ( n29206 ) & (n29207 )  ;
assign n29209 =  ( n29208 ) & (wr )  ;
assign n29210 =  ( n29209 ) ? ( n4906 ) : ( iram_254 ) ;
assign n29211 = wr_addr[7:7] ;
assign n29212 =  ( n29211 ) == ( bv_1_0_n53 )  ;
assign n29213 =  ( wr_addr ) == ( bv_8_254_n577 )  ;
assign n29214 =  ( n29212 ) & (n29213 )  ;
assign n29215 =  ( n29214 ) & (wr )  ;
assign n29216 =  ( n29215 ) ? ( n5485 ) : ( iram_254 ) ;
assign n29217 = wr_addr[7:7] ;
assign n29218 =  ( n29217 ) == ( bv_1_0_n53 )  ;
assign n29219 =  ( wr_addr ) == ( bv_8_254_n577 )  ;
assign n29220 =  ( n29218 ) & (n29219 )  ;
assign n29221 =  ( n29220 ) & (wr )  ;
assign n29222 =  ( n29221 ) ? ( n5512 ) : ( iram_254 ) ;
assign n29223 = wr_addr[7:7] ;
assign n29224 =  ( n29223 ) == ( bv_1_0_n53 )  ;
assign n29225 =  ( wr_addr ) == ( bv_8_254_n577 )  ;
assign n29226 =  ( n29224 ) & (n29225 )  ;
assign n29227 =  ( n29226 ) & (wr )  ;
assign n29228 =  ( n29227 ) ? ( bv_8_0_n69 ) : ( iram_254 ) ;
assign n29229 = wr_addr[7:7] ;
assign n29230 =  ( n29229 ) == ( bv_1_0_n53 )  ;
assign n29231 =  ( wr_addr ) == ( bv_8_254_n577 )  ;
assign n29232 =  ( n29230 ) & (n29231 )  ;
assign n29233 =  ( n29232 ) & (wr )  ;
assign n29234 =  ( n29233 ) ? ( n5071 ) : ( iram_254 ) ;
assign n29235 = wr_addr[7:7] ;
assign n29236 =  ( n29235 ) == ( bv_1_0_n53 )  ;
assign n29237 =  ( wr_addr ) == ( bv_8_254_n577 )  ;
assign n29238 =  ( n29236 ) & (n29237 )  ;
assign n29239 =  ( n29238 ) & (wr )  ;
assign n29240 =  ( n29239 ) ? ( n5096 ) : ( iram_254 ) ;
assign n29241 = wr_addr[7:7] ;
assign n29242 =  ( n29241 ) == ( bv_1_0_n53 )  ;
assign n29243 =  ( wr_addr ) == ( bv_8_254_n577 )  ;
assign n29244 =  ( n29242 ) & (n29243 )  ;
assign n29245 =  ( n29244 ) & (wr )  ;
assign n29246 =  ( n29245 ) ? ( n5123 ) : ( iram_254 ) ;
assign n29247 = wr_addr[7:7] ;
assign n29248 =  ( n29247 ) == ( bv_1_0_n53 )  ;
assign n29249 =  ( wr_addr ) == ( bv_8_254_n577 )  ;
assign n29250 =  ( n29248 ) & (n29249 )  ;
assign n29251 =  ( n29250 ) & (wr )  ;
assign n29252 =  ( n29251 ) ? ( n5165 ) : ( iram_254 ) ;
assign n29253 = wr_addr[7:7] ;
assign n29254 =  ( n29253 ) == ( bv_1_0_n53 )  ;
assign n29255 =  ( wr_addr ) == ( bv_8_254_n577 )  ;
assign n29256 =  ( n29254 ) & (n29255 )  ;
assign n29257 =  ( n29256 ) & (wr )  ;
assign n29258 =  ( n29257 ) ? ( n5204 ) : ( iram_254 ) ;
assign n29259 = wr_addr[7:7] ;
assign n29260 =  ( n29259 ) == ( bv_1_0_n53 )  ;
assign n29261 =  ( wr_addr ) == ( bv_8_254_n577 )  ;
assign n29262 =  ( n29260 ) & (n29261 )  ;
assign n29263 =  ( n29262 ) & (wr )  ;
assign n29264 =  ( n29263 ) ? ( n5262 ) : ( iram_254 ) ;
assign n29265 = wr_addr[7:7] ;
assign n29266 =  ( n29265 ) == ( bv_1_0_n53 )  ;
assign n29267 =  ( wr_addr ) == ( bv_8_254_n577 )  ;
assign n29268 =  ( n29266 ) & (n29267 )  ;
assign n29269 =  ( n29268 ) & (wr )  ;
assign n29270 =  ( n29269 ) ? ( n5298 ) : ( iram_254 ) ;
assign n29271 = wr_addr[7:7] ;
assign n29272 =  ( n29271 ) == ( bv_1_0_n53 )  ;
assign n29273 =  ( wr_addr ) == ( bv_8_254_n577 )  ;
assign n29274 =  ( n29272 ) & (n29273 )  ;
assign n29275 =  ( n29274 ) & (wr )  ;
assign n29276 =  ( n29275 ) ? ( n5325 ) : ( iram_254 ) ;
assign n29277 = wr_addr[7:7] ;
assign n29278 =  ( n29277 ) == ( bv_1_0_n53 )  ;
assign bv_8_255_n29279 = 8'hff ;
assign n29280 =  ( wr_addr ) == ( bv_8_255_n29279 )  ;
assign n29281 =  ( n29278 ) & (n29280 )  ;
assign n29282 =  ( n29281 ) & (wr )  ;
assign n29283 =  ( n29282 ) ? ( n4782 ) : ( iram_255 ) ;
assign n29284 = wr_addr[7:7] ;
assign n29285 =  ( n29284 ) == ( bv_1_0_n53 )  ;
assign n29286 =  ( wr_addr ) == ( bv_8_255_n29279 )  ;
assign n29287 =  ( n29285 ) & (n29286 )  ;
assign n29288 =  ( n29287 ) & (wr )  ;
assign n29289 =  ( n29288 ) ? ( n4841 ) : ( iram_255 ) ;
assign n29290 = wr_addr[7:7] ;
assign n29291 =  ( n29290 ) == ( bv_1_0_n53 )  ;
assign n29292 =  ( wr_addr ) == ( bv_8_255_n29279 )  ;
assign n29293 =  ( n29291 ) & (n29292 )  ;
assign n29294 =  ( n29293 ) & (wr )  ;
assign n29295 =  ( n29294 ) ? ( n5449 ) : ( iram_255 ) ;
assign n29296 = wr_addr[7:7] ;
assign n29297 =  ( n29296 ) == ( bv_1_0_n53 )  ;
assign n29298 =  ( wr_addr ) == ( bv_8_255_n29279 )  ;
assign n29299 =  ( n29297 ) & (n29298 )  ;
assign n29300 =  ( n29299 ) & (wr )  ;
assign n29301 =  ( n29300 ) ? ( n4906 ) : ( iram_255 ) ;
assign n29302 = wr_addr[7:7] ;
assign n29303 =  ( n29302 ) == ( bv_1_0_n53 )  ;
assign n29304 =  ( wr_addr ) == ( bv_8_255_n29279 )  ;
assign n29305 =  ( n29303 ) & (n29304 )  ;
assign n29306 =  ( n29305 ) & (wr )  ;
assign n29307 =  ( n29306 ) ? ( n5485 ) : ( iram_255 ) ;
assign n29308 = wr_addr[7:7] ;
assign n29309 =  ( n29308 ) == ( bv_1_0_n53 )  ;
assign n29310 =  ( wr_addr ) == ( bv_8_255_n29279 )  ;
assign n29311 =  ( n29309 ) & (n29310 )  ;
assign n29312 =  ( n29311 ) & (wr )  ;
assign n29313 =  ( n29312 ) ? ( n5512 ) : ( iram_255 ) ;
assign n29314 = wr_addr[7:7] ;
assign n29315 =  ( n29314 ) == ( bv_1_0_n53 )  ;
assign n29316 =  ( wr_addr ) == ( bv_8_255_n29279 )  ;
assign n29317 =  ( n29315 ) & (n29316 )  ;
assign n29318 =  ( n29317 ) & (wr )  ;
assign n29319 =  ( n29318 ) ? ( bv_8_0_n69 ) : ( iram_255 ) ;
assign n29320 = wr_addr[7:7] ;
assign n29321 =  ( n29320 ) == ( bv_1_0_n53 )  ;
assign n29322 =  ( wr_addr ) == ( bv_8_255_n29279 )  ;
assign n29323 =  ( n29321 ) & (n29322 )  ;
assign n29324 =  ( n29323 ) & (wr )  ;
assign n29325 =  ( n29324 ) ? ( n5071 ) : ( iram_255 ) ;
assign n29326 = wr_addr[7:7] ;
assign n29327 =  ( n29326 ) == ( bv_1_0_n53 )  ;
assign n29328 =  ( wr_addr ) == ( bv_8_255_n29279 )  ;
assign n29329 =  ( n29327 ) & (n29328 )  ;
assign n29330 =  ( n29329 ) & (wr )  ;
assign n29331 =  ( n29330 ) ? ( n5096 ) : ( iram_255 ) ;
assign n29332 = wr_addr[7:7] ;
assign n29333 =  ( n29332 ) == ( bv_1_0_n53 )  ;
assign n29334 =  ( wr_addr ) == ( bv_8_255_n29279 )  ;
assign n29335 =  ( n29333 ) & (n29334 )  ;
assign n29336 =  ( n29335 ) & (wr )  ;
assign n29337 =  ( n29336 ) ? ( n5123 ) : ( iram_255 ) ;
assign n29338 = wr_addr[7:7] ;
assign n29339 =  ( n29338 ) == ( bv_1_0_n53 )  ;
assign n29340 =  ( wr_addr ) == ( bv_8_255_n29279 )  ;
assign n29341 =  ( n29339 ) & (n29340 )  ;
assign n29342 =  ( n29341 ) & (wr )  ;
assign n29343 =  ( n29342 ) ? ( n5165 ) : ( iram_255 ) ;
assign n29344 = wr_addr[7:7] ;
assign n29345 =  ( n29344 ) == ( bv_1_0_n53 )  ;
assign n29346 =  ( wr_addr ) == ( bv_8_255_n29279 )  ;
assign n29347 =  ( n29345 ) & (n29346 )  ;
assign n29348 =  ( n29347 ) & (wr )  ;
assign n29349 =  ( n29348 ) ? ( n5204 ) : ( iram_255 ) ;
assign n29350 = wr_addr[7:7] ;
assign n29351 =  ( n29350 ) == ( bv_1_0_n53 )  ;
assign n29352 =  ( wr_addr ) == ( bv_8_255_n29279 )  ;
assign n29353 =  ( n29351 ) & (n29352 )  ;
assign n29354 =  ( n29353 ) & (wr )  ;
assign n29355 =  ( n29354 ) ? ( n5262 ) : ( iram_255 ) ;
assign n29356 = wr_addr[7:7] ;
assign n29357 =  ( n29356 ) == ( bv_1_0_n53 )  ;
assign n29358 =  ( wr_addr ) == ( bv_8_255_n29279 )  ;
assign n29359 =  ( n29357 ) & (n29358 )  ;
assign n29360 =  ( n29359 ) & (wr )  ;
assign n29361 =  ( n29360 ) ? ( n5298 ) : ( iram_255 ) ;
assign n29362 = wr_addr[7:7] ;
assign n29363 =  ( n29362 ) == ( bv_1_0_n53 )  ;
assign n29364 =  ( wr_addr ) == ( bv_8_255_n29279 )  ;
assign n29365 =  ( n29363 ) & (n29364 )  ;
assign n29366 =  ( n29365 ) & (wr )  ;
assign n29367 =  ( n29366 ) ? ( n5325 ) : ( iram_255 ) ;
always @(posedge clk) begin
   if(rst) begin
   end
   else if(__ILA_DATAPATH_valid__) begin
       if ( __ILA_DATAPATH_decode_of_read_data__ && __ILA_DATAPATH_grant__[15] ) begin
           bit_addr_r <= bit_addr;
       end else if ( __ILA_DATAPATH_decode_of_no_wr__ && __ILA_DATAPATH_grant__[16] ) begin
           bit_addr_r <= bit_addr;
       end else if ( __ILA_DATAPATH_decode_of_wr_sfr__ && __ILA_DATAPATH_grant__[17] ) begin
           bit_addr_r <= bit_addr;
       end else if ( __ILA_DATAPATH_decode_of_wr_ram__ && __ILA_DATAPATH_grant__[18] ) begin
           bit_addr_r <= bit_addr;
       end else if ( __ILA_DATAPATH_decode_of_wr_sfr_ram__ && __ILA_DATAPATH_grant__[19] ) begin
           bit_addr_r <= bit_addr;
       end
       if ( __ILA_DATAPATH_decode_of_read_data__ && __ILA_DATAPATH_grant__[15] ) begin
           bit_address <= n56;
       end else if ( __ILA_DATAPATH_decode_of_no_wr__ && __ILA_DATAPATH_grant__[16] ) begin
           bit_address <= n57;
       end else if ( __ILA_DATAPATH_decode_of_wr_sfr__ && __ILA_DATAPATH_grant__[17] ) begin
           bit_address <= n58;
       end else if ( __ILA_DATAPATH_decode_of_wr_ram__ && __ILA_DATAPATH_grant__[18] ) begin
           bit_address <= n59;
       end else if ( __ILA_DATAPATH_decode_of_wr_sfr_ram__ && __ILA_DATAPATH_grant__[19] ) begin
           bit_address <= n60;
       end
       if ( __ILA_DATAPATH_decode_of_read_data__ && __ILA_DATAPATH_grant__[15] ) begin
           ram_rd_data <= n1344;
       end else if ( __ILA_DATAPATH_decode_of_no_wr__ && __ILA_DATAPATH_grant__[16] ) begin
           ram_rd_data <= n1864;
       end else if ( __ILA_DATAPATH_decode_of_wr_sfr__ && __ILA_DATAPATH_grant__[17] ) begin
           ram_rd_data <= n2384;
       end else if ( __ILA_DATAPATH_decode_of_wr_ram__ && __ILA_DATAPATH_grant__[18] ) begin
           ram_rd_data <= n2915;
       end else if ( __ILA_DATAPATH_decode_of_wr_sfr_ram__ && __ILA_DATAPATH_grant__[19] ) begin
           ram_rd_data <= n3437;
       end
       if ( __ILA_DATAPATH_decode_of_read_data__ && __ILA_DATAPATH_grant__[15] ) begin
           sfr_rd_data <= n3494;
       end else if ( __ILA_DATAPATH_decode_of_no_wr__ && __ILA_DATAPATH_grant__[16] ) begin
           sfr_rd_data <= n3527;
       end else if ( __ILA_DATAPATH_decode_of_wr_sfr__ && __ILA_DATAPATH_grant__[17] ) begin
           sfr_rd_data <= n3573;
       end else if ( __ILA_DATAPATH_decode_of_wr_ram__ && __ILA_DATAPATH_grant__[18] ) begin
           sfr_rd_data <= n3599;
       end else if ( __ILA_DATAPATH_decode_of_wr_sfr_ram__ && __ILA_DATAPATH_grant__[19] ) begin
           sfr_rd_data <= n3644;
       end
       if ( __ILA_DATAPATH_decode_of_no_wr__ && __ILA_DATAPATH_grant__[16] ) begin
           sfr_bit_rd_data <= n3904;
       end else if ( __ILA_DATAPATH_decode_of_wr_sfr__ && __ILA_DATAPATH_grant__[17] ) begin
           sfr_bit_rd_data <= n4208;
       end else if ( __ILA_DATAPATH_decode_of_wr_ram__ && __ILA_DATAPATH_grant__[18] ) begin
           sfr_bit_rd_data <= n4452;
       end else if ( __ILA_DATAPATH_decode_of_wr_sfr_ram__ && __ILA_DATAPATH_grant__[19] ) begin
           sfr_bit_rd_data <= n4732;
       end
       if ( __ILA_DATAPATH_decode_of_read_data__ && __ILA_DATAPATH_grant__[15] ) begin
           rd_addr_r <= n4733;
       end else if ( __ILA_DATAPATH_decode_of_no_wr__ && __ILA_DATAPATH_grant__[16] ) begin
           rd_addr_r <= n4734;
       end else if ( __ILA_DATAPATH_decode_of_wr_sfr__ && __ILA_DATAPATH_grant__[17] ) begin
           rd_addr_r <= n4735;
       end else if ( __ILA_DATAPATH_decode_of_wr_ram__ && __ILA_DATAPATH_grant__[18] ) begin
           rd_addr_r <= n4736;
       end else if ( __ILA_DATAPATH_decode_of_wr_sfr_ram__ && __ILA_DATAPATH_grant__[19] ) begin
           rd_addr_r <= n4737;
       end
       if ( __ILA_DATAPATH_decode_of_read_data__ && __ILA_DATAPATH_grant__[15] ) begin
           wr_addr_r <= wr_addr;
       end
       if ( __ILA_DATAPATH_decode_of_read_data__ && __ILA_DATAPATH_grant__[15] ) begin
           rd_ind <= n4738;
       end else if ( __ILA_DATAPATH_decode_of_no_wr__ && __ILA_DATAPATH_grant__[16] ) begin
           rd_ind <= n4741;
       end else if ( __ILA_DATAPATH_decode_of_wr_sfr__ && __ILA_DATAPATH_grant__[17] ) begin
           rd_ind <= n4744;
       end else if ( __ILA_DATAPATH_decode_of_wr_ram__ && __ILA_DATAPATH_grant__[18] ) begin
           rd_ind <= n4747;
       end else if ( __ILA_DATAPATH_decode_of_wr_sfr_ram__ && __ILA_DATAPATH_grant__[19] ) begin
           rd_ind <= n4750;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           acc <= n4787;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           acc <= n4846;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           acc <= n4872;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           acc <= n4942;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           acc <= n4953;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           acc <= n4964;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           acc <= n5040;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           acc <= n5076;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           acc <= n5104;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           acc <= n5145;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           acc <= n5173;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           acc <= n5211;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           acc <= n5267;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           acc <= n5303;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           acc <= n5383;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           b_reg <= n5386;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           b_reg <= n5389;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           b_reg <= n5392;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           b_reg <= n5395;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           b_reg <= n5398;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           b_reg <= n5401;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           b_reg <= n5404;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           b_reg <= n5407;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           b_reg <= n5410;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           b_reg <= n5413;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           b_reg <= n5416;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           b_reg <= n5419;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           b_reg <= n5422;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           b_reg <= n5425;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           b_reg <= n5428;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           sp <= n5437;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           sp <= n5446;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           sp <= n5456;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           sp <= n5465;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           sp <= n5492;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           sp <= n5519;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           sp <= n5528;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           sp <= n5537;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           sp <= n5546;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           sp <= n5555;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           sp <= n5564;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           sp <= n5573;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           sp <= n5582;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           sp <= n5591;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           dptr_hi <= n5596;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           dptr_hi <= n5601;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           dptr_hi <= n5606;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           dptr_hi <= n5611;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           dptr_hi <= n5616;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           dptr_hi <= n5621;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           dptr_hi <= n5626;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           dptr_hi <= n5631;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           dptr_hi <= n5636;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           dptr_hi <= n5641;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           dptr_hi <= n5646;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           dptr_hi <= n5651;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           dptr_hi <= n5656;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           dptr_hi <= n5661;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           dptr_hi <= n5666;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           dptr_lo <= n5671;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           dptr_lo <= n5676;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           dptr_lo <= n5681;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           dptr_lo <= n5686;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           dptr_lo <= n5691;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           dptr_lo <= n5696;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           dptr_lo <= n5701;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           dptr_lo <= n5706;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           dptr_lo <= n5711;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           dptr_lo <= n5716;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           dptr_lo <= n5721;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           dptr_lo <= n5726;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           dptr_lo <= n5731;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           dptr_lo <= n5736;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           dptr_lo <= n5741;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           p0 <= n5744;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           p0 <= n5747;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           p0 <= n5750;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           p0 <= n5753;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           p0 <= n5756;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           p0 <= n5759;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           p0 <= n5762;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           p0 <= n5765;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           p0 <= n5768;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           p0 <= n5771;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           p0 <= n5774;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           p0 <= n5777;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           p0 <= n5780;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           p0 <= n5783;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           p0 <= n5786;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           p1 <= n5789;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           p1 <= n5792;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           p1 <= n5795;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           p1 <= n5798;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           p1 <= n5801;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           p1 <= n5804;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           p1 <= n5807;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           p1 <= n5810;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           p1 <= n5813;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           p1 <= n5816;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           p1 <= n5819;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           p1 <= n5822;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           p1 <= n5825;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           p1 <= n5828;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           p1 <= n5831;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           p2 <= n5834;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           p2 <= n5837;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           p2 <= n5840;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           p2 <= n5843;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           p2 <= n5846;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           p2 <= n5849;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           p2 <= n5852;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           p2 <= n5855;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           p2 <= n5858;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           p2 <= n5861;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           p2 <= n5864;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           p2 <= n5867;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           p2 <= n5870;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           p2 <= n5873;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           p2 <= n5876;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           p3 <= n5879;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           p3 <= n5882;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           p3 <= n5885;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           p3 <= n5888;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           p3 <= n5891;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           p3 <= n5894;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           p3 <= n5897;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           p3 <= n5900;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           p3 <= n5903;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           p3 <= n5906;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           p3 <= n5909;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           p3 <= n5912;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           p3 <= n5915;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           p3 <= n5918;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           p3 <= n5921;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           tcon <= n5924;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           tcon <= n5927;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           tcon <= n5930;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           tcon <= n5933;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           tcon <= n5936;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           tcon <= n5939;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           tcon <= n5942;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           tcon <= n5945;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           tcon <= n5948;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           tcon <= n5951;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           tcon <= n5954;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           tcon <= n5957;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           tcon <= n5960;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           tcon <= n5963;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           tcon <= n5966;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           scon <= n5969;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           scon <= n5972;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           scon <= n5975;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           scon <= n5978;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           scon <= n5981;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           scon <= n5984;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           scon <= n5987;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           scon <= n5990;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           scon <= n5993;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           scon <= n5996;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           scon <= n5999;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           scon <= n6002;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           scon <= n6005;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           scon <= n6008;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           scon <= n6011;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           pcon <= n6014;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           pcon <= n6017;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           pcon <= n6020;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           pcon <= n6023;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           pcon <= n6026;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           pcon <= n6029;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           pcon <= n6032;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           pcon <= n6035;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           pcon <= n6038;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           pcon <= n6041;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           pcon <= n6044;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           pcon <= n6047;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           pcon <= n6050;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           pcon <= n6053;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           pcon <= n6056;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           sbuf <= n6059;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           sbuf <= n6062;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           sbuf <= n6065;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           sbuf <= n6068;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           sbuf <= n6071;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           sbuf <= n6074;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           sbuf <= n6077;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           sbuf <= n6080;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           sbuf <= n6083;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           sbuf <= n6086;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           sbuf <= n6089;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           sbuf <= n6092;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           sbuf <= n6095;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           sbuf <= n6098;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           sbuf <= n6101;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           th0 <= n6104;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           th0 <= n6107;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           th0 <= n6110;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           th0 <= n6113;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           th0 <= n6116;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           th0 <= n6119;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           th0 <= n6122;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           th0 <= n6125;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           th0 <= n6128;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           th0 <= n6131;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           th0 <= n6134;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           th0 <= n6137;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           th0 <= n6140;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           th0 <= n6143;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           th0 <= n6146;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           th1 <= n6149;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           th1 <= n6152;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           th1 <= n6155;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           th1 <= n6158;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           th1 <= n6161;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           th1 <= n6164;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           th1 <= n6167;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           th1 <= n6170;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           th1 <= n6173;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           th1 <= n6176;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           th1 <= n6179;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           th1 <= n6182;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           th1 <= n6185;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           th1 <= n6188;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           th1 <= n6191;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           tl0 <= n6194;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           tl0 <= n6197;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           tl0 <= n6200;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           tl0 <= n6203;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           tl0 <= n6206;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           tl0 <= n6209;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           tl0 <= n6212;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           tl0 <= n6215;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           tl0 <= n6218;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           tl0 <= n6221;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           tl0 <= n6224;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           tl0 <= n6227;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           tl0 <= n6230;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           tl0 <= n6233;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           tl0 <= n6236;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           tl1 <= n6239;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           tl1 <= n6242;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           tl1 <= n6245;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           tl1 <= n6248;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           tl1 <= n6251;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           tl1 <= n6254;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           tl1 <= n6257;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           tl1 <= n6260;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           tl1 <= n6263;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           tl1 <= n6266;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           tl1 <= n6269;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           tl1 <= n6272;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           tl1 <= n6275;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           tl1 <= n6278;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           tl1 <= n6281;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           tmod <= n6284;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           tmod <= n6287;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           tmod <= n6290;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           tmod <= n6293;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           tmod <= n6296;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           tmod <= n6299;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           tmod <= n6302;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           tmod <= n6305;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           tmod <= n6308;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           tmod <= n6311;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           tmod <= n6314;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           tmod <= n6317;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           tmod <= n6320;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           tmod <= n6323;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           tmod <= n6326;
       end
       if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           op2_reg <= op2;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           op2_reg <= op2;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           op2_reg <= op2;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           op2_reg <= op2;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           op2_reg <= op2;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           op2_reg <= op2;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           op2_reg <= op2;
       end else if ( __ILA_DATAPATH_decode_of_read_data__ && __ILA_DATAPATH_grant__[15] ) begin
           op2_reg <= op2;
       end else if ( __ILA_DATAPATH_decode_of_no_wr__ && __ILA_DATAPATH_grant__[16] ) begin
           op2_reg <= op2;
       end else if ( __ILA_DATAPATH_decode_of_wr_sfr__ && __ILA_DATAPATH_grant__[17] ) begin
           op2_reg <= op2;
       end else if ( __ILA_DATAPATH_decode_of_wr_ram__ && __ILA_DATAPATH_grant__[18] ) begin
           op2_reg <= op2;
       end else if ( __ILA_DATAPATH_decode_of_wr_sfr_ram__ && __ILA_DATAPATH_grant__[19] ) begin
           op2_reg <= op2;
       end
       if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           op3_reg <= op3;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           op3_reg <= op3;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           op3_reg <= op3;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           op3_reg <= op3;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           op3_reg <= op3;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           op3_reg <= op3;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           op3_reg <= op3;
       end else if ( __ILA_DATAPATH_decode_of_read_data__ && __ILA_DATAPATH_grant__[15] ) begin
           op3_reg <= op3;
       end else if ( __ILA_DATAPATH_decode_of_no_wr__ && __ILA_DATAPATH_grant__[16] ) begin
           op3_reg <= op3;
       end else if ( __ILA_DATAPATH_decode_of_wr_sfr__ && __ILA_DATAPATH_grant__[17] ) begin
           op3_reg <= op3;
       end else if ( __ILA_DATAPATH_decode_of_wr_ram__ && __ILA_DATAPATH_grant__[18] ) begin
           op3_reg <= op3;
       end else if ( __ILA_DATAPATH_decode_of_wr_sfr_ram__ && __ILA_DATAPATH_grant__[19] ) begin
           op3_reg <= op3;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_0 <= n6332;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_0 <= n6338;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_0 <= n6344;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_0 <= n6350;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_0 <= n6356;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_0 <= n6362;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_0 <= n6368;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_0 <= n6374;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_0 <= n6380;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_0 <= n6386;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_0 <= n6392;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_0 <= n6398;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_0 <= n6404;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_0 <= n6410;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_0 <= n6416;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_1 <= n6422;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_1 <= n6428;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_1 <= n6434;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_1 <= n6440;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_1 <= n6446;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_1 <= n6452;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_1 <= n6458;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_1 <= n6464;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_1 <= n6470;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_1 <= n6476;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_1 <= n6482;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_1 <= n6488;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_1 <= n6494;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_1 <= n6500;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_1 <= n6506;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_2 <= n6512;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_2 <= n6518;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_2 <= n6524;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_2 <= n6530;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_2 <= n6536;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_2 <= n6542;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_2 <= n6548;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_2 <= n6554;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_2 <= n6560;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_2 <= n6566;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_2 <= n6572;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_2 <= n6578;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_2 <= n6584;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_2 <= n6590;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_2 <= n6596;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_3 <= n6602;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_3 <= n6608;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_3 <= n6614;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_3 <= n6620;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_3 <= n6626;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_3 <= n6632;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_3 <= n6638;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_3 <= n6644;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_3 <= n6650;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_3 <= n6656;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_3 <= n6662;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_3 <= n6668;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_3 <= n6674;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_3 <= n6680;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_3 <= n6686;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_4 <= n6692;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_4 <= n6698;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_4 <= n6704;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_4 <= n6710;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_4 <= n6716;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_4 <= n6722;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_4 <= n6728;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_4 <= n6734;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_4 <= n6740;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_4 <= n6746;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_4 <= n6752;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_4 <= n6758;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_4 <= n6764;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_4 <= n6770;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_4 <= n6776;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_5 <= n6782;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_5 <= n6788;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_5 <= n6794;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_5 <= n6800;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_5 <= n6806;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_5 <= n6812;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_5 <= n6818;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_5 <= n6824;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_5 <= n6830;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_5 <= n6836;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_5 <= n6842;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_5 <= n6848;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_5 <= n6854;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_5 <= n6860;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_5 <= n6866;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_6 <= n6872;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_6 <= n6878;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_6 <= n6884;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_6 <= n6890;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_6 <= n6896;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_6 <= n6902;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_6 <= n6908;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_6 <= n6914;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_6 <= n6920;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_6 <= n6926;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_6 <= n6932;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_6 <= n6938;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_6 <= n6944;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_6 <= n6950;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_6 <= n6956;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_7 <= n6962;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_7 <= n6968;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_7 <= n6974;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_7 <= n6980;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_7 <= n6986;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_7 <= n6992;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_7 <= n6998;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_7 <= n7004;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_7 <= n7010;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_7 <= n7016;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_7 <= n7022;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_7 <= n7028;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_7 <= n7034;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_7 <= n7040;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_7 <= n7046;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_8 <= n7052;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_8 <= n7058;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_8 <= n7064;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_8 <= n7070;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_8 <= n7076;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_8 <= n7082;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_8 <= n7088;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_8 <= n7094;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_8 <= n7100;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_8 <= n7106;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_8 <= n7112;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_8 <= n7118;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_8 <= n7124;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_8 <= n7130;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_8 <= n7136;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_9 <= n7142;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_9 <= n7148;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_9 <= n7154;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_9 <= n7160;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_9 <= n7166;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_9 <= n7172;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_9 <= n7178;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_9 <= n7184;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_9 <= n7190;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_9 <= n7196;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_9 <= n7202;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_9 <= n7208;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_9 <= n7214;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_9 <= n7220;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_9 <= n7226;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_10 <= n7232;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_10 <= n7238;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_10 <= n7244;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_10 <= n7250;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_10 <= n7256;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_10 <= n7262;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_10 <= n7268;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_10 <= n7274;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_10 <= n7280;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_10 <= n7286;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_10 <= n7292;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_10 <= n7298;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_10 <= n7304;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_10 <= n7310;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_10 <= n7316;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_11 <= n7322;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_11 <= n7328;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_11 <= n7334;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_11 <= n7340;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_11 <= n7346;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_11 <= n7352;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_11 <= n7358;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_11 <= n7364;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_11 <= n7370;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_11 <= n7376;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_11 <= n7382;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_11 <= n7388;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_11 <= n7394;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_11 <= n7400;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_11 <= n7406;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_12 <= n7412;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_12 <= n7418;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_12 <= n7424;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_12 <= n7430;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_12 <= n7436;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_12 <= n7442;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_12 <= n7448;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_12 <= n7454;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_12 <= n7460;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_12 <= n7466;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_12 <= n7472;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_12 <= n7478;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_12 <= n7484;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_12 <= n7490;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_12 <= n7496;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_13 <= n7502;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_13 <= n7508;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_13 <= n7514;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_13 <= n7520;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_13 <= n7526;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_13 <= n7532;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_13 <= n7538;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_13 <= n7544;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_13 <= n7550;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_13 <= n7556;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_13 <= n7562;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_13 <= n7568;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_13 <= n7574;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_13 <= n7580;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_13 <= n7586;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_14 <= n7592;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_14 <= n7598;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_14 <= n7604;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_14 <= n7610;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_14 <= n7616;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_14 <= n7622;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_14 <= n7628;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_14 <= n7634;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_14 <= n7640;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_14 <= n7646;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_14 <= n7652;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_14 <= n7658;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_14 <= n7664;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_14 <= n7670;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_14 <= n7676;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_15 <= n7682;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_15 <= n7688;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_15 <= n7694;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_15 <= n7700;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_15 <= n7706;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_15 <= n7712;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_15 <= n7718;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_15 <= n7724;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_15 <= n7730;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_15 <= n7736;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_15 <= n7742;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_15 <= n7748;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_15 <= n7754;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_15 <= n7760;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_15 <= n7766;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_16 <= n7772;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_16 <= n7778;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_16 <= n7784;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_16 <= n7790;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_16 <= n7796;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_16 <= n7802;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_16 <= n7808;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_16 <= n7814;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_16 <= n7820;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_16 <= n7826;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_16 <= n7832;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_16 <= n7838;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_16 <= n7844;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_16 <= n7850;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_16 <= n7856;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_17 <= n7862;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_17 <= n7868;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_17 <= n7874;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_17 <= n7880;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_17 <= n7886;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_17 <= n7892;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_17 <= n7898;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_17 <= n7904;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_17 <= n7910;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_17 <= n7916;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_17 <= n7922;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_17 <= n7928;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_17 <= n7934;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_17 <= n7940;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_17 <= n7946;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_18 <= n7952;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_18 <= n7958;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_18 <= n7964;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_18 <= n7970;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_18 <= n7976;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_18 <= n7982;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_18 <= n7988;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_18 <= n7994;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_18 <= n8000;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_18 <= n8006;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_18 <= n8012;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_18 <= n8018;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_18 <= n8024;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_18 <= n8030;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_18 <= n8036;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_19 <= n8042;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_19 <= n8048;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_19 <= n8054;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_19 <= n8060;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_19 <= n8066;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_19 <= n8072;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_19 <= n8078;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_19 <= n8084;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_19 <= n8090;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_19 <= n8096;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_19 <= n8102;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_19 <= n8108;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_19 <= n8114;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_19 <= n8120;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_19 <= n8126;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_20 <= n8132;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_20 <= n8138;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_20 <= n8144;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_20 <= n8150;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_20 <= n8156;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_20 <= n8162;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_20 <= n8168;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_20 <= n8174;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_20 <= n8180;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_20 <= n8186;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_20 <= n8192;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_20 <= n8198;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_20 <= n8204;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_20 <= n8210;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_20 <= n8216;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_21 <= n8222;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_21 <= n8228;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_21 <= n8234;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_21 <= n8240;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_21 <= n8246;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_21 <= n8252;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_21 <= n8258;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_21 <= n8264;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_21 <= n8270;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_21 <= n8276;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_21 <= n8282;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_21 <= n8288;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_21 <= n8294;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_21 <= n8300;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_21 <= n8306;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_22 <= n8312;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_22 <= n8318;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_22 <= n8324;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_22 <= n8330;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_22 <= n8336;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_22 <= n8342;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_22 <= n8348;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_22 <= n8354;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_22 <= n8360;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_22 <= n8366;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_22 <= n8372;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_22 <= n8378;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_22 <= n8384;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_22 <= n8390;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_22 <= n8396;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_23 <= n8402;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_23 <= n8408;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_23 <= n8414;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_23 <= n8420;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_23 <= n8426;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_23 <= n8432;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_23 <= n8438;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_23 <= n8444;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_23 <= n8450;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_23 <= n8456;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_23 <= n8462;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_23 <= n8468;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_23 <= n8474;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_23 <= n8480;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_23 <= n8486;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_24 <= n8492;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_24 <= n8498;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_24 <= n8504;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_24 <= n8510;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_24 <= n8516;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_24 <= n8522;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_24 <= n8528;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_24 <= n8534;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_24 <= n8540;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_24 <= n8546;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_24 <= n8552;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_24 <= n8558;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_24 <= n8564;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_24 <= n8570;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_24 <= n8576;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_25 <= n8582;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_25 <= n8588;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_25 <= n8594;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_25 <= n8600;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_25 <= n8606;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_25 <= n8612;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_25 <= n8618;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_25 <= n8624;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_25 <= n8630;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_25 <= n8636;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_25 <= n8642;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_25 <= n8648;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_25 <= n8654;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_25 <= n8660;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_25 <= n8666;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_26 <= n8672;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_26 <= n8678;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_26 <= n8684;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_26 <= n8690;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_26 <= n8696;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_26 <= n8702;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_26 <= n8708;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_26 <= n8714;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_26 <= n8720;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_26 <= n8726;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_26 <= n8732;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_26 <= n8738;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_26 <= n8744;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_26 <= n8750;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_26 <= n8756;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_27 <= n8762;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_27 <= n8768;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_27 <= n8774;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_27 <= n8780;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_27 <= n8786;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_27 <= n8792;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_27 <= n8798;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_27 <= n8804;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_27 <= n8810;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_27 <= n8816;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_27 <= n8822;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_27 <= n8828;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_27 <= n8834;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_27 <= n8840;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_27 <= n8846;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_28 <= n8852;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_28 <= n8858;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_28 <= n8864;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_28 <= n8870;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_28 <= n8876;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_28 <= n8882;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_28 <= n8888;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_28 <= n8894;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_28 <= n8900;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_28 <= n8906;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_28 <= n8912;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_28 <= n8918;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_28 <= n8924;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_28 <= n8930;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_28 <= n8936;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_29 <= n8942;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_29 <= n8948;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_29 <= n8954;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_29 <= n8960;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_29 <= n8966;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_29 <= n8972;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_29 <= n8978;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_29 <= n8984;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_29 <= n8990;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_29 <= n8996;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_29 <= n9002;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_29 <= n9008;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_29 <= n9014;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_29 <= n9020;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_29 <= n9026;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_30 <= n9032;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_30 <= n9038;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_30 <= n9044;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_30 <= n9050;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_30 <= n9056;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_30 <= n9062;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_30 <= n9068;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_30 <= n9074;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_30 <= n9080;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_30 <= n9086;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_30 <= n9092;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_30 <= n9098;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_30 <= n9104;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_30 <= n9110;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_30 <= n9116;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_31 <= n9122;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_31 <= n9128;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_31 <= n9134;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_31 <= n9140;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_31 <= n9146;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_31 <= n9152;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_31 <= n9158;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_31 <= n9164;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_31 <= n9170;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_31 <= n9176;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_31 <= n9182;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_31 <= n9188;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_31 <= n9194;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_31 <= n9200;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_31 <= n9206;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_32 <= n9212;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_32 <= n9218;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_32 <= n9224;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_32 <= n9230;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_32 <= n9236;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_32 <= n9242;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_32 <= n9248;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_32 <= n9254;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_32 <= n9260;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_32 <= n9266;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_32 <= n9272;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_32 <= n9278;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_32 <= n9284;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_32 <= n9290;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_32 <= n9296;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_33 <= n9302;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_33 <= n9308;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_33 <= n9314;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_33 <= n9320;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_33 <= n9326;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_33 <= n9332;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_33 <= n9338;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_33 <= n9344;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_33 <= n9350;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_33 <= n9356;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_33 <= n9362;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_33 <= n9368;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_33 <= n9374;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_33 <= n9380;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_33 <= n9386;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_34 <= n9392;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_34 <= n9398;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_34 <= n9404;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_34 <= n9410;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_34 <= n9416;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_34 <= n9422;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_34 <= n9428;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_34 <= n9434;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_34 <= n9440;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_34 <= n9446;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_34 <= n9452;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_34 <= n9458;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_34 <= n9464;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_34 <= n9470;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_34 <= n9476;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_35 <= n9482;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_35 <= n9488;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_35 <= n9494;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_35 <= n9500;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_35 <= n9506;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_35 <= n9512;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_35 <= n9518;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_35 <= n9524;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_35 <= n9530;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_35 <= n9536;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_35 <= n9542;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_35 <= n9548;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_35 <= n9554;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_35 <= n9560;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_35 <= n9566;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_36 <= n9572;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_36 <= n9578;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_36 <= n9584;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_36 <= n9590;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_36 <= n9596;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_36 <= n9602;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_36 <= n9608;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_36 <= n9614;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_36 <= n9620;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_36 <= n9626;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_36 <= n9632;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_36 <= n9638;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_36 <= n9644;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_36 <= n9650;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_36 <= n9656;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_37 <= n9662;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_37 <= n9668;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_37 <= n9674;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_37 <= n9680;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_37 <= n9686;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_37 <= n9692;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_37 <= n9698;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_37 <= n9704;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_37 <= n9710;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_37 <= n9716;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_37 <= n9722;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_37 <= n9728;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_37 <= n9734;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_37 <= n9740;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_37 <= n9746;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_38 <= n9752;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_38 <= n9758;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_38 <= n9764;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_38 <= n9770;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_38 <= n9776;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_38 <= n9782;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_38 <= n9788;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_38 <= n9794;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_38 <= n9800;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_38 <= n9806;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_38 <= n9812;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_38 <= n9818;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_38 <= n9824;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_38 <= n9830;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_38 <= n9836;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_39 <= n9842;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_39 <= n9848;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_39 <= n9854;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_39 <= n9860;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_39 <= n9866;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_39 <= n9872;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_39 <= n9878;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_39 <= n9884;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_39 <= n9890;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_39 <= n9896;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_39 <= n9902;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_39 <= n9908;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_39 <= n9914;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_39 <= n9920;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_39 <= n9926;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_40 <= n9932;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_40 <= n9938;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_40 <= n9944;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_40 <= n9950;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_40 <= n9956;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_40 <= n9962;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_40 <= n9968;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_40 <= n9974;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_40 <= n9980;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_40 <= n9986;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_40 <= n9992;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_40 <= n9998;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_40 <= n10004;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_40 <= n10010;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_40 <= n10016;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_41 <= n10022;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_41 <= n10028;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_41 <= n10034;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_41 <= n10040;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_41 <= n10046;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_41 <= n10052;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_41 <= n10058;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_41 <= n10064;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_41 <= n10070;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_41 <= n10076;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_41 <= n10082;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_41 <= n10088;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_41 <= n10094;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_41 <= n10100;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_41 <= n10106;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_42 <= n10112;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_42 <= n10118;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_42 <= n10124;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_42 <= n10130;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_42 <= n10136;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_42 <= n10142;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_42 <= n10148;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_42 <= n10154;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_42 <= n10160;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_42 <= n10166;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_42 <= n10172;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_42 <= n10178;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_42 <= n10184;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_42 <= n10190;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_42 <= n10196;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_43 <= n10202;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_43 <= n10208;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_43 <= n10214;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_43 <= n10220;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_43 <= n10226;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_43 <= n10232;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_43 <= n10238;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_43 <= n10244;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_43 <= n10250;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_43 <= n10256;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_43 <= n10262;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_43 <= n10268;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_43 <= n10274;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_43 <= n10280;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_43 <= n10286;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_44 <= n10292;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_44 <= n10298;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_44 <= n10304;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_44 <= n10310;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_44 <= n10316;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_44 <= n10322;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_44 <= n10328;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_44 <= n10334;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_44 <= n10340;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_44 <= n10346;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_44 <= n10352;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_44 <= n10358;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_44 <= n10364;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_44 <= n10370;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_44 <= n10376;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_45 <= n10382;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_45 <= n10388;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_45 <= n10394;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_45 <= n10400;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_45 <= n10406;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_45 <= n10412;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_45 <= n10418;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_45 <= n10424;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_45 <= n10430;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_45 <= n10436;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_45 <= n10442;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_45 <= n10448;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_45 <= n10454;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_45 <= n10460;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_45 <= n10466;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_46 <= n10472;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_46 <= n10478;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_46 <= n10484;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_46 <= n10490;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_46 <= n10496;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_46 <= n10502;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_46 <= n10508;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_46 <= n10514;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_46 <= n10520;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_46 <= n10526;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_46 <= n10532;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_46 <= n10538;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_46 <= n10544;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_46 <= n10550;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_46 <= n10556;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_47 <= n10562;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_47 <= n10568;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_47 <= n10574;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_47 <= n10580;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_47 <= n10586;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_47 <= n10592;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_47 <= n10598;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_47 <= n10604;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_47 <= n10610;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_47 <= n10616;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_47 <= n10622;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_47 <= n10628;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_47 <= n10634;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_47 <= n10640;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_47 <= n10646;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_48 <= n10652;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_48 <= n10658;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_48 <= n10664;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_48 <= n10670;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_48 <= n10676;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_48 <= n10682;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_48 <= n10688;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_48 <= n10694;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_48 <= n10700;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_48 <= n10706;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_48 <= n10712;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_48 <= n10718;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_48 <= n10724;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_48 <= n10730;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_48 <= n10736;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_49 <= n10742;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_49 <= n10748;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_49 <= n10754;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_49 <= n10760;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_49 <= n10766;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_49 <= n10772;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_49 <= n10778;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_49 <= n10784;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_49 <= n10790;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_49 <= n10796;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_49 <= n10802;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_49 <= n10808;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_49 <= n10814;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_49 <= n10820;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_49 <= n10826;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_50 <= n10832;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_50 <= n10838;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_50 <= n10844;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_50 <= n10850;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_50 <= n10856;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_50 <= n10862;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_50 <= n10868;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_50 <= n10874;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_50 <= n10880;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_50 <= n10886;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_50 <= n10892;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_50 <= n10898;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_50 <= n10904;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_50 <= n10910;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_50 <= n10916;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_51 <= n10922;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_51 <= n10928;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_51 <= n10934;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_51 <= n10940;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_51 <= n10946;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_51 <= n10952;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_51 <= n10958;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_51 <= n10964;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_51 <= n10970;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_51 <= n10976;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_51 <= n10982;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_51 <= n10988;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_51 <= n10994;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_51 <= n11000;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_51 <= n11006;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_52 <= n11012;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_52 <= n11018;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_52 <= n11024;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_52 <= n11030;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_52 <= n11036;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_52 <= n11042;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_52 <= n11048;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_52 <= n11054;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_52 <= n11060;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_52 <= n11066;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_52 <= n11072;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_52 <= n11078;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_52 <= n11084;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_52 <= n11090;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_52 <= n11096;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_53 <= n11102;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_53 <= n11108;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_53 <= n11114;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_53 <= n11120;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_53 <= n11126;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_53 <= n11132;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_53 <= n11138;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_53 <= n11144;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_53 <= n11150;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_53 <= n11156;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_53 <= n11162;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_53 <= n11168;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_53 <= n11174;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_53 <= n11180;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_53 <= n11186;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_54 <= n11192;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_54 <= n11198;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_54 <= n11204;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_54 <= n11210;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_54 <= n11216;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_54 <= n11222;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_54 <= n11228;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_54 <= n11234;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_54 <= n11240;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_54 <= n11246;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_54 <= n11252;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_54 <= n11258;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_54 <= n11264;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_54 <= n11270;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_54 <= n11276;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_55 <= n11282;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_55 <= n11288;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_55 <= n11294;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_55 <= n11300;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_55 <= n11306;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_55 <= n11312;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_55 <= n11318;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_55 <= n11324;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_55 <= n11330;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_55 <= n11336;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_55 <= n11342;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_55 <= n11348;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_55 <= n11354;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_55 <= n11360;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_55 <= n11366;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_56 <= n11372;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_56 <= n11378;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_56 <= n11384;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_56 <= n11390;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_56 <= n11396;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_56 <= n11402;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_56 <= n11408;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_56 <= n11414;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_56 <= n11420;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_56 <= n11426;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_56 <= n11432;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_56 <= n11438;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_56 <= n11444;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_56 <= n11450;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_56 <= n11456;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_57 <= n11462;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_57 <= n11468;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_57 <= n11474;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_57 <= n11480;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_57 <= n11486;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_57 <= n11492;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_57 <= n11498;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_57 <= n11504;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_57 <= n11510;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_57 <= n11516;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_57 <= n11522;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_57 <= n11528;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_57 <= n11534;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_57 <= n11540;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_57 <= n11546;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_58 <= n11552;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_58 <= n11558;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_58 <= n11564;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_58 <= n11570;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_58 <= n11576;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_58 <= n11582;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_58 <= n11588;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_58 <= n11594;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_58 <= n11600;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_58 <= n11606;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_58 <= n11612;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_58 <= n11618;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_58 <= n11624;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_58 <= n11630;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_58 <= n11636;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_59 <= n11642;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_59 <= n11648;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_59 <= n11654;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_59 <= n11660;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_59 <= n11666;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_59 <= n11672;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_59 <= n11678;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_59 <= n11684;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_59 <= n11690;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_59 <= n11696;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_59 <= n11702;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_59 <= n11708;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_59 <= n11714;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_59 <= n11720;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_59 <= n11726;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_60 <= n11732;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_60 <= n11738;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_60 <= n11744;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_60 <= n11750;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_60 <= n11756;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_60 <= n11762;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_60 <= n11768;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_60 <= n11774;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_60 <= n11780;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_60 <= n11786;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_60 <= n11792;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_60 <= n11798;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_60 <= n11804;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_60 <= n11810;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_60 <= n11816;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_61 <= n11822;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_61 <= n11828;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_61 <= n11834;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_61 <= n11840;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_61 <= n11846;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_61 <= n11852;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_61 <= n11858;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_61 <= n11864;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_61 <= n11870;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_61 <= n11876;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_61 <= n11882;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_61 <= n11888;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_61 <= n11894;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_61 <= n11900;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_61 <= n11906;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_62 <= n11912;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_62 <= n11918;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_62 <= n11924;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_62 <= n11930;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_62 <= n11936;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_62 <= n11942;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_62 <= n11948;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_62 <= n11954;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_62 <= n11960;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_62 <= n11966;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_62 <= n11972;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_62 <= n11978;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_62 <= n11984;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_62 <= n11990;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_62 <= n11996;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_63 <= n12002;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_63 <= n12008;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_63 <= n12014;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_63 <= n12020;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_63 <= n12026;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_63 <= n12032;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_63 <= n12038;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_63 <= n12044;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_63 <= n12050;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_63 <= n12056;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_63 <= n12062;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_63 <= n12068;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_63 <= n12074;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_63 <= n12080;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_63 <= n12086;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_64 <= n12092;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_64 <= n12098;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_64 <= n12104;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_64 <= n12110;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_64 <= n12116;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_64 <= n12122;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_64 <= n12128;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_64 <= n12134;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_64 <= n12140;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_64 <= n12146;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_64 <= n12152;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_64 <= n12158;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_64 <= n12164;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_64 <= n12170;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_64 <= n12176;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_65 <= n12182;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_65 <= n12188;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_65 <= n12194;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_65 <= n12200;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_65 <= n12206;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_65 <= n12212;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_65 <= n12218;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_65 <= n12224;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_65 <= n12230;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_65 <= n12236;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_65 <= n12242;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_65 <= n12248;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_65 <= n12254;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_65 <= n12260;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_65 <= n12266;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_66 <= n12272;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_66 <= n12278;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_66 <= n12284;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_66 <= n12290;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_66 <= n12296;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_66 <= n12302;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_66 <= n12308;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_66 <= n12314;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_66 <= n12320;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_66 <= n12326;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_66 <= n12332;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_66 <= n12338;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_66 <= n12344;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_66 <= n12350;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_66 <= n12356;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_67 <= n12362;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_67 <= n12368;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_67 <= n12374;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_67 <= n12380;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_67 <= n12386;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_67 <= n12392;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_67 <= n12398;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_67 <= n12404;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_67 <= n12410;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_67 <= n12416;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_67 <= n12422;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_67 <= n12428;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_67 <= n12434;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_67 <= n12440;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_67 <= n12446;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_68 <= n12452;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_68 <= n12458;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_68 <= n12464;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_68 <= n12470;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_68 <= n12476;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_68 <= n12482;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_68 <= n12488;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_68 <= n12494;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_68 <= n12500;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_68 <= n12506;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_68 <= n12512;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_68 <= n12518;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_68 <= n12524;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_68 <= n12530;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_68 <= n12536;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_69 <= n12542;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_69 <= n12548;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_69 <= n12554;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_69 <= n12560;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_69 <= n12566;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_69 <= n12572;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_69 <= n12578;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_69 <= n12584;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_69 <= n12590;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_69 <= n12596;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_69 <= n12602;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_69 <= n12608;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_69 <= n12614;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_69 <= n12620;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_69 <= n12626;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_70 <= n12632;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_70 <= n12638;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_70 <= n12644;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_70 <= n12650;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_70 <= n12656;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_70 <= n12662;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_70 <= n12668;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_70 <= n12674;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_70 <= n12680;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_70 <= n12686;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_70 <= n12692;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_70 <= n12698;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_70 <= n12704;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_70 <= n12710;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_70 <= n12716;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_71 <= n12722;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_71 <= n12728;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_71 <= n12734;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_71 <= n12740;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_71 <= n12746;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_71 <= n12752;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_71 <= n12758;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_71 <= n12764;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_71 <= n12770;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_71 <= n12776;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_71 <= n12782;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_71 <= n12788;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_71 <= n12794;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_71 <= n12800;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_71 <= n12806;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_72 <= n12812;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_72 <= n12818;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_72 <= n12824;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_72 <= n12830;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_72 <= n12836;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_72 <= n12842;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_72 <= n12848;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_72 <= n12854;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_72 <= n12860;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_72 <= n12866;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_72 <= n12872;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_72 <= n12878;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_72 <= n12884;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_72 <= n12890;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_72 <= n12896;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_73 <= n12902;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_73 <= n12908;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_73 <= n12914;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_73 <= n12920;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_73 <= n12926;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_73 <= n12932;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_73 <= n12938;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_73 <= n12944;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_73 <= n12950;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_73 <= n12956;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_73 <= n12962;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_73 <= n12968;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_73 <= n12974;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_73 <= n12980;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_73 <= n12986;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_74 <= n12992;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_74 <= n12998;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_74 <= n13004;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_74 <= n13010;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_74 <= n13016;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_74 <= n13022;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_74 <= n13028;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_74 <= n13034;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_74 <= n13040;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_74 <= n13046;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_74 <= n13052;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_74 <= n13058;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_74 <= n13064;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_74 <= n13070;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_74 <= n13076;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_75 <= n13082;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_75 <= n13088;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_75 <= n13094;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_75 <= n13100;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_75 <= n13106;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_75 <= n13112;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_75 <= n13118;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_75 <= n13124;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_75 <= n13130;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_75 <= n13136;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_75 <= n13142;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_75 <= n13148;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_75 <= n13154;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_75 <= n13160;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_75 <= n13166;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_76 <= n13172;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_76 <= n13178;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_76 <= n13184;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_76 <= n13190;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_76 <= n13196;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_76 <= n13202;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_76 <= n13208;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_76 <= n13214;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_76 <= n13220;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_76 <= n13226;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_76 <= n13232;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_76 <= n13238;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_76 <= n13244;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_76 <= n13250;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_76 <= n13256;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_77 <= n13262;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_77 <= n13268;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_77 <= n13274;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_77 <= n13280;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_77 <= n13286;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_77 <= n13292;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_77 <= n13298;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_77 <= n13304;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_77 <= n13310;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_77 <= n13316;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_77 <= n13322;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_77 <= n13328;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_77 <= n13334;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_77 <= n13340;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_77 <= n13346;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_78 <= n13352;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_78 <= n13358;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_78 <= n13364;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_78 <= n13370;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_78 <= n13376;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_78 <= n13382;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_78 <= n13388;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_78 <= n13394;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_78 <= n13400;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_78 <= n13406;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_78 <= n13412;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_78 <= n13418;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_78 <= n13424;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_78 <= n13430;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_78 <= n13436;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_79 <= n13442;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_79 <= n13448;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_79 <= n13454;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_79 <= n13460;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_79 <= n13466;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_79 <= n13472;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_79 <= n13478;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_79 <= n13484;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_79 <= n13490;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_79 <= n13496;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_79 <= n13502;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_79 <= n13508;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_79 <= n13514;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_79 <= n13520;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_79 <= n13526;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_80 <= n13532;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_80 <= n13538;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_80 <= n13544;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_80 <= n13550;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_80 <= n13556;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_80 <= n13562;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_80 <= n13568;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_80 <= n13574;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_80 <= n13580;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_80 <= n13586;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_80 <= n13592;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_80 <= n13598;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_80 <= n13604;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_80 <= n13610;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_80 <= n13616;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_81 <= n13622;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_81 <= n13628;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_81 <= n13634;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_81 <= n13640;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_81 <= n13646;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_81 <= n13652;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_81 <= n13658;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_81 <= n13664;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_81 <= n13670;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_81 <= n13676;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_81 <= n13682;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_81 <= n13688;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_81 <= n13694;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_81 <= n13700;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_81 <= n13706;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_82 <= n13712;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_82 <= n13718;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_82 <= n13724;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_82 <= n13730;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_82 <= n13736;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_82 <= n13742;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_82 <= n13748;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_82 <= n13754;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_82 <= n13760;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_82 <= n13766;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_82 <= n13772;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_82 <= n13778;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_82 <= n13784;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_82 <= n13790;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_82 <= n13796;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_83 <= n13802;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_83 <= n13808;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_83 <= n13814;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_83 <= n13820;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_83 <= n13826;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_83 <= n13832;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_83 <= n13838;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_83 <= n13844;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_83 <= n13850;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_83 <= n13856;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_83 <= n13862;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_83 <= n13868;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_83 <= n13874;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_83 <= n13880;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_83 <= n13886;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_84 <= n13892;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_84 <= n13898;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_84 <= n13904;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_84 <= n13910;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_84 <= n13916;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_84 <= n13922;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_84 <= n13928;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_84 <= n13934;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_84 <= n13940;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_84 <= n13946;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_84 <= n13952;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_84 <= n13958;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_84 <= n13964;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_84 <= n13970;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_84 <= n13976;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_85 <= n13982;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_85 <= n13988;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_85 <= n13994;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_85 <= n14000;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_85 <= n14006;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_85 <= n14012;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_85 <= n14018;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_85 <= n14024;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_85 <= n14030;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_85 <= n14036;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_85 <= n14042;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_85 <= n14048;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_85 <= n14054;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_85 <= n14060;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_85 <= n14066;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_86 <= n14072;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_86 <= n14078;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_86 <= n14084;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_86 <= n14090;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_86 <= n14096;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_86 <= n14102;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_86 <= n14108;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_86 <= n14114;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_86 <= n14120;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_86 <= n14126;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_86 <= n14132;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_86 <= n14138;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_86 <= n14144;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_86 <= n14150;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_86 <= n14156;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_87 <= n14162;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_87 <= n14168;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_87 <= n14174;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_87 <= n14180;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_87 <= n14186;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_87 <= n14192;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_87 <= n14198;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_87 <= n14204;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_87 <= n14210;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_87 <= n14216;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_87 <= n14222;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_87 <= n14228;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_87 <= n14234;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_87 <= n14240;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_87 <= n14246;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_88 <= n14252;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_88 <= n14258;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_88 <= n14264;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_88 <= n14270;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_88 <= n14276;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_88 <= n14282;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_88 <= n14288;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_88 <= n14294;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_88 <= n14300;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_88 <= n14306;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_88 <= n14312;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_88 <= n14318;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_88 <= n14324;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_88 <= n14330;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_88 <= n14336;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_89 <= n14342;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_89 <= n14348;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_89 <= n14354;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_89 <= n14360;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_89 <= n14366;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_89 <= n14372;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_89 <= n14378;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_89 <= n14384;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_89 <= n14390;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_89 <= n14396;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_89 <= n14402;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_89 <= n14408;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_89 <= n14414;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_89 <= n14420;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_89 <= n14426;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_90 <= n14432;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_90 <= n14438;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_90 <= n14444;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_90 <= n14450;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_90 <= n14456;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_90 <= n14462;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_90 <= n14468;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_90 <= n14474;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_90 <= n14480;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_90 <= n14486;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_90 <= n14492;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_90 <= n14498;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_90 <= n14504;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_90 <= n14510;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_90 <= n14516;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_91 <= n14522;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_91 <= n14528;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_91 <= n14534;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_91 <= n14540;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_91 <= n14546;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_91 <= n14552;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_91 <= n14558;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_91 <= n14564;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_91 <= n14570;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_91 <= n14576;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_91 <= n14582;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_91 <= n14588;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_91 <= n14594;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_91 <= n14600;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_91 <= n14606;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_92 <= n14612;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_92 <= n14618;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_92 <= n14624;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_92 <= n14630;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_92 <= n14636;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_92 <= n14642;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_92 <= n14648;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_92 <= n14654;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_92 <= n14660;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_92 <= n14666;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_92 <= n14672;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_92 <= n14678;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_92 <= n14684;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_92 <= n14690;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_92 <= n14696;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_93 <= n14702;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_93 <= n14708;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_93 <= n14714;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_93 <= n14720;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_93 <= n14726;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_93 <= n14732;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_93 <= n14738;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_93 <= n14744;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_93 <= n14750;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_93 <= n14756;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_93 <= n14762;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_93 <= n14768;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_93 <= n14774;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_93 <= n14780;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_93 <= n14786;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_94 <= n14792;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_94 <= n14798;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_94 <= n14804;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_94 <= n14810;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_94 <= n14816;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_94 <= n14822;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_94 <= n14828;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_94 <= n14834;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_94 <= n14840;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_94 <= n14846;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_94 <= n14852;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_94 <= n14858;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_94 <= n14864;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_94 <= n14870;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_94 <= n14876;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_95 <= n14882;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_95 <= n14888;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_95 <= n14894;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_95 <= n14900;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_95 <= n14906;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_95 <= n14912;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_95 <= n14918;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_95 <= n14924;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_95 <= n14930;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_95 <= n14936;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_95 <= n14942;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_95 <= n14948;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_95 <= n14954;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_95 <= n14960;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_95 <= n14966;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_96 <= n14972;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_96 <= n14978;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_96 <= n14984;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_96 <= n14990;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_96 <= n14996;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_96 <= n15002;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_96 <= n15008;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_96 <= n15014;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_96 <= n15020;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_96 <= n15026;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_96 <= n15032;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_96 <= n15038;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_96 <= n15044;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_96 <= n15050;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_96 <= n15056;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_97 <= n15062;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_97 <= n15068;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_97 <= n15074;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_97 <= n15080;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_97 <= n15086;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_97 <= n15092;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_97 <= n15098;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_97 <= n15104;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_97 <= n15110;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_97 <= n15116;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_97 <= n15122;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_97 <= n15128;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_97 <= n15134;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_97 <= n15140;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_97 <= n15146;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_98 <= n15152;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_98 <= n15158;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_98 <= n15164;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_98 <= n15170;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_98 <= n15176;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_98 <= n15182;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_98 <= n15188;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_98 <= n15194;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_98 <= n15200;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_98 <= n15206;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_98 <= n15212;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_98 <= n15218;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_98 <= n15224;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_98 <= n15230;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_98 <= n15236;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_99 <= n15242;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_99 <= n15248;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_99 <= n15254;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_99 <= n15260;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_99 <= n15266;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_99 <= n15272;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_99 <= n15278;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_99 <= n15284;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_99 <= n15290;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_99 <= n15296;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_99 <= n15302;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_99 <= n15308;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_99 <= n15314;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_99 <= n15320;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_99 <= n15326;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_100 <= n15332;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_100 <= n15338;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_100 <= n15344;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_100 <= n15350;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_100 <= n15356;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_100 <= n15362;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_100 <= n15368;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_100 <= n15374;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_100 <= n15380;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_100 <= n15386;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_100 <= n15392;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_100 <= n15398;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_100 <= n15404;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_100 <= n15410;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_100 <= n15416;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_101 <= n15422;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_101 <= n15428;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_101 <= n15434;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_101 <= n15440;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_101 <= n15446;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_101 <= n15452;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_101 <= n15458;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_101 <= n15464;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_101 <= n15470;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_101 <= n15476;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_101 <= n15482;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_101 <= n15488;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_101 <= n15494;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_101 <= n15500;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_101 <= n15506;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_102 <= n15512;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_102 <= n15518;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_102 <= n15524;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_102 <= n15530;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_102 <= n15536;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_102 <= n15542;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_102 <= n15548;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_102 <= n15554;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_102 <= n15560;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_102 <= n15566;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_102 <= n15572;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_102 <= n15578;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_102 <= n15584;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_102 <= n15590;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_102 <= n15596;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_103 <= n15602;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_103 <= n15608;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_103 <= n15614;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_103 <= n15620;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_103 <= n15626;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_103 <= n15632;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_103 <= n15638;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_103 <= n15644;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_103 <= n15650;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_103 <= n15656;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_103 <= n15662;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_103 <= n15668;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_103 <= n15674;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_103 <= n15680;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_103 <= n15686;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_104 <= n15692;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_104 <= n15698;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_104 <= n15704;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_104 <= n15710;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_104 <= n15716;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_104 <= n15722;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_104 <= n15728;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_104 <= n15734;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_104 <= n15740;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_104 <= n15746;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_104 <= n15752;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_104 <= n15758;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_104 <= n15764;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_104 <= n15770;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_104 <= n15776;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_105 <= n15782;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_105 <= n15788;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_105 <= n15794;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_105 <= n15800;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_105 <= n15806;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_105 <= n15812;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_105 <= n15818;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_105 <= n15824;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_105 <= n15830;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_105 <= n15836;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_105 <= n15842;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_105 <= n15848;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_105 <= n15854;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_105 <= n15860;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_105 <= n15866;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_106 <= n15872;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_106 <= n15878;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_106 <= n15884;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_106 <= n15890;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_106 <= n15896;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_106 <= n15902;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_106 <= n15908;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_106 <= n15914;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_106 <= n15920;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_106 <= n15926;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_106 <= n15932;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_106 <= n15938;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_106 <= n15944;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_106 <= n15950;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_106 <= n15956;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_107 <= n15962;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_107 <= n15968;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_107 <= n15974;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_107 <= n15980;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_107 <= n15986;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_107 <= n15992;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_107 <= n15998;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_107 <= n16004;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_107 <= n16010;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_107 <= n16016;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_107 <= n16022;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_107 <= n16028;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_107 <= n16034;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_107 <= n16040;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_107 <= n16046;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_108 <= n16052;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_108 <= n16058;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_108 <= n16064;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_108 <= n16070;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_108 <= n16076;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_108 <= n16082;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_108 <= n16088;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_108 <= n16094;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_108 <= n16100;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_108 <= n16106;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_108 <= n16112;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_108 <= n16118;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_108 <= n16124;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_108 <= n16130;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_108 <= n16136;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_109 <= n16142;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_109 <= n16148;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_109 <= n16154;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_109 <= n16160;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_109 <= n16166;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_109 <= n16172;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_109 <= n16178;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_109 <= n16184;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_109 <= n16190;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_109 <= n16196;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_109 <= n16202;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_109 <= n16208;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_109 <= n16214;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_109 <= n16220;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_109 <= n16226;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_110 <= n16232;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_110 <= n16238;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_110 <= n16244;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_110 <= n16250;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_110 <= n16256;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_110 <= n16262;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_110 <= n16268;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_110 <= n16274;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_110 <= n16280;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_110 <= n16286;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_110 <= n16292;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_110 <= n16298;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_110 <= n16304;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_110 <= n16310;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_110 <= n16316;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_111 <= n16322;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_111 <= n16328;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_111 <= n16334;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_111 <= n16340;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_111 <= n16346;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_111 <= n16352;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_111 <= n16358;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_111 <= n16364;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_111 <= n16370;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_111 <= n16376;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_111 <= n16382;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_111 <= n16388;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_111 <= n16394;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_111 <= n16400;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_111 <= n16406;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_112 <= n16412;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_112 <= n16418;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_112 <= n16424;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_112 <= n16430;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_112 <= n16436;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_112 <= n16442;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_112 <= n16448;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_112 <= n16454;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_112 <= n16460;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_112 <= n16466;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_112 <= n16472;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_112 <= n16478;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_112 <= n16484;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_112 <= n16490;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_112 <= n16496;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_113 <= n16502;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_113 <= n16508;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_113 <= n16514;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_113 <= n16520;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_113 <= n16526;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_113 <= n16532;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_113 <= n16538;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_113 <= n16544;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_113 <= n16550;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_113 <= n16556;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_113 <= n16562;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_113 <= n16568;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_113 <= n16574;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_113 <= n16580;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_113 <= n16586;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_114 <= n16592;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_114 <= n16598;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_114 <= n16604;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_114 <= n16610;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_114 <= n16616;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_114 <= n16622;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_114 <= n16628;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_114 <= n16634;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_114 <= n16640;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_114 <= n16646;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_114 <= n16652;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_114 <= n16658;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_114 <= n16664;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_114 <= n16670;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_114 <= n16676;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_115 <= n16682;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_115 <= n16688;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_115 <= n16694;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_115 <= n16700;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_115 <= n16706;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_115 <= n16712;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_115 <= n16718;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_115 <= n16724;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_115 <= n16730;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_115 <= n16736;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_115 <= n16742;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_115 <= n16748;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_115 <= n16754;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_115 <= n16760;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_115 <= n16766;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_116 <= n16772;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_116 <= n16778;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_116 <= n16784;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_116 <= n16790;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_116 <= n16796;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_116 <= n16802;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_116 <= n16808;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_116 <= n16814;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_116 <= n16820;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_116 <= n16826;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_116 <= n16832;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_116 <= n16838;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_116 <= n16844;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_116 <= n16850;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_116 <= n16856;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_117 <= n16862;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_117 <= n16868;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_117 <= n16874;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_117 <= n16880;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_117 <= n16886;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_117 <= n16892;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_117 <= n16898;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_117 <= n16904;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_117 <= n16910;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_117 <= n16916;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_117 <= n16922;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_117 <= n16928;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_117 <= n16934;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_117 <= n16940;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_117 <= n16946;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_118 <= n16952;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_118 <= n16958;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_118 <= n16964;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_118 <= n16970;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_118 <= n16976;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_118 <= n16982;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_118 <= n16988;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_118 <= n16994;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_118 <= n17000;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_118 <= n17006;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_118 <= n17012;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_118 <= n17018;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_118 <= n17024;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_118 <= n17030;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_118 <= n17036;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_119 <= n17042;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_119 <= n17048;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_119 <= n17054;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_119 <= n17060;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_119 <= n17066;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_119 <= n17072;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_119 <= n17078;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_119 <= n17084;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_119 <= n17090;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_119 <= n17096;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_119 <= n17102;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_119 <= n17108;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_119 <= n17114;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_119 <= n17120;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_119 <= n17126;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_120 <= n17132;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_120 <= n17138;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_120 <= n17144;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_120 <= n17150;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_120 <= n17156;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_120 <= n17162;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_120 <= n17168;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_120 <= n17174;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_120 <= n17180;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_120 <= n17186;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_120 <= n17192;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_120 <= n17198;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_120 <= n17204;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_120 <= n17210;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_120 <= n17216;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_121 <= n17222;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_121 <= n17228;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_121 <= n17234;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_121 <= n17240;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_121 <= n17246;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_121 <= n17252;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_121 <= n17258;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_121 <= n17264;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_121 <= n17270;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_121 <= n17276;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_121 <= n17282;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_121 <= n17288;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_121 <= n17294;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_121 <= n17300;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_121 <= n17306;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_122 <= n17312;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_122 <= n17318;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_122 <= n17324;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_122 <= n17330;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_122 <= n17336;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_122 <= n17342;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_122 <= n17348;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_122 <= n17354;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_122 <= n17360;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_122 <= n17366;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_122 <= n17372;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_122 <= n17378;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_122 <= n17384;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_122 <= n17390;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_122 <= n17396;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_123 <= n17402;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_123 <= n17408;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_123 <= n17414;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_123 <= n17420;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_123 <= n17426;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_123 <= n17432;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_123 <= n17438;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_123 <= n17444;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_123 <= n17450;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_123 <= n17456;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_123 <= n17462;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_123 <= n17468;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_123 <= n17474;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_123 <= n17480;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_123 <= n17486;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_124 <= n17492;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_124 <= n17498;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_124 <= n17504;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_124 <= n17510;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_124 <= n17516;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_124 <= n17522;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_124 <= n17528;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_124 <= n17534;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_124 <= n17540;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_124 <= n17546;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_124 <= n17552;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_124 <= n17558;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_124 <= n17564;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_124 <= n17570;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_124 <= n17576;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_125 <= n17582;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_125 <= n17588;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_125 <= n17594;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_125 <= n17600;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_125 <= n17606;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_125 <= n17612;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_125 <= n17618;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_125 <= n17624;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_125 <= n17630;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_125 <= n17636;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_125 <= n17642;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_125 <= n17648;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_125 <= n17654;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_125 <= n17660;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_125 <= n17666;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_126 <= n17672;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_126 <= n17678;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_126 <= n17684;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_126 <= n17690;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_126 <= n17696;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_126 <= n17702;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_126 <= n17708;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_126 <= n17714;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_126 <= n17720;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_126 <= n17726;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_126 <= n17732;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_126 <= n17738;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_126 <= n17744;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_126 <= n17750;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_126 <= n17756;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_127 <= n17762;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_127 <= n17768;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_127 <= n17774;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_127 <= n17780;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_127 <= n17786;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_127 <= n17792;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_127 <= n17798;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_127 <= n17804;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_127 <= n17810;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_127 <= n17816;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_127 <= n17822;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_127 <= n17828;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_127 <= n17834;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_127 <= n17840;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_127 <= n17846;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_128 <= n17852;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_128 <= n17858;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_128 <= n17864;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_128 <= n17870;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_128 <= n17876;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_128 <= n17882;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_128 <= n17888;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_128 <= n17894;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_128 <= n17900;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_128 <= n17906;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_128 <= n17912;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_128 <= n17918;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_128 <= n17924;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_128 <= n17930;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_128 <= n17936;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_129 <= n17942;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_129 <= n17948;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_129 <= n17954;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_129 <= n17960;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_129 <= n17966;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_129 <= n17972;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_129 <= n17978;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_129 <= n17984;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_129 <= n17990;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_129 <= n17996;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_129 <= n18002;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_129 <= n18008;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_129 <= n18014;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_129 <= n18020;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_129 <= n18026;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_130 <= n18032;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_130 <= n18038;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_130 <= n18044;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_130 <= n18050;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_130 <= n18056;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_130 <= n18062;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_130 <= n18068;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_130 <= n18074;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_130 <= n18080;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_130 <= n18086;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_130 <= n18092;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_130 <= n18098;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_130 <= n18104;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_130 <= n18110;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_130 <= n18116;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_131 <= n18122;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_131 <= n18128;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_131 <= n18134;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_131 <= n18140;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_131 <= n18146;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_131 <= n18152;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_131 <= n18158;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_131 <= n18164;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_131 <= n18170;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_131 <= n18176;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_131 <= n18182;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_131 <= n18188;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_131 <= n18194;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_131 <= n18200;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_131 <= n18206;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_132 <= n18212;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_132 <= n18218;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_132 <= n18224;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_132 <= n18230;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_132 <= n18236;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_132 <= n18242;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_132 <= n18248;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_132 <= n18254;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_132 <= n18260;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_132 <= n18266;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_132 <= n18272;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_132 <= n18278;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_132 <= n18284;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_132 <= n18290;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_132 <= n18296;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_133 <= n18302;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_133 <= n18308;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_133 <= n18314;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_133 <= n18320;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_133 <= n18326;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_133 <= n18332;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_133 <= n18338;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_133 <= n18344;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_133 <= n18350;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_133 <= n18356;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_133 <= n18362;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_133 <= n18368;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_133 <= n18374;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_133 <= n18380;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_133 <= n18386;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_134 <= n18392;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_134 <= n18398;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_134 <= n18404;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_134 <= n18410;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_134 <= n18416;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_134 <= n18422;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_134 <= n18428;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_134 <= n18434;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_134 <= n18440;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_134 <= n18446;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_134 <= n18452;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_134 <= n18458;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_134 <= n18464;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_134 <= n18470;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_134 <= n18476;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_135 <= n18482;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_135 <= n18488;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_135 <= n18494;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_135 <= n18500;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_135 <= n18506;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_135 <= n18512;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_135 <= n18518;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_135 <= n18524;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_135 <= n18530;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_135 <= n18536;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_135 <= n18542;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_135 <= n18548;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_135 <= n18554;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_135 <= n18560;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_135 <= n18566;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_136 <= n18572;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_136 <= n18578;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_136 <= n18584;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_136 <= n18590;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_136 <= n18596;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_136 <= n18602;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_136 <= n18608;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_136 <= n18614;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_136 <= n18620;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_136 <= n18626;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_136 <= n18632;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_136 <= n18638;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_136 <= n18644;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_136 <= n18650;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_136 <= n18656;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_137 <= n18662;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_137 <= n18668;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_137 <= n18674;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_137 <= n18680;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_137 <= n18686;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_137 <= n18692;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_137 <= n18698;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_137 <= n18704;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_137 <= n18710;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_137 <= n18716;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_137 <= n18722;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_137 <= n18728;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_137 <= n18734;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_137 <= n18740;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_137 <= n18746;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_138 <= n18752;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_138 <= n18758;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_138 <= n18764;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_138 <= n18770;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_138 <= n18776;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_138 <= n18782;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_138 <= n18788;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_138 <= n18794;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_138 <= n18800;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_138 <= n18806;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_138 <= n18812;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_138 <= n18818;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_138 <= n18824;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_138 <= n18830;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_138 <= n18836;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_139 <= n18842;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_139 <= n18848;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_139 <= n18854;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_139 <= n18860;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_139 <= n18866;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_139 <= n18872;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_139 <= n18878;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_139 <= n18884;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_139 <= n18890;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_139 <= n18896;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_139 <= n18902;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_139 <= n18908;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_139 <= n18914;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_139 <= n18920;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_139 <= n18926;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_140 <= n18932;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_140 <= n18938;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_140 <= n18944;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_140 <= n18950;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_140 <= n18956;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_140 <= n18962;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_140 <= n18968;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_140 <= n18974;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_140 <= n18980;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_140 <= n18986;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_140 <= n18992;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_140 <= n18998;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_140 <= n19004;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_140 <= n19010;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_140 <= n19016;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_141 <= n19022;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_141 <= n19028;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_141 <= n19034;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_141 <= n19040;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_141 <= n19046;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_141 <= n19052;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_141 <= n19058;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_141 <= n19064;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_141 <= n19070;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_141 <= n19076;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_141 <= n19082;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_141 <= n19088;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_141 <= n19094;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_141 <= n19100;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_141 <= n19106;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_142 <= n19112;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_142 <= n19118;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_142 <= n19124;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_142 <= n19130;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_142 <= n19136;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_142 <= n19142;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_142 <= n19148;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_142 <= n19154;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_142 <= n19160;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_142 <= n19166;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_142 <= n19172;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_142 <= n19178;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_142 <= n19184;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_142 <= n19190;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_142 <= n19196;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_143 <= n19202;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_143 <= n19208;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_143 <= n19214;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_143 <= n19220;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_143 <= n19226;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_143 <= n19232;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_143 <= n19238;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_143 <= n19244;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_143 <= n19250;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_143 <= n19256;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_143 <= n19262;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_143 <= n19268;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_143 <= n19274;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_143 <= n19280;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_143 <= n19286;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_144 <= n19292;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_144 <= n19298;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_144 <= n19304;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_144 <= n19310;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_144 <= n19316;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_144 <= n19322;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_144 <= n19328;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_144 <= n19334;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_144 <= n19340;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_144 <= n19346;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_144 <= n19352;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_144 <= n19358;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_144 <= n19364;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_144 <= n19370;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_144 <= n19376;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_145 <= n19382;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_145 <= n19388;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_145 <= n19394;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_145 <= n19400;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_145 <= n19406;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_145 <= n19412;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_145 <= n19418;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_145 <= n19424;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_145 <= n19430;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_145 <= n19436;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_145 <= n19442;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_145 <= n19448;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_145 <= n19454;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_145 <= n19460;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_145 <= n19466;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_146 <= n19472;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_146 <= n19478;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_146 <= n19484;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_146 <= n19490;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_146 <= n19496;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_146 <= n19502;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_146 <= n19508;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_146 <= n19514;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_146 <= n19520;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_146 <= n19526;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_146 <= n19532;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_146 <= n19538;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_146 <= n19544;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_146 <= n19550;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_146 <= n19556;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_147 <= n19562;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_147 <= n19568;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_147 <= n19574;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_147 <= n19580;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_147 <= n19586;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_147 <= n19592;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_147 <= n19598;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_147 <= n19604;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_147 <= n19610;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_147 <= n19616;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_147 <= n19622;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_147 <= n19628;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_147 <= n19634;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_147 <= n19640;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_147 <= n19646;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_148 <= n19652;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_148 <= n19658;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_148 <= n19664;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_148 <= n19670;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_148 <= n19676;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_148 <= n19682;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_148 <= n19688;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_148 <= n19694;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_148 <= n19700;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_148 <= n19706;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_148 <= n19712;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_148 <= n19718;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_148 <= n19724;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_148 <= n19730;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_148 <= n19736;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_149 <= n19742;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_149 <= n19748;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_149 <= n19754;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_149 <= n19760;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_149 <= n19766;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_149 <= n19772;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_149 <= n19778;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_149 <= n19784;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_149 <= n19790;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_149 <= n19796;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_149 <= n19802;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_149 <= n19808;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_149 <= n19814;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_149 <= n19820;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_149 <= n19826;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_150 <= n19832;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_150 <= n19838;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_150 <= n19844;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_150 <= n19850;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_150 <= n19856;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_150 <= n19862;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_150 <= n19868;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_150 <= n19874;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_150 <= n19880;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_150 <= n19886;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_150 <= n19892;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_150 <= n19898;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_150 <= n19904;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_150 <= n19910;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_150 <= n19916;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_151 <= n19922;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_151 <= n19928;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_151 <= n19934;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_151 <= n19940;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_151 <= n19946;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_151 <= n19952;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_151 <= n19958;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_151 <= n19964;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_151 <= n19970;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_151 <= n19976;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_151 <= n19982;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_151 <= n19988;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_151 <= n19994;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_151 <= n20000;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_151 <= n20006;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_152 <= n20012;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_152 <= n20018;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_152 <= n20024;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_152 <= n20030;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_152 <= n20036;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_152 <= n20042;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_152 <= n20048;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_152 <= n20054;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_152 <= n20060;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_152 <= n20066;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_152 <= n20072;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_152 <= n20078;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_152 <= n20084;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_152 <= n20090;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_152 <= n20096;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_153 <= n20102;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_153 <= n20108;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_153 <= n20114;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_153 <= n20120;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_153 <= n20126;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_153 <= n20132;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_153 <= n20138;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_153 <= n20144;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_153 <= n20150;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_153 <= n20156;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_153 <= n20162;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_153 <= n20168;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_153 <= n20174;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_153 <= n20180;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_153 <= n20186;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_154 <= n20192;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_154 <= n20198;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_154 <= n20204;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_154 <= n20210;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_154 <= n20216;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_154 <= n20222;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_154 <= n20228;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_154 <= n20234;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_154 <= n20240;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_154 <= n20246;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_154 <= n20252;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_154 <= n20258;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_154 <= n20264;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_154 <= n20270;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_154 <= n20276;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_155 <= n20282;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_155 <= n20288;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_155 <= n20294;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_155 <= n20300;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_155 <= n20306;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_155 <= n20312;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_155 <= n20318;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_155 <= n20324;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_155 <= n20330;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_155 <= n20336;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_155 <= n20342;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_155 <= n20348;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_155 <= n20354;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_155 <= n20360;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_155 <= n20366;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_156 <= n20372;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_156 <= n20378;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_156 <= n20384;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_156 <= n20390;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_156 <= n20396;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_156 <= n20402;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_156 <= n20408;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_156 <= n20414;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_156 <= n20420;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_156 <= n20426;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_156 <= n20432;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_156 <= n20438;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_156 <= n20444;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_156 <= n20450;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_156 <= n20456;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_157 <= n20462;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_157 <= n20468;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_157 <= n20474;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_157 <= n20480;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_157 <= n20486;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_157 <= n20492;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_157 <= n20498;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_157 <= n20504;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_157 <= n20510;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_157 <= n20516;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_157 <= n20522;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_157 <= n20528;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_157 <= n20534;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_157 <= n20540;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_157 <= n20546;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_158 <= n20552;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_158 <= n20558;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_158 <= n20564;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_158 <= n20570;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_158 <= n20576;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_158 <= n20582;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_158 <= n20588;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_158 <= n20594;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_158 <= n20600;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_158 <= n20606;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_158 <= n20612;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_158 <= n20618;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_158 <= n20624;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_158 <= n20630;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_158 <= n20636;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_159 <= n20642;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_159 <= n20648;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_159 <= n20654;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_159 <= n20660;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_159 <= n20666;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_159 <= n20672;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_159 <= n20678;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_159 <= n20684;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_159 <= n20690;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_159 <= n20696;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_159 <= n20702;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_159 <= n20708;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_159 <= n20714;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_159 <= n20720;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_159 <= n20726;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_160 <= n20732;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_160 <= n20738;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_160 <= n20744;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_160 <= n20750;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_160 <= n20756;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_160 <= n20762;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_160 <= n20768;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_160 <= n20774;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_160 <= n20780;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_160 <= n20786;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_160 <= n20792;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_160 <= n20798;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_160 <= n20804;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_160 <= n20810;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_160 <= n20816;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_161 <= n20822;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_161 <= n20828;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_161 <= n20834;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_161 <= n20840;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_161 <= n20846;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_161 <= n20852;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_161 <= n20858;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_161 <= n20864;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_161 <= n20870;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_161 <= n20876;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_161 <= n20882;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_161 <= n20888;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_161 <= n20894;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_161 <= n20900;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_161 <= n20906;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_162 <= n20912;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_162 <= n20918;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_162 <= n20924;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_162 <= n20930;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_162 <= n20936;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_162 <= n20942;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_162 <= n20948;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_162 <= n20954;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_162 <= n20960;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_162 <= n20966;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_162 <= n20972;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_162 <= n20978;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_162 <= n20984;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_162 <= n20990;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_162 <= n20996;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_163 <= n21002;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_163 <= n21008;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_163 <= n21014;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_163 <= n21020;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_163 <= n21026;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_163 <= n21032;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_163 <= n21038;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_163 <= n21044;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_163 <= n21050;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_163 <= n21056;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_163 <= n21062;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_163 <= n21068;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_163 <= n21074;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_163 <= n21080;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_163 <= n21086;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_164 <= n21092;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_164 <= n21098;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_164 <= n21104;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_164 <= n21110;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_164 <= n21116;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_164 <= n21122;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_164 <= n21128;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_164 <= n21134;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_164 <= n21140;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_164 <= n21146;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_164 <= n21152;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_164 <= n21158;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_164 <= n21164;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_164 <= n21170;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_164 <= n21176;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_165 <= n21182;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_165 <= n21188;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_165 <= n21194;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_165 <= n21200;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_165 <= n21206;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_165 <= n21212;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_165 <= n21218;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_165 <= n21224;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_165 <= n21230;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_165 <= n21236;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_165 <= n21242;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_165 <= n21248;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_165 <= n21254;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_165 <= n21260;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_165 <= n21266;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_166 <= n21272;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_166 <= n21278;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_166 <= n21284;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_166 <= n21290;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_166 <= n21296;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_166 <= n21302;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_166 <= n21308;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_166 <= n21314;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_166 <= n21320;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_166 <= n21326;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_166 <= n21332;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_166 <= n21338;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_166 <= n21344;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_166 <= n21350;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_166 <= n21356;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_167 <= n21362;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_167 <= n21368;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_167 <= n21374;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_167 <= n21380;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_167 <= n21386;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_167 <= n21392;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_167 <= n21398;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_167 <= n21404;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_167 <= n21410;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_167 <= n21416;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_167 <= n21422;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_167 <= n21428;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_167 <= n21434;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_167 <= n21440;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_167 <= n21446;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_168 <= n21452;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_168 <= n21458;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_168 <= n21464;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_168 <= n21470;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_168 <= n21476;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_168 <= n21482;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_168 <= n21488;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_168 <= n21494;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_168 <= n21500;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_168 <= n21506;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_168 <= n21512;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_168 <= n21518;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_168 <= n21524;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_168 <= n21530;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_168 <= n21536;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_169 <= n21542;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_169 <= n21548;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_169 <= n21554;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_169 <= n21560;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_169 <= n21566;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_169 <= n21572;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_169 <= n21578;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_169 <= n21584;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_169 <= n21590;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_169 <= n21596;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_169 <= n21602;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_169 <= n21608;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_169 <= n21614;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_169 <= n21620;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_169 <= n21626;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_170 <= n21632;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_170 <= n21638;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_170 <= n21644;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_170 <= n21650;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_170 <= n21656;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_170 <= n21662;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_170 <= n21668;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_170 <= n21674;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_170 <= n21680;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_170 <= n21686;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_170 <= n21692;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_170 <= n21698;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_170 <= n21704;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_170 <= n21710;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_170 <= n21716;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_171 <= n21722;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_171 <= n21728;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_171 <= n21734;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_171 <= n21740;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_171 <= n21746;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_171 <= n21752;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_171 <= n21758;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_171 <= n21764;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_171 <= n21770;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_171 <= n21776;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_171 <= n21782;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_171 <= n21788;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_171 <= n21794;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_171 <= n21800;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_171 <= n21806;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_172 <= n21812;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_172 <= n21818;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_172 <= n21824;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_172 <= n21830;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_172 <= n21836;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_172 <= n21842;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_172 <= n21848;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_172 <= n21854;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_172 <= n21860;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_172 <= n21866;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_172 <= n21872;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_172 <= n21878;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_172 <= n21884;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_172 <= n21890;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_172 <= n21896;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_173 <= n21902;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_173 <= n21908;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_173 <= n21914;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_173 <= n21920;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_173 <= n21926;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_173 <= n21932;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_173 <= n21938;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_173 <= n21944;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_173 <= n21950;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_173 <= n21956;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_173 <= n21962;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_173 <= n21968;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_173 <= n21974;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_173 <= n21980;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_173 <= n21986;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_174 <= n21992;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_174 <= n21998;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_174 <= n22004;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_174 <= n22010;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_174 <= n22016;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_174 <= n22022;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_174 <= n22028;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_174 <= n22034;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_174 <= n22040;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_174 <= n22046;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_174 <= n22052;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_174 <= n22058;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_174 <= n22064;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_174 <= n22070;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_174 <= n22076;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_175 <= n22082;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_175 <= n22088;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_175 <= n22094;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_175 <= n22100;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_175 <= n22106;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_175 <= n22112;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_175 <= n22118;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_175 <= n22124;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_175 <= n22130;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_175 <= n22136;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_175 <= n22142;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_175 <= n22148;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_175 <= n22154;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_175 <= n22160;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_175 <= n22166;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_176 <= n22172;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_176 <= n22178;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_176 <= n22184;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_176 <= n22190;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_176 <= n22196;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_176 <= n22202;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_176 <= n22208;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_176 <= n22214;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_176 <= n22220;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_176 <= n22226;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_176 <= n22232;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_176 <= n22238;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_176 <= n22244;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_176 <= n22250;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_176 <= n22256;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_177 <= n22262;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_177 <= n22268;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_177 <= n22274;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_177 <= n22280;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_177 <= n22286;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_177 <= n22292;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_177 <= n22298;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_177 <= n22304;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_177 <= n22310;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_177 <= n22316;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_177 <= n22322;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_177 <= n22328;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_177 <= n22334;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_177 <= n22340;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_177 <= n22346;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_178 <= n22352;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_178 <= n22358;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_178 <= n22364;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_178 <= n22370;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_178 <= n22376;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_178 <= n22382;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_178 <= n22388;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_178 <= n22394;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_178 <= n22400;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_178 <= n22406;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_178 <= n22412;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_178 <= n22418;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_178 <= n22424;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_178 <= n22430;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_178 <= n22436;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_179 <= n22442;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_179 <= n22448;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_179 <= n22454;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_179 <= n22460;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_179 <= n22466;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_179 <= n22472;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_179 <= n22478;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_179 <= n22484;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_179 <= n22490;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_179 <= n22496;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_179 <= n22502;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_179 <= n22508;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_179 <= n22514;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_179 <= n22520;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_179 <= n22526;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_180 <= n22532;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_180 <= n22538;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_180 <= n22544;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_180 <= n22550;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_180 <= n22556;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_180 <= n22562;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_180 <= n22568;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_180 <= n22574;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_180 <= n22580;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_180 <= n22586;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_180 <= n22592;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_180 <= n22598;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_180 <= n22604;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_180 <= n22610;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_180 <= n22616;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_181 <= n22622;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_181 <= n22628;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_181 <= n22634;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_181 <= n22640;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_181 <= n22646;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_181 <= n22652;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_181 <= n22658;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_181 <= n22664;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_181 <= n22670;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_181 <= n22676;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_181 <= n22682;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_181 <= n22688;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_181 <= n22694;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_181 <= n22700;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_181 <= n22706;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_182 <= n22712;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_182 <= n22718;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_182 <= n22724;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_182 <= n22730;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_182 <= n22736;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_182 <= n22742;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_182 <= n22748;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_182 <= n22754;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_182 <= n22760;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_182 <= n22766;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_182 <= n22772;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_182 <= n22778;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_182 <= n22784;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_182 <= n22790;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_182 <= n22796;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_183 <= n22802;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_183 <= n22808;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_183 <= n22814;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_183 <= n22820;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_183 <= n22826;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_183 <= n22832;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_183 <= n22838;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_183 <= n22844;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_183 <= n22850;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_183 <= n22856;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_183 <= n22862;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_183 <= n22868;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_183 <= n22874;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_183 <= n22880;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_183 <= n22886;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_184 <= n22892;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_184 <= n22898;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_184 <= n22904;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_184 <= n22910;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_184 <= n22916;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_184 <= n22922;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_184 <= n22928;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_184 <= n22934;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_184 <= n22940;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_184 <= n22946;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_184 <= n22952;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_184 <= n22958;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_184 <= n22964;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_184 <= n22970;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_184 <= n22976;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_185 <= n22982;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_185 <= n22988;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_185 <= n22994;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_185 <= n23000;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_185 <= n23006;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_185 <= n23012;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_185 <= n23018;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_185 <= n23024;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_185 <= n23030;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_185 <= n23036;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_185 <= n23042;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_185 <= n23048;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_185 <= n23054;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_185 <= n23060;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_185 <= n23066;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_186 <= n23072;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_186 <= n23078;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_186 <= n23084;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_186 <= n23090;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_186 <= n23096;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_186 <= n23102;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_186 <= n23108;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_186 <= n23114;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_186 <= n23120;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_186 <= n23126;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_186 <= n23132;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_186 <= n23138;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_186 <= n23144;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_186 <= n23150;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_186 <= n23156;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_187 <= n23162;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_187 <= n23168;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_187 <= n23174;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_187 <= n23180;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_187 <= n23186;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_187 <= n23192;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_187 <= n23198;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_187 <= n23204;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_187 <= n23210;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_187 <= n23216;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_187 <= n23222;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_187 <= n23228;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_187 <= n23234;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_187 <= n23240;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_187 <= n23246;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_188 <= n23252;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_188 <= n23258;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_188 <= n23264;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_188 <= n23270;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_188 <= n23276;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_188 <= n23282;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_188 <= n23288;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_188 <= n23294;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_188 <= n23300;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_188 <= n23306;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_188 <= n23312;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_188 <= n23318;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_188 <= n23324;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_188 <= n23330;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_188 <= n23336;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_189 <= n23342;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_189 <= n23348;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_189 <= n23354;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_189 <= n23360;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_189 <= n23366;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_189 <= n23372;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_189 <= n23378;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_189 <= n23384;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_189 <= n23390;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_189 <= n23396;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_189 <= n23402;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_189 <= n23408;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_189 <= n23414;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_189 <= n23420;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_189 <= n23426;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_190 <= n23432;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_190 <= n23438;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_190 <= n23444;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_190 <= n23450;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_190 <= n23456;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_190 <= n23462;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_190 <= n23468;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_190 <= n23474;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_190 <= n23480;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_190 <= n23486;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_190 <= n23492;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_190 <= n23498;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_190 <= n23504;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_190 <= n23510;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_190 <= n23516;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_191 <= n23522;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_191 <= n23528;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_191 <= n23534;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_191 <= n23540;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_191 <= n23546;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_191 <= n23552;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_191 <= n23558;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_191 <= n23564;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_191 <= n23570;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_191 <= n23576;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_191 <= n23582;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_191 <= n23588;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_191 <= n23594;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_191 <= n23600;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_191 <= n23606;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_192 <= n23612;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_192 <= n23618;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_192 <= n23624;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_192 <= n23630;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_192 <= n23636;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_192 <= n23642;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_192 <= n23648;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_192 <= n23654;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_192 <= n23660;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_192 <= n23666;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_192 <= n23672;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_192 <= n23678;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_192 <= n23684;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_192 <= n23690;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_192 <= n23696;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_193 <= n23702;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_193 <= n23708;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_193 <= n23714;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_193 <= n23720;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_193 <= n23726;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_193 <= n23732;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_193 <= n23738;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_193 <= n23744;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_193 <= n23750;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_193 <= n23756;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_193 <= n23762;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_193 <= n23768;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_193 <= n23774;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_193 <= n23780;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_193 <= n23786;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_194 <= n23792;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_194 <= n23798;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_194 <= n23804;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_194 <= n23810;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_194 <= n23816;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_194 <= n23822;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_194 <= n23828;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_194 <= n23834;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_194 <= n23840;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_194 <= n23846;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_194 <= n23852;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_194 <= n23858;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_194 <= n23864;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_194 <= n23870;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_194 <= n23876;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_195 <= n23882;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_195 <= n23888;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_195 <= n23894;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_195 <= n23900;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_195 <= n23906;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_195 <= n23912;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_195 <= n23918;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_195 <= n23924;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_195 <= n23930;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_195 <= n23936;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_195 <= n23942;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_195 <= n23948;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_195 <= n23954;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_195 <= n23960;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_195 <= n23966;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_196 <= n23972;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_196 <= n23978;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_196 <= n23984;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_196 <= n23990;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_196 <= n23996;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_196 <= n24002;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_196 <= n24008;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_196 <= n24014;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_196 <= n24020;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_196 <= n24026;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_196 <= n24032;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_196 <= n24038;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_196 <= n24044;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_196 <= n24050;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_196 <= n24056;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_197 <= n24062;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_197 <= n24068;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_197 <= n24074;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_197 <= n24080;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_197 <= n24086;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_197 <= n24092;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_197 <= n24098;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_197 <= n24104;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_197 <= n24110;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_197 <= n24116;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_197 <= n24122;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_197 <= n24128;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_197 <= n24134;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_197 <= n24140;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_197 <= n24146;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_198 <= n24152;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_198 <= n24158;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_198 <= n24164;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_198 <= n24170;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_198 <= n24176;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_198 <= n24182;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_198 <= n24188;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_198 <= n24194;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_198 <= n24200;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_198 <= n24206;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_198 <= n24212;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_198 <= n24218;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_198 <= n24224;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_198 <= n24230;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_198 <= n24236;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_199 <= n24242;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_199 <= n24248;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_199 <= n24254;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_199 <= n24260;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_199 <= n24266;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_199 <= n24272;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_199 <= n24278;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_199 <= n24284;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_199 <= n24290;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_199 <= n24296;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_199 <= n24302;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_199 <= n24308;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_199 <= n24314;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_199 <= n24320;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_199 <= n24326;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_200 <= n24332;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_200 <= n24338;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_200 <= n24344;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_200 <= n24350;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_200 <= n24356;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_200 <= n24362;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_200 <= n24368;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_200 <= n24374;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_200 <= n24380;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_200 <= n24386;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_200 <= n24392;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_200 <= n24398;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_200 <= n24404;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_200 <= n24410;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_200 <= n24416;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_201 <= n24422;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_201 <= n24428;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_201 <= n24434;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_201 <= n24440;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_201 <= n24446;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_201 <= n24452;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_201 <= n24458;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_201 <= n24464;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_201 <= n24470;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_201 <= n24476;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_201 <= n24482;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_201 <= n24488;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_201 <= n24494;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_201 <= n24500;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_201 <= n24506;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_202 <= n24512;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_202 <= n24518;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_202 <= n24524;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_202 <= n24530;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_202 <= n24536;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_202 <= n24542;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_202 <= n24548;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_202 <= n24554;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_202 <= n24560;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_202 <= n24566;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_202 <= n24572;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_202 <= n24578;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_202 <= n24584;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_202 <= n24590;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_202 <= n24596;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_203 <= n24602;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_203 <= n24608;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_203 <= n24614;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_203 <= n24620;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_203 <= n24626;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_203 <= n24632;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_203 <= n24638;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_203 <= n24644;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_203 <= n24650;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_203 <= n24656;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_203 <= n24662;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_203 <= n24668;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_203 <= n24674;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_203 <= n24680;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_203 <= n24686;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_204 <= n24692;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_204 <= n24698;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_204 <= n24704;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_204 <= n24710;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_204 <= n24716;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_204 <= n24722;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_204 <= n24728;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_204 <= n24734;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_204 <= n24740;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_204 <= n24746;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_204 <= n24752;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_204 <= n24758;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_204 <= n24764;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_204 <= n24770;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_204 <= n24776;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_205 <= n24782;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_205 <= n24788;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_205 <= n24794;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_205 <= n24800;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_205 <= n24806;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_205 <= n24812;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_205 <= n24818;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_205 <= n24824;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_205 <= n24830;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_205 <= n24836;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_205 <= n24842;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_205 <= n24848;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_205 <= n24854;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_205 <= n24860;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_205 <= n24866;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_206 <= n24872;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_206 <= n24878;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_206 <= n24884;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_206 <= n24890;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_206 <= n24896;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_206 <= n24902;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_206 <= n24908;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_206 <= n24914;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_206 <= n24920;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_206 <= n24926;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_206 <= n24932;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_206 <= n24938;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_206 <= n24944;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_206 <= n24950;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_206 <= n24956;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_207 <= n24962;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_207 <= n24968;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_207 <= n24974;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_207 <= n24980;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_207 <= n24986;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_207 <= n24992;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_207 <= n24998;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_207 <= n25004;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_207 <= n25010;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_207 <= n25016;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_207 <= n25022;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_207 <= n25028;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_207 <= n25034;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_207 <= n25040;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_207 <= n25046;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_208 <= n25052;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_208 <= n25058;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_208 <= n25064;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_208 <= n25070;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_208 <= n25076;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_208 <= n25082;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_208 <= n25088;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_208 <= n25094;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_208 <= n25100;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_208 <= n25106;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_208 <= n25112;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_208 <= n25118;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_208 <= n25124;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_208 <= n25130;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_208 <= n25136;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_209 <= n25142;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_209 <= n25148;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_209 <= n25154;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_209 <= n25160;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_209 <= n25166;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_209 <= n25172;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_209 <= n25178;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_209 <= n25184;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_209 <= n25190;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_209 <= n25196;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_209 <= n25202;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_209 <= n25208;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_209 <= n25214;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_209 <= n25220;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_209 <= n25226;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_210 <= n25232;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_210 <= n25238;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_210 <= n25244;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_210 <= n25250;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_210 <= n25256;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_210 <= n25262;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_210 <= n25268;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_210 <= n25274;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_210 <= n25280;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_210 <= n25286;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_210 <= n25292;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_210 <= n25298;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_210 <= n25304;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_210 <= n25310;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_210 <= n25316;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_211 <= n25322;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_211 <= n25328;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_211 <= n25334;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_211 <= n25340;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_211 <= n25346;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_211 <= n25352;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_211 <= n25358;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_211 <= n25364;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_211 <= n25370;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_211 <= n25376;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_211 <= n25382;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_211 <= n25388;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_211 <= n25394;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_211 <= n25400;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_211 <= n25406;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_212 <= n25412;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_212 <= n25418;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_212 <= n25424;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_212 <= n25430;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_212 <= n25436;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_212 <= n25442;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_212 <= n25448;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_212 <= n25454;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_212 <= n25460;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_212 <= n25466;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_212 <= n25472;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_212 <= n25478;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_212 <= n25484;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_212 <= n25490;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_212 <= n25496;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_213 <= n25502;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_213 <= n25508;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_213 <= n25514;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_213 <= n25520;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_213 <= n25526;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_213 <= n25532;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_213 <= n25538;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_213 <= n25544;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_213 <= n25550;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_213 <= n25556;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_213 <= n25562;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_213 <= n25568;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_213 <= n25574;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_213 <= n25580;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_213 <= n25586;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_214 <= n25592;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_214 <= n25598;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_214 <= n25604;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_214 <= n25610;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_214 <= n25616;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_214 <= n25622;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_214 <= n25628;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_214 <= n25634;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_214 <= n25640;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_214 <= n25646;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_214 <= n25652;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_214 <= n25658;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_214 <= n25664;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_214 <= n25670;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_214 <= n25676;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_215 <= n25682;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_215 <= n25688;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_215 <= n25694;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_215 <= n25700;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_215 <= n25706;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_215 <= n25712;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_215 <= n25718;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_215 <= n25724;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_215 <= n25730;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_215 <= n25736;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_215 <= n25742;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_215 <= n25748;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_215 <= n25754;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_215 <= n25760;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_215 <= n25766;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_216 <= n25772;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_216 <= n25778;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_216 <= n25784;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_216 <= n25790;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_216 <= n25796;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_216 <= n25802;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_216 <= n25808;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_216 <= n25814;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_216 <= n25820;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_216 <= n25826;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_216 <= n25832;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_216 <= n25838;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_216 <= n25844;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_216 <= n25850;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_216 <= n25856;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_217 <= n25862;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_217 <= n25868;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_217 <= n25874;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_217 <= n25880;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_217 <= n25886;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_217 <= n25892;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_217 <= n25898;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_217 <= n25904;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_217 <= n25910;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_217 <= n25916;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_217 <= n25922;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_217 <= n25928;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_217 <= n25934;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_217 <= n25940;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_217 <= n25946;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_218 <= n25952;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_218 <= n25958;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_218 <= n25964;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_218 <= n25970;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_218 <= n25976;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_218 <= n25982;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_218 <= n25988;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_218 <= n25994;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_218 <= n26000;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_218 <= n26006;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_218 <= n26012;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_218 <= n26018;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_218 <= n26024;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_218 <= n26030;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_218 <= n26036;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_219 <= n26042;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_219 <= n26048;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_219 <= n26054;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_219 <= n26060;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_219 <= n26066;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_219 <= n26072;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_219 <= n26078;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_219 <= n26084;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_219 <= n26090;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_219 <= n26096;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_219 <= n26102;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_219 <= n26108;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_219 <= n26114;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_219 <= n26120;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_219 <= n26126;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_220 <= n26132;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_220 <= n26138;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_220 <= n26144;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_220 <= n26150;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_220 <= n26156;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_220 <= n26162;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_220 <= n26168;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_220 <= n26174;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_220 <= n26180;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_220 <= n26186;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_220 <= n26192;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_220 <= n26198;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_220 <= n26204;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_220 <= n26210;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_220 <= n26216;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_221 <= n26222;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_221 <= n26228;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_221 <= n26234;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_221 <= n26240;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_221 <= n26246;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_221 <= n26252;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_221 <= n26258;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_221 <= n26264;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_221 <= n26270;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_221 <= n26276;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_221 <= n26282;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_221 <= n26288;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_221 <= n26294;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_221 <= n26300;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_221 <= n26306;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_222 <= n26312;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_222 <= n26318;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_222 <= n26324;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_222 <= n26330;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_222 <= n26336;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_222 <= n26342;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_222 <= n26348;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_222 <= n26354;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_222 <= n26360;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_222 <= n26366;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_222 <= n26372;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_222 <= n26378;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_222 <= n26384;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_222 <= n26390;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_222 <= n26396;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_223 <= n26402;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_223 <= n26408;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_223 <= n26414;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_223 <= n26420;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_223 <= n26426;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_223 <= n26432;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_223 <= n26438;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_223 <= n26444;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_223 <= n26450;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_223 <= n26456;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_223 <= n26462;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_223 <= n26468;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_223 <= n26474;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_223 <= n26480;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_223 <= n26486;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_224 <= n26492;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_224 <= n26498;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_224 <= n26504;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_224 <= n26510;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_224 <= n26516;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_224 <= n26522;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_224 <= n26528;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_224 <= n26534;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_224 <= n26540;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_224 <= n26546;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_224 <= n26552;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_224 <= n26558;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_224 <= n26564;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_224 <= n26570;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_224 <= n26576;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_225 <= n26582;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_225 <= n26588;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_225 <= n26594;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_225 <= n26600;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_225 <= n26606;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_225 <= n26612;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_225 <= n26618;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_225 <= n26624;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_225 <= n26630;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_225 <= n26636;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_225 <= n26642;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_225 <= n26648;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_225 <= n26654;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_225 <= n26660;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_225 <= n26666;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_226 <= n26672;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_226 <= n26678;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_226 <= n26684;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_226 <= n26690;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_226 <= n26696;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_226 <= n26702;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_226 <= n26708;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_226 <= n26714;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_226 <= n26720;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_226 <= n26726;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_226 <= n26732;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_226 <= n26738;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_226 <= n26744;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_226 <= n26750;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_226 <= n26756;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_227 <= n26762;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_227 <= n26768;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_227 <= n26774;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_227 <= n26780;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_227 <= n26786;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_227 <= n26792;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_227 <= n26798;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_227 <= n26804;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_227 <= n26810;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_227 <= n26816;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_227 <= n26822;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_227 <= n26828;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_227 <= n26834;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_227 <= n26840;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_227 <= n26846;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_228 <= n26852;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_228 <= n26858;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_228 <= n26864;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_228 <= n26870;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_228 <= n26876;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_228 <= n26882;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_228 <= n26888;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_228 <= n26894;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_228 <= n26900;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_228 <= n26906;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_228 <= n26912;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_228 <= n26918;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_228 <= n26924;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_228 <= n26930;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_228 <= n26936;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_229 <= n26942;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_229 <= n26948;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_229 <= n26954;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_229 <= n26960;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_229 <= n26966;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_229 <= n26972;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_229 <= n26978;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_229 <= n26984;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_229 <= n26990;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_229 <= n26996;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_229 <= n27002;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_229 <= n27008;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_229 <= n27014;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_229 <= n27020;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_229 <= n27026;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_230 <= n27032;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_230 <= n27038;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_230 <= n27044;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_230 <= n27050;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_230 <= n27056;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_230 <= n27062;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_230 <= n27068;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_230 <= n27074;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_230 <= n27080;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_230 <= n27086;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_230 <= n27092;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_230 <= n27098;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_230 <= n27104;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_230 <= n27110;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_230 <= n27116;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_231 <= n27122;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_231 <= n27128;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_231 <= n27134;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_231 <= n27140;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_231 <= n27146;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_231 <= n27152;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_231 <= n27158;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_231 <= n27164;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_231 <= n27170;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_231 <= n27176;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_231 <= n27182;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_231 <= n27188;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_231 <= n27194;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_231 <= n27200;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_231 <= n27206;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_232 <= n27212;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_232 <= n27218;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_232 <= n27224;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_232 <= n27230;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_232 <= n27236;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_232 <= n27242;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_232 <= n27248;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_232 <= n27254;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_232 <= n27260;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_232 <= n27266;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_232 <= n27272;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_232 <= n27278;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_232 <= n27284;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_232 <= n27290;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_232 <= n27296;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_233 <= n27302;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_233 <= n27308;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_233 <= n27314;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_233 <= n27320;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_233 <= n27326;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_233 <= n27332;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_233 <= n27338;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_233 <= n27344;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_233 <= n27350;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_233 <= n27356;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_233 <= n27362;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_233 <= n27368;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_233 <= n27374;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_233 <= n27380;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_233 <= n27386;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_234 <= n27392;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_234 <= n27398;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_234 <= n27404;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_234 <= n27410;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_234 <= n27416;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_234 <= n27422;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_234 <= n27428;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_234 <= n27434;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_234 <= n27440;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_234 <= n27446;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_234 <= n27452;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_234 <= n27458;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_234 <= n27464;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_234 <= n27470;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_234 <= n27476;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_235 <= n27482;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_235 <= n27488;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_235 <= n27494;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_235 <= n27500;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_235 <= n27506;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_235 <= n27512;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_235 <= n27518;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_235 <= n27524;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_235 <= n27530;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_235 <= n27536;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_235 <= n27542;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_235 <= n27548;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_235 <= n27554;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_235 <= n27560;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_235 <= n27566;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_236 <= n27572;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_236 <= n27578;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_236 <= n27584;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_236 <= n27590;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_236 <= n27596;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_236 <= n27602;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_236 <= n27608;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_236 <= n27614;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_236 <= n27620;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_236 <= n27626;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_236 <= n27632;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_236 <= n27638;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_236 <= n27644;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_236 <= n27650;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_236 <= n27656;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_237 <= n27662;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_237 <= n27668;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_237 <= n27674;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_237 <= n27680;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_237 <= n27686;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_237 <= n27692;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_237 <= n27698;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_237 <= n27704;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_237 <= n27710;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_237 <= n27716;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_237 <= n27722;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_237 <= n27728;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_237 <= n27734;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_237 <= n27740;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_237 <= n27746;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_238 <= n27752;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_238 <= n27758;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_238 <= n27764;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_238 <= n27770;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_238 <= n27776;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_238 <= n27782;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_238 <= n27788;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_238 <= n27794;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_238 <= n27800;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_238 <= n27806;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_238 <= n27812;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_238 <= n27818;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_238 <= n27824;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_238 <= n27830;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_238 <= n27836;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_239 <= n27842;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_239 <= n27848;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_239 <= n27854;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_239 <= n27860;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_239 <= n27866;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_239 <= n27872;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_239 <= n27878;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_239 <= n27884;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_239 <= n27890;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_239 <= n27896;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_239 <= n27902;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_239 <= n27908;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_239 <= n27914;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_239 <= n27920;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_239 <= n27926;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_240 <= n27932;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_240 <= n27938;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_240 <= n27944;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_240 <= n27950;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_240 <= n27956;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_240 <= n27962;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_240 <= n27968;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_240 <= n27974;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_240 <= n27980;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_240 <= n27986;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_240 <= n27992;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_240 <= n27998;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_240 <= n28004;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_240 <= n28010;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_240 <= n28016;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_241 <= n28022;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_241 <= n28028;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_241 <= n28034;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_241 <= n28040;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_241 <= n28046;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_241 <= n28052;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_241 <= n28058;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_241 <= n28064;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_241 <= n28070;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_241 <= n28076;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_241 <= n28082;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_241 <= n28088;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_241 <= n28094;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_241 <= n28100;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_241 <= n28106;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_242 <= n28112;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_242 <= n28118;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_242 <= n28124;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_242 <= n28130;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_242 <= n28136;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_242 <= n28142;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_242 <= n28148;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_242 <= n28154;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_242 <= n28160;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_242 <= n28166;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_242 <= n28172;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_242 <= n28178;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_242 <= n28184;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_242 <= n28190;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_242 <= n28196;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_243 <= n28202;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_243 <= n28208;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_243 <= n28214;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_243 <= n28220;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_243 <= n28226;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_243 <= n28232;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_243 <= n28238;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_243 <= n28244;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_243 <= n28250;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_243 <= n28256;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_243 <= n28262;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_243 <= n28268;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_243 <= n28274;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_243 <= n28280;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_243 <= n28286;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_244 <= n28292;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_244 <= n28298;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_244 <= n28304;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_244 <= n28310;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_244 <= n28316;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_244 <= n28322;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_244 <= n28328;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_244 <= n28334;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_244 <= n28340;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_244 <= n28346;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_244 <= n28352;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_244 <= n28358;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_244 <= n28364;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_244 <= n28370;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_244 <= n28376;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_245 <= n28382;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_245 <= n28388;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_245 <= n28394;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_245 <= n28400;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_245 <= n28406;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_245 <= n28412;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_245 <= n28418;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_245 <= n28424;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_245 <= n28430;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_245 <= n28436;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_245 <= n28442;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_245 <= n28448;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_245 <= n28454;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_245 <= n28460;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_245 <= n28466;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_246 <= n28472;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_246 <= n28478;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_246 <= n28484;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_246 <= n28490;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_246 <= n28496;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_246 <= n28502;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_246 <= n28508;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_246 <= n28514;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_246 <= n28520;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_246 <= n28526;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_246 <= n28532;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_246 <= n28538;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_246 <= n28544;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_246 <= n28550;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_246 <= n28556;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_247 <= n28562;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_247 <= n28568;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_247 <= n28574;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_247 <= n28580;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_247 <= n28586;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_247 <= n28592;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_247 <= n28598;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_247 <= n28604;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_247 <= n28610;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_247 <= n28616;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_247 <= n28622;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_247 <= n28628;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_247 <= n28634;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_247 <= n28640;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_247 <= n28646;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_248 <= n28652;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_248 <= n28658;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_248 <= n28664;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_248 <= n28670;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_248 <= n28676;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_248 <= n28682;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_248 <= n28688;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_248 <= n28694;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_248 <= n28700;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_248 <= n28706;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_248 <= n28712;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_248 <= n28718;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_248 <= n28724;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_248 <= n28730;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_248 <= n28736;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_249 <= n28742;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_249 <= n28748;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_249 <= n28754;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_249 <= n28760;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_249 <= n28766;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_249 <= n28772;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_249 <= n28778;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_249 <= n28784;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_249 <= n28790;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_249 <= n28796;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_249 <= n28802;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_249 <= n28808;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_249 <= n28814;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_249 <= n28820;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_249 <= n28826;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_250 <= n28832;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_250 <= n28838;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_250 <= n28844;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_250 <= n28850;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_250 <= n28856;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_250 <= n28862;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_250 <= n28868;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_250 <= n28874;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_250 <= n28880;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_250 <= n28886;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_250 <= n28892;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_250 <= n28898;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_250 <= n28904;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_250 <= n28910;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_250 <= n28916;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_251 <= n28922;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_251 <= n28928;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_251 <= n28934;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_251 <= n28940;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_251 <= n28946;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_251 <= n28952;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_251 <= n28958;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_251 <= n28964;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_251 <= n28970;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_251 <= n28976;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_251 <= n28982;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_251 <= n28988;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_251 <= n28994;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_251 <= n29000;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_251 <= n29006;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_252 <= n29012;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_252 <= n29018;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_252 <= n29024;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_252 <= n29030;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_252 <= n29036;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_252 <= n29042;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_252 <= n29048;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_252 <= n29054;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_252 <= n29060;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_252 <= n29066;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_252 <= n29072;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_252 <= n29078;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_252 <= n29084;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_252 <= n29090;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_252 <= n29096;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_253 <= n29102;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_253 <= n29108;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_253 <= n29114;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_253 <= n29120;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_253 <= n29126;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_253 <= n29132;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_253 <= n29138;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_253 <= n29144;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_253 <= n29150;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_253 <= n29156;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_253 <= n29162;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_253 <= n29168;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_253 <= n29174;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_253 <= n29180;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_253 <= n29186;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_254 <= n29192;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_254 <= n29198;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_254 <= n29204;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_254 <= n29210;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_254 <= n29216;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_254 <= n29222;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_254 <= n29228;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_254 <= n29234;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_254 <= n29240;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_254 <= n29246;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_254 <= n29252;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_254 <= n29258;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_254 <= n29264;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_254 <= n29270;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_254 <= n29276;
       end
       if ( __ILA_DATAPATH_decode_of_alu_and__ && __ILA_DATAPATH_grant__[0] ) begin
           iram_255 <= n29283;
       end else if ( __ILA_DATAPATH_decode_of_alu_inc__ && __ILA_DATAPATH_grant__[1] ) begin
           iram_255 <= n29289;
       end else if ( __ILA_DATAPATH_decode_of_alu_not__ && __ILA_DATAPATH_grant__[2] ) begin
           iram_255 <= n29295;
       end else if ( __ILA_DATAPATH_decode_of_alu_da__ && __ILA_DATAPATH_grant__[3] ) begin
           iram_255 <= n29301;
       end else if ( __ILA_DATAPATH_decode_of_alu_mul__ && __ILA_DATAPATH_grant__[4] ) begin
           iram_255 <= n29307;
       end else if ( __ILA_DATAPATH_decode_of_alu_div__ && __ILA_DATAPATH_grant__[5] ) begin
           iram_255 <= n29313;
       end else if ( __ILA_DATAPATH_decode_of_alu_sub__ && __ILA_DATAPATH_grant__[6] ) begin
           iram_255 <= n29319;
       end else if ( __ILA_DATAPATH_decode_of_alu_or__ && __ILA_DATAPATH_grant__[7] ) begin
           iram_255 <= n29325;
       end else if ( __ILA_DATAPATH_decode_of_alu_rl__ && __ILA_DATAPATH_grant__[8] ) begin
           iram_255 <= n29331;
       end else if ( __ILA_DATAPATH_decode_of_alu_rlc__ && __ILA_DATAPATH_grant__[9] ) begin
           iram_255 <= n29337;
       end else if ( __ILA_DATAPATH_decode_of_alu_rr__ && __ILA_DATAPATH_grant__[10] ) begin
           iram_255 <= n29343;
       end else if ( __ILA_DATAPATH_decode_of_alu_rrc__ && __ILA_DATAPATH_grant__[11] ) begin
           iram_255 <= n29349;
       end else if ( __ILA_DATAPATH_decode_of_alu_xch__ && __ILA_DATAPATH_grant__[12] ) begin
           iram_255 <= n29355;
       end else if ( __ILA_DATAPATH_decode_of_alu_xor__ && __ILA_DATAPATH_grant__[13] ) begin
           iram_255 <= n29361;
       end else if ( __ILA_DATAPATH_decode_of_alu_add__ && __ILA_DATAPATH_grant__[14] ) begin
           iram_255 <= n29367;
       end
   end
end
endmodule
