module AES(
__ILA_AES_grant__,
clk,
cmd,
cmdaddr,
cmddata,
nondet_unknown0_n83,
nondet_unknown1_n86,
nondet_unknown2_n203,
rst,
__ILA_AES_acc_decode__,
__ILA_AES_decode_of_GET_STATUS__,
__ILA_AES_decode_of_READ_ADDRESS__,
__ILA_AES_decode_of_READ_COUNTER__,
__ILA_AES_decode_of_READ_KEY__,
__ILA_AES_decode_of_READ_LENGTH__,
__ILA_AES_decode_of_START_ENCRYPT__,
__ILA_AES_decode_of_WRITE_ADDRESS__,
__ILA_AES_decode_of_WRITE_COUNTER__,
__ILA_AES_decode_of_WRITE_KEY__,
__ILA_AES_decode_of_WRITE_LENGTH__,
__ILA_AES_valid__,
aes_status,
aes_address,
aes_length,
aes_counter,
aes_key,
outdata
);
input      [9:0] __ILA_AES_grant__;
input            clk;
input      [1:0] cmd;
input     [15:0] cmdaddr;
input      [7:0] cmddata;
input      [1:0] nondet_unknown0_n83;
input      [1:0] nondet_unknown1_n86;
input    [127:0] nondet_unknown2_n203;
input            rst;
output      [9:0] __ILA_AES_acc_decode__;
output            __ILA_AES_decode_of_GET_STATUS__;
output            __ILA_AES_decode_of_READ_ADDRESS__;
output            __ILA_AES_decode_of_READ_COUNTER__;
output            __ILA_AES_decode_of_READ_KEY__;
output            __ILA_AES_decode_of_READ_LENGTH__;
output            __ILA_AES_decode_of_START_ENCRYPT__;
output            __ILA_AES_decode_of_WRITE_ADDRESS__;
output            __ILA_AES_decode_of_WRITE_COUNTER__;
output            __ILA_AES_decode_of_WRITE_KEY__;
output            __ILA_AES_decode_of_WRITE_LENGTH__;
output            __ILA_AES_valid__;
output reg      [1:0] aes_status;
output reg     [15:0] aes_address;
output reg     [15:0] aes_length;
output reg    [127:0] aes_counter;
output reg    [127:0] aes_key;
output reg      [7:0] outdata;
wire      [9:0] __ILA_AES_acc_decode__;
wire            __ILA_AES_decode_of_GET_STATUS__;
wire            __ILA_AES_decode_of_READ_ADDRESS__;
wire            __ILA_AES_decode_of_READ_COUNTER__;
wire            __ILA_AES_decode_of_READ_KEY__;
wire            __ILA_AES_decode_of_READ_LENGTH__;
wire            __ILA_AES_decode_of_START_ENCRYPT__;
wire            __ILA_AES_decode_of_WRITE_ADDRESS__;
wire            __ILA_AES_decode_of_WRITE_COUNTER__;
wire            __ILA_AES_decode_of_WRITE_KEY__;
wire            __ILA_AES_decode_of_WRITE_LENGTH__;
wire      [9:0] __ILA_AES_grant__;
wire            __ILA_AES_valid__;
wire     [15:0] bv_16_0_n104;
wire     [15:0] bv_16_10_n136;
wire     [15:0] bv_16_11_n131;
wire     [15:0] bv_16_12_n126;
wire     [15:0] bv_16_13_n121;
wire     [15:0] bv_16_14_n116;
wire     [15:0] bv_16_15_n111;
wire     [15:0] bv_16_1_n99;
wire     [15:0] bv_16_2_n176;
wire     [15:0] bv_16_3_n171;
wire     [15:0] bv_16_4_n166;
wire     [15:0] bv_16_5_n161;
wire     [15:0] bv_16_65280_n15;
wire     [15:0] bv_16_65282_n6;
wire     [15:0] bv_16_65283_n89;
wire     [15:0] bv_16_65284_n11;
wire     [15:0] bv_16_65286_n26;
wire     [15:0] bv_16_65296_n46;
wire     [15:0] bv_16_65312_n37;
wire     [15:0] bv_16_65328_n42;
wire     [15:0] bv_16_6_n156;
wire     [15:0] bv_16_7_n151;
wire     [15:0] bv_16_8_n146;
wire     [15:0] bv_16_9_n141;
wire      [1:0] bv_2_0_n81;
wire      [1:0] bv_2_1_n0;
wire      [1:0] bv_2_2_n2;
wire      [7:0] bv_8_1_n18;
wire            clk;
wire      [1:0] cmd;
wire     [15:0] cmdaddr;
wire      [7:0] cmddata;
wire            n1;
wire            n10;
wire            n100;
wire      [7:0] n101;
wire      [7:0] n102;
wire     [15:0] n103;
wire            n105;
wire      [7:0] n106;
wire      [7:0] n107;
wire     [15:0] n108;
wire     [15:0] n109;
wire     [15:0] n110;
wire            n112;
wire      [7:0] n113;
wire      [7:0] n114;
wire     [15:0] n115;
wire            n117;
wire      [7:0] n118;
wire      [7:0] n119;
wire            n12;
wire     [15:0] n120;
wire            n122;
wire      [7:0] n123;
wire      [7:0] n124;
wire     [15:0] n125;
wire            n127;
wire      [7:0] n128;
wire      [7:0] n129;
wire            n13;
wire     [15:0] n130;
wire            n132;
wire      [7:0] n133;
wire      [7:0] n134;
wire     [15:0] n135;
wire            n137;
wire      [7:0] n138;
wire      [7:0] n139;
wire            n14;
wire     [15:0] n140;
wire            n142;
wire      [7:0] n143;
wire      [7:0] n144;
wire     [15:0] n145;
wire            n147;
wire      [7:0] n148;
wire      [7:0] n149;
wire     [15:0] n150;
wire            n152;
wire      [7:0] n153;
wire      [7:0] n154;
wire     [15:0] n155;
wire            n157;
wire      [7:0] n158;
wire      [7:0] n159;
wire            n16;
wire     [15:0] n160;
wire            n162;
wire      [7:0] n163;
wire      [7:0] n164;
wire     [15:0] n165;
wire            n167;
wire      [7:0] n168;
wire      [7:0] n169;
wire            n17;
wire     [15:0] n170;
wire            n172;
wire      [7:0] n173;
wire      [7:0] n174;
wire     [15:0] n175;
wire            n177;
wire      [7:0] n178;
wire      [7:0] n179;
wire     [15:0] n180;
wire            n181;
wire      [7:0] n182;
wire      [7:0] n183;
wire     [15:0] n184;
wire            n185;
wire      [7:0] n186;
wire      [7:0] n187;
wire     [15:0] n188;
wire     [23:0] n189;
wire            n19;
wire     [31:0] n190;
wire     [39:0] n191;
wire     [47:0] n192;
wire     [55:0] n193;
wire     [63:0] n194;
wire     [71:0] n195;
wire     [79:0] n196;
wire     [87:0] n197;
wire     [95:0] n198;
wire    [103:0] n199;
wire            n20;
wire    [111:0] n200;
wire    [119:0] n201;
wire    [127:0] n202;
wire    [127:0] n204;
wire    [127:0] n205;
wire     [15:0] n206;
wire            n207;
wire      [7:0] n208;
wire      [7:0] n209;
wire            n21;
wire     [15:0] n210;
wire            n211;
wire      [7:0] n212;
wire      [7:0] n213;
wire     [15:0] n214;
wire            n215;
wire      [7:0] n216;
wire      [7:0] n217;
wire     [15:0] n218;
wire            n219;
wire            n22;
wire      [7:0] n220;
wire      [7:0] n221;
wire     [15:0] n222;
wire            n223;
wire      [7:0] n224;
wire      [7:0] n225;
wire     [15:0] n226;
wire            n227;
wire      [7:0] n228;
wire      [7:0] n229;
wire            n23;
wire     [15:0] n230;
wire            n231;
wire      [7:0] n232;
wire      [7:0] n233;
wire     [15:0] n234;
wire            n235;
wire      [7:0] n236;
wire      [7:0] n237;
wire     [15:0] n238;
wire            n239;
wire            n24;
wire      [7:0] n240;
wire      [7:0] n241;
wire     [15:0] n242;
wire            n243;
wire      [7:0] n244;
wire      [7:0] n245;
wire     [15:0] n246;
wire            n247;
wire      [7:0] n248;
wire      [7:0] n249;
wire            n25;
wire     [15:0] n250;
wire            n251;
wire      [7:0] n252;
wire      [7:0] n253;
wire     [15:0] n254;
wire            n255;
wire      [7:0] n256;
wire      [7:0] n257;
wire     [15:0] n258;
wire            n259;
wire      [7:0] n260;
wire      [7:0] n261;
wire     [15:0] n262;
wire            n263;
wire      [7:0] n264;
wire      [7:0] n265;
wire     [15:0] n266;
wire            n267;
wire      [7:0] n268;
wire      [7:0] n269;
wire            n27;
wire     [15:0] n270;
wire     [23:0] n271;
wire     [31:0] n272;
wire     [39:0] n273;
wire     [47:0] n274;
wire     [55:0] n275;
wire     [63:0] n276;
wire     [71:0] n277;
wire     [79:0] n278;
wire     [87:0] n279;
wire            n28;
wire     [95:0] n280;
wire    [103:0] n281;
wire    [111:0] n282;
wire    [119:0] n283;
wire    [127:0] n284;
wire    [127:0] n285;
wire     [15:0] n286;
wire            n287;
wire      [7:0] n288;
wire      [7:0] n289;
wire            n29;
wire      [7:0] n290;
wire     [15:0] n291;
wire            n292;
wire      [7:0] n293;
wire      [7:0] n294;
wire      [7:0] n295;
wire     [15:0] n296;
wire            n297;
wire      [7:0] n298;
wire     [15:0] n299;
wire            n3;
wire            n30;
wire            n300;
wire      [7:0] n301;
wire     [15:0] n302;
wire            n303;
wire      [7:0] n304;
wire     [15:0] n305;
wire            n306;
wire      [7:0] n307;
wire     [15:0] n308;
wire            n309;
wire            n31;
wire      [7:0] n310;
wire     [15:0] n311;
wire            n312;
wire      [7:0] n313;
wire     [15:0] n314;
wire            n315;
wire      [7:0] n316;
wire     [15:0] n317;
wire            n318;
wire      [7:0] n319;
wire            n32;
wire     [15:0] n320;
wire            n321;
wire      [7:0] n322;
wire     [15:0] n323;
wire            n324;
wire      [7:0] n325;
wire     [15:0] n326;
wire            n327;
wire      [7:0] n328;
wire     [15:0] n329;
wire            n33;
wire            n330;
wire      [7:0] n331;
wire     [15:0] n332;
wire            n333;
wire      [7:0] n334;
wire     [15:0] n335;
wire            n336;
wire      [7:0] n337;
wire     [15:0] n338;
wire            n339;
wire            n34;
wire      [7:0] n340;
wire      [7:0] n341;
wire      [7:0] n342;
wire      [7:0] n343;
wire      [7:0] n344;
wire      [7:0] n345;
wire      [7:0] n346;
wire      [7:0] n347;
wire      [7:0] n348;
wire      [7:0] n349;
wire            n35;
wire      [7:0] n350;
wire      [7:0] n351;
wire      [7:0] n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire     [15:0] n357;
wire            n358;
wire      [7:0] n359;
wire            n36;
wire     [15:0] n360;
wire            n361;
wire      [7:0] n362;
wire     [15:0] n363;
wire            n364;
wire      [7:0] n365;
wire     [15:0] n366;
wire            n367;
wire      [7:0] n368;
wire     [15:0] n369;
wire            n370;
wire      [7:0] n371;
wire     [15:0] n372;
wire            n373;
wire      [7:0] n374;
wire     [15:0] n375;
wire            n376;
wire      [7:0] n377;
wire     [15:0] n378;
wire            n379;
wire            n38;
wire      [7:0] n380;
wire     [15:0] n381;
wire            n382;
wire      [7:0] n383;
wire     [15:0] n384;
wire            n385;
wire      [7:0] n386;
wire     [15:0] n387;
wire            n388;
wire      [7:0] n389;
wire            n39;
wire     [15:0] n390;
wire            n391;
wire      [7:0] n392;
wire     [15:0] n393;
wire            n394;
wire      [7:0] n395;
wire     [15:0] n396;
wire            n397;
wire      [7:0] n398;
wire     [15:0] n399;
wire            n4;
wire            n40;
wire            n400;
wire      [7:0] n401;
wire      [7:0] n402;
wire      [7:0] n403;
wire      [7:0] n404;
wire      [7:0] n405;
wire      [7:0] n406;
wire      [7:0] n407;
wire      [7:0] n408;
wire      [7:0] n409;
wire            n41;
wire      [7:0] n410;
wire      [7:0] n411;
wire      [7:0] n412;
wire      [7:0] n413;
wire      [7:0] n414;
wire      [7:0] n415;
wire      [7:0] n416;
wire      [7:0] n417;
wire     [15:0] n418;
wire            n419;
wire      [7:0] n420;
wire     [15:0] n421;
wire            n422;
wire      [7:0] n423;
wire     [15:0] n424;
wire            n425;
wire      [7:0] n426;
wire     [15:0] n427;
wire            n428;
wire      [7:0] n429;
wire            n43;
wire     [15:0] n430;
wire            n431;
wire      [7:0] n432;
wire     [15:0] n433;
wire            n434;
wire      [7:0] n435;
wire     [15:0] n436;
wire            n437;
wire      [7:0] n438;
wire     [15:0] n439;
wire            n44;
wire            n440;
wire      [7:0] n441;
wire     [15:0] n442;
wire            n443;
wire      [7:0] n444;
wire     [15:0] n445;
wire            n446;
wire      [7:0] n447;
wire     [15:0] n448;
wire            n449;
wire            n45;
wire      [7:0] n450;
wire     [15:0] n451;
wire            n452;
wire      [7:0] n453;
wire     [15:0] n454;
wire            n455;
wire      [7:0] n456;
wire     [15:0] n457;
wire            n458;
wire      [7:0] n459;
wire     [15:0] n460;
wire            n461;
wire      [7:0] n462;
wire      [7:0] n463;
wire      [7:0] n464;
wire      [7:0] n465;
wire      [7:0] n466;
wire      [7:0] n467;
wire      [7:0] n468;
wire      [7:0] n469;
wire            n47;
wire      [7:0] n470;
wire      [7:0] n471;
wire      [7:0] n472;
wire      [7:0] n473;
wire      [7:0] n474;
wire      [7:0] n475;
wire      [7:0] n476;
wire      [7:0] n477;
wire      [7:0] n478;
wire            n48;
wire            n49;
wire            n5;
wire            n50;
wire            n51;
wire            n52;
wire            n53;
wire            n54;
wire            n55;
wire            n56;
wire            n57;
wire            n58;
wire            n59;
wire            n60;
wire            n61;
wire            n62;
wire            n63;
wire            n64;
wire            n65;
wire            n66;
wire            n67;
wire            n68;
wire            n69;
wire            n7;
wire            n70;
wire            n71;
wire            n72;
wire            n73;
wire            n74;
wire            n75;
wire            n76;
wire            n77;
wire            n78;
wire            n79;
wire            n8;
wire            n80;
wire            n82;
wire      [1:0] n84;
wire      [1:0] n85;
wire      [1:0] n87;
wire      [1:0] n88;
wire            n9;
wire            n90;
wire      [7:0] n91;
wire      [7:0] n92;
wire            n93;
wire      [7:0] n94;
wire      [7:0] n95;
wire     [15:0] n96;
wire     [15:0] n97;
wire     [15:0] n98;
wire      [1:0] nondet_unknown0_n83;
wire      [1:0] nondet_unknown1_n86;
wire    [127:0] nondet_unknown2_n203;
wire            rst;
assign bv_2_1_n0 = 2'h1 ;
assign n1 =  ( cmd ) == ( bv_2_1_n0 )  ;
assign bv_2_2_n2 = 2'h2 ;
assign n3 =  ( cmd ) == ( bv_2_2_n2 )  ;
assign n4 =  ( n1 ) | ( n3 )  ;
assign __ILA_AES_valid__ = n4 ;
assign n5 =  ( cmd ) == ( bv_2_2_n2 )  ;
assign bv_16_65282_n6 = 16'hff02 ;
assign n7 =  ( cmdaddr ) == ( bv_16_65282_n6 )  ;
assign n8 =  ( cmdaddr ) > ( bv_16_65282_n6 )  ;
assign n9 =  ( n7 ) | ( n8 )  ;
assign n10 =  ( n5 ) & (n9 )  ;
assign bv_16_65284_n11 = 16'hff04 ;
assign n12 =  ( cmdaddr ) < ( bv_16_65284_n11 )  ;
assign n13 =  ( n10 ) & (n12 )  ;
assign __ILA_AES_decode_of_WRITE_ADDRESS__ = n13 ;
assign __ILA_AES_acc_decode__[0] = __ILA_AES_decode_of_WRITE_ADDRESS__ ;
assign n14 =  ( cmd ) == ( bv_2_2_n2 )  ;
assign bv_16_65280_n15 = 16'hff00 ;
assign n16 =  ( cmdaddr ) == ( bv_16_65280_n15 )  ;
assign n17 =  ( n14 ) & (n16 )  ;
assign bv_8_1_n18 = 8'h1 ;
assign n19 =  ( cmddata ) == ( bv_8_1_n18 )  ;
assign n20 =  ( n17 ) & (n19 )  ;
assign __ILA_AES_decode_of_START_ENCRYPT__ = n20 ;
assign __ILA_AES_acc_decode__[1] = __ILA_AES_decode_of_START_ENCRYPT__ ;
assign n21 =  ( cmd ) == ( bv_2_1_n0 )  ;
assign n22 =  ( cmdaddr ) == ( bv_16_65284_n11 )  ;
assign n23 =  ( cmdaddr ) > ( bv_16_65284_n11 )  ;
assign n24 =  ( n22 ) | ( n23 )  ;
assign n25 =  ( n21 ) & (n24 )  ;
assign bv_16_65286_n26 = 16'hff06 ;
assign n27 =  ( cmdaddr ) < ( bv_16_65286_n26 )  ;
assign n28 =  ( n25 ) & (n27 )  ;
assign __ILA_AES_decode_of_READ_LENGTH__ = n28 ;
assign __ILA_AES_acc_decode__[2] = __ILA_AES_decode_of_READ_LENGTH__ ;
assign n29 =  ( cmd ) == ( bv_2_1_n0 )  ;
assign n30 =  ( cmdaddr ) == ( bv_16_65282_n6 )  ;
assign n31 =  ( cmdaddr ) > ( bv_16_65282_n6 )  ;
assign n32 =  ( n30 ) | ( n31 )  ;
assign n33 =  ( n29 ) & (n32 )  ;
assign n34 =  ( cmdaddr ) < ( bv_16_65284_n11 )  ;
assign n35 =  ( n33 ) & (n34 )  ;
assign __ILA_AES_decode_of_READ_ADDRESS__ = n35 ;
assign __ILA_AES_acc_decode__[3] = __ILA_AES_decode_of_READ_ADDRESS__ ;
assign n36 =  ( cmd ) == ( bv_2_1_n0 )  ;
assign bv_16_65312_n37 = 16'hff20 ;
assign n38 =  ( cmdaddr ) == ( bv_16_65312_n37 )  ;
assign n39 =  ( cmdaddr ) > ( bv_16_65312_n37 )  ;
assign n40 =  ( n38 ) | ( n39 )  ;
assign n41 =  ( n36 ) & (n40 )  ;
assign bv_16_65328_n42 = 16'hff30 ;
assign n43 =  ( cmdaddr ) < ( bv_16_65328_n42 )  ;
assign n44 =  ( n41 ) & (n43 )  ;
assign __ILA_AES_decode_of_READ_KEY__ = n44 ;
assign __ILA_AES_acc_decode__[4] = __ILA_AES_decode_of_READ_KEY__ ;
assign n45 =  ( cmd ) == ( bv_2_1_n0 )  ;
assign bv_16_65296_n46 = 16'hff10 ;
assign n47 =  ( cmdaddr ) == ( bv_16_65296_n46 )  ;
assign n48 =  ( cmdaddr ) > ( bv_16_65296_n46 )  ;
assign n49 =  ( n47 ) | ( n48 )  ;
assign n50 =  ( n45 ) & (n49 )  ;
assign n51 =  ( cmdaddr ) < ( bv_16_65312_n37 )  ;
assign n52 =  ( n50 ) & (n51 )  ;
assign __ILA_AES_decode_of_READ_COUNTER__ = n52 ;
assign __ILA_AES_acc_decode__[5] = __ILA_AES_decode_of_READ_COUNTER__ ;
assign n53 =  ( cmd ) == ( bv_2_1_n0 )  ;
assign n54 =  ( cmdaddr ) == ( bv_16_65296_n46 )  ;
assign n55 =  ( cmdaddr ) > ( bv_16_65296_n46 )  ;
assign n56 =  ( n54 ) | ( n55 )  ;
assign n57 =  ( n53 ) & (n56 )  ;
assign n58 =  ( cmdaddr ) < ( bv_16_65312_n37 )  ;
assign n59 =  ( n57 ) & (n58 )  ;
assign __ILA_AES_decode_of_GET_STATUS__ = n59 ;
assign __ILA_AES_acc_decode__[6] = __ILA_AES_decode_of_GET_STATUS__ ;
assign n60 =  ( cmd ) == ( bv_2_2_n2 )  ;
assign n61 =  ( cmdaddr ) == ( bv_16_65284_n11 )  ;
assign n62 =  ( cmdaddr ) > ( bv_16_65284_n11 )  ;
assign n63 =  ( n61 ) | ( n62 )  ;
assign n64 =  ( n60 ) & (n63 )  ;
assign n65 =  ( cmdaddr ) < ( bv_16_65286_n26 )  ;
assign n66 =  ( n64 ) & (n65 )  ;
assign __ILA_AES_decode_of_WRITE_LENGTH__ = n66 ;
assign __ILA_AES_acc_decode__[7] = __ILA_AES_decode_of_WRITE_LENGTH__ ;
assign n67 =  ( cmd ) == ( bv_2_2_n2 )  ;
assign n68 =  ( cmdaddr ) == ( bv_16_65312_n37 )  ;
assign n69 =  ( cmdaddr ) > ( bv_16_65312_n37 )  ;
assign n70 =  ( n68 ) | ( n69 )  ;
assign n71 =  ( n67 ) & (n70 )  ;
assign n72 =  ( cmdaddr ) < ( bv_16_65328_n42 )  ;
assign n73 =  ( n71 ) & (n72 )  ;
assign __ILA_AES_decode_of_WRITE_KEY__ = n73 ;
assign __ILA_AES_acc_decode__[8] = __ILA_AES_decode_of_WRITE_KEY__ ;
assign n74 =  ( cmd ) == ( bv_2_2_n2 )  ;
assign n75 =  ( cmdaddr ) == ( bv_16_65296_n46 )  ;
assign n76 =  ( cmdaddr ) > ( bv_16_65296_n46 )  ;
assign n77 =  ( n75 ) | ( n76 )  ;
assign n78 =  ( n74 ) & (n77 )  ;
assign n79 =  ( cmdaddr ) < ( bv_16_65312_n37 )  ;
assign n80 =  ( n78 ) & (n79 )  ;
assign __ILA_AES_decode_of_WRITE_COUNTER__ = n80 ;
assign __ILA_AES_acc_decode__[9] = __ILA_AES_decode_of_WRITE_COUNTER__ ;
assign bv_2_0_n81 = 2'h0 ;
assign n82 =  ( aes_status ) == ( bv_2_0_n81 )  ;
assign n84 = nondet_unknown0_n83 ;
assign n85 =  ( n82 ) ? ( bv_2_1_n0 ) : ( n84 ) ;
assign n87 = nondet_unknown1_n86 ;
assign n88 =  ( n82 ) ? ( aes_status ) : ( n87 ) ;
assign bv_16_65283_n89 = 16'hff03 ;
assign n90 =  ( cmdaddr ) == ( bv_16_65283_n89 )  ;
assign n91 = aes_address[15:8] ;
assign n92 =  ( n90 ) ? ( cmddata ) : ( n91 ) ;
assign n93 =  ( cmdaddr ) == ( bv_16_65282_n6 )  ;
assign n94 = aes_address[7:0] ;
assign n95 =  ( n93 ) ? ( cmddata ) : ( n94 ) ;
assign n96 =  { ( n92 ) , ( n95 ) }  ;
assign n97 =  ( n82 ) ? ( n96 ) : ( aes_address ) ;
assign n98 =  ( cmdaddr ) - ( bv_16_65284_n11 )  ;
assign bv_16_1_n99 = 16'h1 ;
assign n100 =  ( n98 ) == ( bv_16_1_n99 )  ;
assign n101 = aes_length[15:8] ;
assign n102 =  ( n100 ) ? ( cmddata ) : ( n101 ) ;
assign n103 =  ( cmdaddr ) - ( bv_16_65284_n11 )  ;
assign bv_16_0_n104 = 16'h0 ;
assign n105 =  ( n103 ) == ( bv_16_0_n104 )  ;
assign n106 = aes_length[7:0] ;
assign n107 =  ( n105 ) ? ( cmddata ) : ( n106 ) ;
assign n108 =  { ( n102 ) , ( n107 ) }  ;
assign n109 =  ( n82 ) ? ( n108 ) : ( aes_length ) ;
assign n110 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign bv_16_15_n111 = 16'hf ;
assign n112 =  ( n110 ) == ( bv_16_15_n111 )  ;
assign n113 = aes_counter[127:120] ;
assign n114 =  ( n112 ) ? ( cmddata ) : ( n113 ) ;
assign n115 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign bv_16_14_n116 = 16'he ;
assign n117 =  ( n115 ) == ( bv_16_14_n116 )  ;
assign n118 = aes_counter[119:112] ;
assign n119 =  ( n117 ) ? ( cmddata ) : ( n118 ) ;
assign n120 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign bv_16_13_n121 = 16'hd ;
assign n122 =  ( n120 ) == ( bv_16_13_n121 )  ;
assign n123 = aes_counter[111:104] ;
assign n124 =  ( n122 ) ? ( cmddata ) : ( n123 ) ;
assign n125 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign bv_16_12_n126 = 16'hc ;
assign n127 =  ( n125 ) == ( bv_16_12_n126 )  ;
assign n128 = aes_counter[103:96] ;
assign n129 =  ( n127 ) ? ( cmddata ) : ( n128 ) ;
assign n130 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign bv_16_11_n131 = 16'hb ;
assign n132 =  ( n130 ) == ( bv_16_11_n131 )  ;
assign n133 = aes_counter[95:88] ;
assign n134 =  ( n132 ) ? ( cmddata ) : ( n133 ) ;
assign n135 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign bv_16_10_n136 = 16'ha ;
assign n137 =  ( n135 ) == ( bv_16_10_n136 )  ;
assign n138 = aes_counter[87:80] ;
assign n139 =  ( n137 ) ? ( cmddata ) : ( n138 ) ;
assign n140 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign bv_16_9_n141 = 16'h9 ;
assign n142 =  ( n140 ) == ( bv_16_9_n141 )  ;
assign n143 = aes_counter[79:72] ;
assign n144 =  ( n142 ) ? ( cmddata ) : ( n143 ) ;
assign n145 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign bv_16_8_n146 = 16'h8 ;
assign n147 =  ( n145 ) == ( bv_16_8_n146 )  ;
assign n148 = aes_counter[71:64] ;
assign n149 =  ( n147 ) ? ( cmddata ) : ( n148 ) ;
assign n150 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign bv_16_7_n151 = 16'h7 ;
assign n152 =  ( n150 ) == ( bv_16_7_n151 )  ;
assign n153 = aes_counter[63:56] ;
assign n154 =  ( n152 ) ? ( cmddata ) : ( n153 ) ;
assign n155 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign bv_16_6_n156 = 16'h6 ;
assign n157 =  ( n155 ) == ( bv_16_6_n156 )  ;
assign n158 = aes_counter[55:48] ;
assign n159 =  ( n157 ) ? ( cmddata ) : ( n158 ) ;
assign n160 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign bv_16_5_n161 = 16'h5 ;
assign n162 =  ( n160 ) == ( bv_16_5_n161 )  ;
assign n163 = aes_counter[47:40] ;
assign n164 =  ( n162 ) ? ( cmddata ) : ( n163 ) ;
assign n165 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign bv_16_4_n166 = 16'h4 ;
assign n167 =  ( n165 ) == ( bv_16_4_n166 )  ;
assign n168 = aes_counter[39:32] ;
assign n169 =  ( n167 ) ? ( cmddata ) : ( n168 ) ;
assign n170 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign bv_16_3_n171 = 16'h3 ;
assign n172 =  ( n170 ) == ( bv_16_3_n171 )  ;
assign n173 = aes_counter[31:24] ;
assign n174 =  ( n172 ) ? ( cmddata ) : ( n173 ) ;
assign n175 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign bv_16_2_n176 = 16'h2 ;
assign n177 =  ( n175 ) == ( bv_16_2_n176 )  ;
assign n178 = aes_counter[23:16] ;
assign n179 =  ( n177 ) ? ( cmddata ) : ( n178 ) ;
assign n180 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n181 =  ( n180 ) == ( bv_16_1_n99 )  ;
assign n182 = aes_counter[15:8] ;
assign n183 =  ( n181 ) ? ( cmddata ) : ( n182 ) ;
assign n184 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n185 =  ( n184 ) == ( bv_16_0_n104 )  ;
assign n186 = aes_counter[7:0] ;
assign n187 =  ( n185 ) ? ( cmddata ) : ( n186 ) ;
assign n188 =  { ( n183 ) , ( n187 ) }  ;
assign n189 =  { ( n179 ) , ( n188 ) }  ;
assign n190 =  { ( n174 ) , ( n189 ) }  ;
assign n191 =  { ( n169 ) , ( n190 ) }  ;
assign n192 =  { ( n164 ) , ( n191 ) }  ;
assign n193 =  { ( n159 ) , ( n192 ) }  ;
assign n194 =  { ( n154 ) , ( n193 ) }  ;
assign n195 =  { ( n149 ) , ( n194 ) }  ;
assign n196 =  { ( n144 ) , ( n195 ) }  ;
assign n197 =  { ( n139 ) , ( n196 ) }  ;
assign n198 =  { ( n134 ) , ( n197 ) }  ;
assign n199 =  { ( n129 ) , ( n198 ) }  ;
assign n200 =  { ( n124 ) , ( n199 ) }  ;
assign n201 =  { ( n119 ) , ( n200 ) }  ;
assign n202 =  { ( n114 ) , ( n201 ) }  ;
assign n204 = nondet_unknown2_n203 ;
assign n205 =  ( n82 ) ? ( n202 ) : ( n204 ) ;
assign n206 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n207 =  ( n206 ) == ( bv_16_15_n111 )  ;
assign n208 = aes_key[127:120] ;
assign n209 =  ( n207 ) ? ( cmddata ) : ( n208 ) ;
assign n210 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n211 =  ( n210 ) == ( bv_16_14_n116 )  ;
assign n212 = aes_key[119:112] ;
assign n213 =  ( n211 ) ? ( cmddata ) : ( n212 ) ;
assign n214 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n215 =  ( n214 ) == ( bv_16_13_n121 )  ;
assign n216 = aes_key[111:104] ;
assign n217 =  ( n215 ) ? ( cmddata ) : ( n216 ) ;
assign n218 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n219 =  ( n218 ) == ( bv_16_12_n126 )  ;
assign n220 = aes_key[103:96] ;
assign n221 =  ( n219 ) ? ( cmddata ) : ( n220 ) ;
assign n222 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n223 =  ( n222 ) == ( bv_16_11_n131 )  ;
assign n224 = aes_key[95:88] ;
assign n225 =  ( n223 ) ? ( cmddata ) : ( n224 ) ;
assign n226 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n227 =  ( n226 ) == ( bv_16_10_n136 )  ;
assign n228 = aes_key[87:80] ;
assign n229 =  ( n227 ) ? ( cmddata ) : ( n228 ) ;
assign n230 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n231 =  ( n230 ) == ( bv_16_9_n141 )  ;
assign n232 = aes_key[79:72] ;
assign n233 =  ( n231 ) ? ( cmddata ) : ( n232 ) ;
assign n234 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n235 =  ( n234 ) == ( bv_16_8_n146 )  ;
assign n236 = aes_key[71:64] ;
assign n237 =  ( n235 ) ? ( cmddata ) : ( n236 ) ;
assign n238 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n239 =  ( n238 ) == ( bv_16_7_n151 )  ;
assign n240 = aes_key[63:56] ;
assign n241 =  ( n239 ) ? ( cmddata ) : ( n240 ) ;
assign n242 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n243 =  ( n242 ) == ( bv_16_6_n156 )  ;
assign n244 = aes_key[55:48] ;
assign n245 =  ( n243 ) ? ( cmddata ) : ( n244 ) ;
assign n246 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n247 =  ( n246 ) == ( bv_16_5_n161 )  ;
assign n248 = aes_key[47:40] ;
assign n249 =  ( n247 ) ? ( cmddata ) : ( n248 ) ;
assign n250 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n251 =  ( n250 ) == ( bv_16_4_n166 )  ;
assign n252 = aes_key[39:32] ;
assign n253 =  ( n251 ) ? ( cmddata ) : ( n252 ) ;
assign n254 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n255 =  ( n254 ) == ( bv_16_3_n171 )  ;
assign n256 = aes_key[31:24] ;
assign n257 =  ( n255 ) ? ( cmddata ) : ( n256 ) ;
assign n258 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n259 =  ( n258 ) == ( bv_16_2_n176 )  ;
assign n260 = aes_key[23:16] ;
assign n261 =  ( n259 ) ? ( cmddata ) : ( n260 ) ;
assign n262 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n263 =  ( n262 ) == ( bv_16_1_n99 )  ;
assign n264 = aes_key[15:8] ;
assign n265 =  ( n263 ) ? ( cmddata ) : ( n264 ) ;
assign n266 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n267 =  ( n266 ) == ( bv_16_0_n104 )  ;
assign n268 = aes_key[7:0] ;
assign n269 =  ( n267 ) ? ( cmddata ) : ( n268 ) ;
assign n270 =  { ( n265 ) , ( n269 ) }  ;
assign n271 =  { ( n261 ) , ( n270 ) }  ;
assign n272 =  { ( n257 ) , ( n271 ) }  ;
assign n273 =  { ( n253 ) , ( n272 ) }  ;
assign n274 =  { ( n249 ) , ( n273 ) }  ;
assign n275 =  { ( n245 ) , ( n274 ) }  ;
assign n276 =  { ( n241 ) , ( n275 ) }  ;
assign n277 =  { ( n237 ) , ( n276 ) }  ;
assign n278 =  { ( n233 ) , ( n277 ) }  ;
assign n279 =  { ( n229 ) , ( n278 ) }  ;
assign n280 =  { ( n225 ) , ( n279 ) }  ;
assign n281 =  { ( n221 ) , ( n280 ) }  ;
assign n282 =  { ( n217 ) , ( n281 ) }  ;
assign n283 =  { ( n213 ) , ( n282 ) }  ;
assign n284 =  { ( n209 ) , ( n283 ) }  ;
assign n285 =  ( n82 ) ? ( n284 ) : ( aes_key ) ;
assign n286 =  ( cmdaddr ) - ( bv_16_65284_n11 )  ;
assign n287 =  ( n286 ) == ( bv_16_1_n99 )  ;
assign n288 = aes_length[15:8] ;
assign n289 = aes_length[7:0] ;
assign n290 =  ( n287 ) ? ( n288 ) : ( n289 ) ;
assign n291 =  ( cmdaddr ) - ( bv_16_65282_n6 )  ;
assign n292 =  ( n291 ) == ( bv_16_1_n99 )  ;
assign n293 = aes_address[15:8] ;
assign n294 = aes_address[7:0] ;
assign n295 =  ( n292 ) ? ( n293 ) : ( n294 ) ;
assign n296 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n297 =  ( n296 ) == ( bv_16_15_n111 )  ;
assign n298 = aes_key[127:120] ;
assign n299 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n300 =  ( n299 ) == ( bv_16_14_n116 )  ;
assign n301 = aes_key[119:112] ;
assign n302 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n303 =  ( n302 ) == ( bv_16_13_n121 )  ;
assign n304 = aes_key[111:104] ;
assign n305 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n306 =  ( n305 ) == ( bv_16_12_n126 )  ;
assign n307 = aes_key[103:96] ;
assign n308 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n309 =  ( n308 ) == ( bv_16_11_n131 )  ;
assign n310 = aes_key[95:88] ;
assign n311 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n312 =  ( n311 ) == ( bv_16_10_n136 )  ;
assign n313 = aes_key[87:80] ;
assign n314 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n315 =  ( n314 ) == ( bv_16_9_n141 )  ;
assign n316 = aes_key[79:72] ;
assign n317 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n318 =  ( n317 ) == ( bv_16_8_n146 )  ;
assign n319 = aes_key[71:64] ;
assign n320 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n321 =  ( n320 ) == ( bv_16_7_n151 )  ;
assign n322 = aes_key[63:56] ;
assign n323 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n324 =  ( n323 ) == ( bv_16_6_n156 )  ;
assign n325 = aes_key[55:48] ;
assign n326 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n327 =  ( n326 ) == ( bv_16_5_n161 )  ;
assign n328 = aes_key[47:40] ;
assign n329 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n330 =  ( n329 ) == ( bv_16_4_n166 )  ;
assign n331 = aes_key[39:32] ;
assign n332 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n333 =  ( n332 ) == ( bv_16_3_n171 )  ;
assign n334 = aes_key[31:24] ;
assign n335 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n336 =  ( n335 ) == ( bv_16_2_n176 )  ;
assign n337 = aes_key[23:16] ;
assign n338 =  ( cmdaddr ) - ( bv_16_65312_n37 )  ;
assign n339 =  ( n338 ) == ( bv_16_1_n99 )  ;
assign n340 = aes_key[15:8] ;
assign n341 = aes_key[7:0] ;
assign n342 =  ( n339 ) ? ( n340 ) : ( n341 ) ;
assign n343 =  ( n336 ) ? ( n337 ) : ( n342 ) ;
assign n344 =  ( n333 ) ? ( n334 ) : ( n343 ) ;
assign n345 =  ( n330 ) ? ( n331 ) : ( n344 ) ;
assign n346 =  ( n327 ) ? ( n328 ) : ( n345 ) ;
assign n347 =  ( n324 ) ? ( n325 ) : ( n346 ) ;
assign n348 =  ( n321 ) ? ( n322 ) : ( n347 ) ;
assign n349 =  ( n318 ) ? ( n319 ) : ( n348 ) ;
assign n350 =  ( n315 ) ? ( n316 ) : ( n349 ) ;
assign n351 =  ( n312 ) ? ( n313 ) : ( n350 ) ;
assign n352 =  ( n309 ) ? ( n310 ) : ( n351 ) ;
assign n353 =  ( n306 ) ? ( n307 ) : ( n352 ) ;
assign n354 =  ( n303 ) ? ( n304 ) : ( n353 ) ;
assign n355 =  ( n300 ) ? ( n301 ) : ( n354 ) ;
assign n356 =  ( n297 ) ? ( n298 ) : ( n355 ) ;
assign n357 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n358 =  ( n357 ) == ( bv_16_15_n111 )  ;
assign n359 = aes_counter[127:120] ;
assign n360 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n361 =  ( n360 ) == ( bv_16_14_n116 )  ;
assign n362 = aes_counter[119:112] ;
assign n363 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n364 =  ( n363 ) == ( bv_16_13_n121 )  ;
assign n365 = aes_counter[111:104] ;
assign n366 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n367 =  ( n366 ) == ( bv_16_12_n126 )  ;
assign n368 = aes_counter[103:96] ;
assign n369 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n370 =  ( n369 ) == ( bv_16_11_n131 )  ;
assign n371 = aes_counter[95:88] ;
assign n372 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n373 =  ( n372 ) == ( bv_16_10_n136 )  ;
assign n374 = aes_counter[87:80] ;
assign n375 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n376 =  ( n375 ) == ( bv_16_9_n141 )  ;
assign n377 = aes_counter[79:72] ;
assign n378 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n379 =  ( n378 ) == ( bv_16_8_n146 )  ;
assign n380 = aes_counter[71:64] ;
assign n381 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n382 =  ( n381 ) == ( bv_16_7_n151 )  ;
assign n383 = aes_counter[63:56] ;
assign n384 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n385 =  ( n384 ) == ( bv_16_6_n156 )  ;
assign n386 = aes_counter[55:48] ;
assign n387 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n388 =  ( n387 ) == ( bv_16_5_n161 )  ;
assign n389 = aes_counter[47:40] ;
assign n390 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n391 =  ( n390 ) == ( bv_16_4_n166 )  ;
assign n392 = aes_counter[39:32] ;
assign n393 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n394 =  ( n393 ) == ( bv_16_3_n171 )  ;
assign n395 = aes_counter[31:24] ;
assign n396 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n397 =  ( n396 ) == ( bv_16_2_n176 )  ;
assign n398 = aes_counter[23:16] ;
assign n399 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n400 =  ( n399 ) == ( bv_16_1_n99 )  ;
assign n401 = aes_counter[15:8] ;
assign n402 = aes_counter[7:0] ;
assign n403 =  ( n400 ) ? ( n401 ) : ( n402 ) ;
assign n404 =  ( n397 ) ? ( n398 ) : ( n403 ) ;
assign n405 =  ( n394 ) ? ( n395 ) : ( n404 ) ;
assign n406 =  ( n391 ) ? ( n392 ) : ( n405 ) ;
assign n407 =  ( n388 ) ? ( n389 ) : ( n406 ) ;
assign n408 =  ( n385 ) ? ( n386 ) : ( n407 ) ;
assign n409 =  ( n382 ) ? ( n383 ) : ( n408 ) ;
assign n410 =  ( n379 ) ? ( n380 ) : ( n409 ) ;
assign n411 =  ( n376 ) ? ( n377 ) : ( n410 ) ;
assign n412 =  ( n373 ) ? ( n374 ) : ( n411 ) ;
assign n413 =  ( n370 ) ? ( n371 ) : ( n412 ) ;
assign n414 =  ( n367 ) ? ( n368 ) : ( n413 ) ;
assign n415 =  ( n364 ) ? ( n365 ) : ( n414 ) ;
assign n416 =  ( n361 ) ? ( n362 ) : ( n415 ) ;
assign n417 =  ( n358 ) ? ( n359 ) : ( n416 ) ;
assign n418 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n419 =  ( n418 ) == ( bv_16_15_n111 )  ;
assign n420 = aes_counter[127:120] ;
assign n421 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n422 =  ( n421 ) == ( bv_16_14_n116 )  ;
assign n423 = aes_counter[119:112] ;
assign n424 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n425 =  ( n424 ) == ( bv_16_13_n121 )  ;
assign n426 = aes_counter[111:104] ;
assign n427 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n428 =  ( n427 ) == ( bv_16_12_n126 )  ;
assign n429 = aes_counter[103:96] ;
assign n430 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n431 =  ( n430 ) == ( bv_16_11_n131 )  ;
assign n432 = aes_counter[95:88] ;
assign n433 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n434 =  ( n433 ) == ( bv_16_10_n136 )  ;
assign n435 = aes_counter[87:80] ;
assign n436 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n437 =  ( n436 ) == ( bv_16_9_n141 )  ;
assign n438 = aes_counter[79:72] ;
assign n439 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n440 =  ( n439 ) == ( bv_16_8_n146 )  ;
assign n441 = aes_counter[71:64] ;
assign n442 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n443 =  ( n442 ) == ( bv_16_7_n151 )  ;
assign n444 = aes_counter[63:56] ;
assign n445 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n446 =  ( n445 ) == ( bv_16_6_n156 )  ;
assign n447 = aes_counter[55:48] ;
assign n448 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n449 =  ( n448 ) == ( bv_16_5_n161 )  ;
assign n450 = aes_counter[47:40] ;
assign n451 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n452 =  ( n451 ) == ( bv_16_4_n166 )  ;
assign n453 = aes_counter[39:32] ;
assign n454 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n455 =  ( n454 ) == ( bv_16_3_n171 )  ;
assign n456 = aes_counter[31:24] ;
assign n457 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n458 =  ( n457 ) == ( bv_16_2_n176 )  ;
assign n459 = aes_counter[23:16] ;
assign n460 =  ( cmdaddr ) - ( bv_16_65296_n46 )  ;
assign n461 =  ( n460 ) == ( bv_16_1_n99 )  ;
assign n462 = aes_counter[15:8] ;
assign n463 = aes_counter[7:0] ;
assign n464 =  ( n461 ) ? ( n462 ) : ( n463 ) ;
assign n465 =  ( n458 ) ? ( n459 ) : ( n464 ) ;
assign n466 =  ( n455 ) ? ( n456 ) : ( n465 ) ;
assign n467 =  ( n452 ) ? ( n453 ) : ( n466 ) ;
assign n468 =  ( n449 ) ? ( n450 ) : ( n467 ) ;
assign n469 =  ( n446 ) ? ( n447 ) : ( n468 ) ;
assign n470 =  ( n443 ) ? ( n444 ) : ( n469 ) ;
assign n471 =  ( n440 ) ? ( n441 ) : ( n470 ) ;
assign n472 =  ( n437 ) ? ( n438 ) : ( n471 ) ;
assign n473 =  ( n434 ) ? ( n435 ) : ( n472 ) ;
assign n474 =  ( n431 ) ? ( n432 ) : ( n473 ) ;
assign n475 =  ( n428 ) ? ( n429 ) : ( n474 ) ;
assign n476 =  ( n425 ) ? ( n426 ) : ( n475 ) ;
assign n477 =  ( n422 ) ? ( n423 ) : ( n476 ) ;
assign n478 =  ( n419 ) ? ( n420 ) : ( n477 ) ;
always @(posedge clk) begin
   if(rst) begin
   end
   else if(__ILA_AES_valid__) begin
       if ( __ILA_AES_decode_of_START_ENCRYPT__ && __ILA_AES_grant__[1] ) begin
           aes_status <= n85;
       end else if ( __ILA_AES_decode_of_WRITE_LENGTH__ && __ILA_AES_grant__[7] ) begin
           aes_status <= n88;
       end
       if ( __ILA_AES_decode_of_WRITE_ADDRESS__ && __ILA_AES_grant__[0] ) begin
           aes_address <= n97;
       end else if ( __ILA_AES_decode_of_READ_LENGTH__ && __ILA_AES_grant__[2] ) begin
           aes_address <= aes_address;
       end else if ( __ILA_AES_decode_of_READ_ADDRESS__ && __ILA_AES_grant__[3] ) begin
           aes_address <= aes_address;
       end else if ( __ILA_AES_decode_of_READ_KEY__ && __ILA_AES_grant__[4] ) begin
           aes_address <= aes_address;
       end else if ( __ILA_AES_decode_of_READ_COUNTER__ && __ILA_AES_grant__[5] ) begin
           aes_address <= aes_address;
       end else if ( __ILA_AES_decode_of_GET_STATUS__ && __ILA_AES_grant__[6] ) begin
           aes_address <= aes_address;
       end else if ( __ILA_AES_decode_of_WRITE_LENGTH__ && __ILA_AES_grant__[7] ) begin
           aes_address <= aes_address;
       end else if ( __ILA_AES_decode_of_WRITE_KEY__ && __ILA_AES_grant__[8] ) begin
           aes_address <= aes_address;
       end else if ( __ILA_AES_decode_of_WRITE_COUNTER__ && __ILA_AES_grant__[9] ) begin
           aes_address <= aes_address;
       end
       if ( __ILA_AES_decode_of_WRITE_ADDRESS__ && __ILA_AES_grant__[0] ) begin
           aes_length <= aes_length;
       end else if ( __ILA_AES_decode_of_READ_LENGTH__ && __ILA_AES_grant__[2] ) begin
           aes_length <= aes_length;
       end else if ( __ILA_AES_decode_of_READ_ADDRESS__ && __ILA_AES_grant__[3] ) begin
           aes_length <= aes_length;
       end else if ( __ILA_AES_decode_of_READ_KEY__ && __ILA_AES_grant__[4] ) begin
           aes_length <= aes_length;
       end else if ( __ILA_AES_decode_of_READ_COUNTER__ && __ILA_AES_grant__[5] ) begin
           aes_length <= aes_length;
       end else if ( __ILA_AES_decode_of_GET_STATUS__ && __ILA_AES_grant__[6] ) begin
           aes_length <= aes_length;
       end else if ( __ILA_AES_decode_of_WRITE_LENGTH__ && __ILA_AES_grant__[7] ) begin
           aes_length <= n109;
       end else if ( __ILA_AES_decode_of_WRITE_KEY__ && __ILA_AES_grant__[8] ) begin
           aes_length <= aes_length;
       end
       if ( __ILA_AES_decode_of_WRITE_ADDRESS__ && __ILA_AES_grant__[0] ) begin
           aes_counter <= aes_counter;
       end else if ( __ILA_AES_decode_of_WRITE_LENGTH__ && __ILA_AES_grant__[7] ) begin
           aes_counter <= aes_counter;
       end else if ( __ILA_AES_decode_of_WRITE_KEY__ && __ILA_AES_grant__[8] ) begin
           aes_counter <= aes_counter;
       end else if ( __ILA_AES_decode_of_WRITE_COUNTER__ && __ILA_AES_grant__[9] ) begin
           aes_counter <= n205;
       end
       if ( __ILA_AES_decode_of_WRITE_ADDRESS__ && __ILA_AES_grant__[0] ) begin
           aes_key <= aes_key;
       end else if ( __ILA_AES_decode_of_READ_LENGTH__ && __ILA_AES_grant__[2] ) begin
           aes_key <= aes_key;
       end else if ( __ILA_AES_decode_of_READ_ADDRESS__ && __ILA_AES_grant__[3] ) begin
           aes_key <= aes_key;
       end else if ( __ILA_AES_decode_of_READ_KEY__ && __ILA_AES_grant__[4] ) begin
           aes_key <= aes_key;
       end else if ( __ILA_AES_decode_of_READ_COUNTER__ && __ILA_AES_grant__[5] ) begin
           aes_key <= aes_key;
       end else if ( __ILA_AES_decode_of_GET_STATUS__ && __ILA_AES_grant__[6] ) begin
           aes_key <= aes_key;
       end else if ( __ILA_AES_decode_of_WRITE_LENGTH__ && __ILA_AES_grant__[7] ) begin
           aes_key <= aes_key;
       end else if ( __ILA_AES_decode_of_WRITE_KEY__ && __ILA_AES_grant__[8] ) begin
           aes_key <= n285;
       end else if ( __ILA_AES_decode_of_WRITE_COUNTER__ && __ILA_AES_grant__[9] ) begin
           aes_key <= aes_key;
       end
       if ( __ILA_AES_decode_of_READ_LENGTH__ && __ILA_AES_grant__[2] ) begin
           outdata <= n290;
       end else if ( __ILA_AES_decode_of_READ_ADDRESS__ && __ILA_AES_grant__[3] ) begin
           outdata <= n295;
       end else if ( __ILA_AES_decode_of_READ_KEY__ && __ILA_AES_grant__[4] ) begin
           outdata <= n356;
       end else if ( __ILA_AES_decode_of_READ_COUNTER__ && __ILA_AES_grant__[5] ) begin
           outdata <= n417;
       end else if ( __ILA_AES_decode_of_GET_STATUS__ && __ILA_AES_grant__[6] ) begin
           outdata <= n478;
       end
   end
end
endmodule
