module NVDLA_CMAC (
__ILA_NVDLA_CMAC_grant__,
clk,
csb_req_pd,
csb_req_valid_i,
data_i0,
data_i1,
data_i10,
data_i100,
data_i101,
data_i102,
data_i103,
data_i104,
data_i105,
data_i106,
data_i107,
data_i108,
data_i109,
data_i11,
data_i110,
data_i111,
data_i112,
data_i113,
data_i114,
data_i115,
data_i116,
data_i117,
data_i118,
data_i119,
data_i12,
data_i120,
data_i121,
data_i122,
data_i123,
data_i124,
data_i125,
data_i126,
data_i127,
data_i13,
data_i14,
data_i15,
data_i16,
data_i17,
data_i18,
data_i19,
data_i2,
data_i20,
data_i21,
data_i22,
data_i23,
data_i24,
data_i25,
data_i26,
data_i27,
data_i28,
data_i29,
data_i3,
data_i30,
data_i31,
data_i32,
data_i33,
data_i34,
data_i35,
data_i36,
data_i37,
data_i38,
data_i39,
data_i4,
data_i40,
data_i41,
data_i42,
data_i43,
data_i44,
data_i45,
data_i46,
data_i47,
data_i48,
data_i49,
data_i5,
data_i50,
data_i51,
data_i52,
data_i53,
data_i54,
data_i55,
data_i56,
data_i57,
data_i58,
data_i59,
data_i6,
data_i60,
data_i61,
data_i62,
data_i63,
data_i64,
data_i65,
data_i66,
data_i67,
data_i68,
data_i69,
data_i7,
data_i70,
data_i71,
data_i72,
data_i73,
data_i74,
data_i75,
data_i76,
data_i77,
data_i78,
data_i79,
data_i8,
data_i80,
data_i81,
data_i82,
data_i83,
data_i84,
data_i85,
data_i86,
data_i87,
data_i88,
data_i89,
data_i9,
data_i90,
data_i91,
data_i92,
data_i93,
data_i94,
data_i95,
data_i96,
data_i97,
data_i98,
data_i99,
data_mask_i,
data_pd_i,
data_valid_i,
nondet_muladd_0_n65,
nondet_muladd_1_n67,
nondet_muladd_2_n69,
nondet_muladd_3_n71,
nondet_muladd_4_n73,
nondet_muladd_5_n75,
nondet_muladd_6_n77,
nondet_muladd_7_n79,
rst,
weight_i0,
weight_i1,
weight_i10,
weight_i100,
weight_i101,
weight_i102,
weight_i103,
weight_i104,
weight_i105,
weight_i106,
weight_i107,
weight_i108,
weight_i109,
weight_i11,
weight_i110,
weight_i111,
weight_i112,
weight_i113,
weight_i114,
weight_i115,
weight_i116,
weight_i117,
weight_i118,
weight_i119,
weight_i12,
weight_i120,
weight_i121,
weight_i122,
weight_i123,
weight_i124,
weight_i125,
weight_i126,
weight_i127,
weight_i13,
weight_i14,
weight_i15,
weight_i16,
weight_i17,
weight_i18,
weight_i19,
weight_i2,
weight_i20,
weight_i21,
weight_i22,
weight_i23,
weight_i24,
weight_i25,
weight_i26,
weight_i27,
weight_i28,
weight_i29,
weight_i3,
weight_i30,
weight_i31,
weight_i32,
weight_i33,
weight_i34,
weight_i35,
weight_i36,
weight_i37,
weight_i38,
weight_i39,
weight_i4,
weight_i40,
weight_i41,
weight_i42,
weight_i43,
weight_i44,
weight_i45,
weight_i46,
weight_i47,
weight_i48,
weight_i49,
weight_i5,
weight_i50,
weight_i51,
weight_i52,
weight_i53,
weight_i54,
weight_i55,
weight_i56,
weight_i57,
weight_i58,
weight_i59,
weight_i6,
weight_i60,
weight_i61,
weight_i62,
weight_i63,
weight_i64,
weight_i65,
weight_i66,
weight_i67,
weight_i68,
weight_i69,
weight_i7,
weight_i70,
weight_i71,
weight_i72,
weight_i73,
weight_i74,
weight_i75,
weight_i76,
weight_i77,
weight_i78,
weight_i79,
weight_i8,
weight_i80,
weight_i81,
weight_i82,
weight_i83,
weight_i84,
weight_i85,
weight_i86,
weight_i87,
weight_i88,
weight_i89,
weight_i9,
weight_i90,
weight_i91,
weight_i92,
weight_i93,
weight_i94,
weight_i95,
weight_i96,
weight_i97,
weight_i98,
weight_i99,
weight_mask_i,
weight_sel_i,
weight_valid_i,
__ILA_NVDLA_CMAC_acc_decode__,
__ILA_NVDLA_CMAC_decode_of_compute__,
__ILA_NVDLA_CMAC_decode_of_set__SPACE__cfg_0__,
__ILA_NVDLA_CMAC_decode_of_set__SPACE__cfg_1__,
__ILA_NVDLA_CMAC_decode_of_set__SPACE__op_enable_0__,
__ILA_NVDLA_CMAC_decode_of_set__SPACE__op_enable_1__,
__ILA_NVDLA_CMAC_decode_of_set__SPACE__pointer__,
__ILA_NVDLA_CMAC_valid__,
producer,
consumer,
conv_mode0,
conv_mode1,
proc_precision0,
proc_precision1,
op_en0,
op_en1,
data_ready_o,
csb_req_ready_o,
csb_resp_valid_o,
csb_resp_pd_o,
data_mask_o,
data_valid_o,
act_data_o0,
act_data_o1,
act_data_o2,
act_data_o3,
act_data_o4,
act_data_o5,
act_data_o6,
act_data_o7,
act_mask_o,
act_pd_o
);
input      [5:0] __ILA_NVDLA_CMAC_grant__;
input            clk;
input     [62:0] csb_req_pd;
input            csb_req_valid_i;
input      [7:0] data_i0;
input      [7:0] data_i1;
input      [7:0] data_i10;
input      [7:0] data_i100;
input      [7:0] data_i101;
input      [7:0] data_i102;
input      [7:0] data_i103;
input      [7:0] data_i104;
input      [7:0] data_i105;
input      [7:0] data_i106;
input      [7:0] data_i107;
input      [7:0] data_i108;
input      [7:0] data_i109;
input      [7:0] data_i11;
input      [7:0] data_i110;
input      [7:0] data_i111;
input      [7:0] data_i112;
input      [7:0] data_i113;
input      [7:0] data_i114;
input      [7:0] data_i115;
input      [7:0] data_i116;
input      [7:0] data_i117;
input      [7:0] data_i118;
input      [7:0] data_i119;
input      [7:0] data_i12;
input      [7:0] data_i120;
input      [7:0] data_i121;
input      [7:0] data_i122;
input      [7:0] data_i123;
input      [7:0] data_i124;
input      [7:0] data_i125;
input      [7:0] data_i126;
input      [7:0] data_i127;
input      [7:0] data_i13;
input      [7:0] data_i14;
input      [7:0] data_i15;
input      [7:0] data_i16;
input      [7:0] data_i17;
input      [7:0] data_i18;
input      [7:0] data_i19;
input      [7:0] data_i2;
input      [7:0] data_i20;
input      [7:0] data_i21;
input      [7:0] data_i22;
input      [7:0] data_i23;
input      [7:0] data_i24;
input      [7:0] data_i25;
input      [7:0] data_i26;
input      [7:0] data_i27;
input      [7:0] data_i28;
input      [7:0] data_i29;
input      [7:0] data_i3;
input      [7:0] data_i30;
input      [7:0] data_i31;
input      [7:0] data_i32;
input      [7:0] data_i33;
input      [7:0] data_i34;
input      [7:0] data_i35;
input      [7:0] data_i36;
input      [7:0] data_i37;
input      [7:0] data_i38;
input      [7:0] data_i39;
input      [7:0] data_i4;
input      [7:0] data_i40;
input      [7:0] data_i41;
input      [7:0] data_i42;
input      [7:0] data_i43;
input      [7:0] data_i44;
input      [7:0] data_i45;
input      [7:0] data_i46;
input      [7:0] data_i47;
input      [7:0] data_i48;
input      [7:0] data_i49;
input      [7:0] data_i5;
input      [7:0] data_i50;
input      [7:0] data_i51;
input      [7:0] data_i52;
input      [7:0] data_i53;
input      [7:0] data_i54;
input      [7:0] data_i55;
input      [7:0] data_i56;
input      [7:0] data_i57;
input      [7:0] data_i58;
input      [7:0] data_i59;
input      [7:0] data_i6;
input      [7:0] data_i60;
input      [7:0] data_i61;
input      [7:0] data_i62;
input      [7:0] data_i63;
input      [7:0] data_i64;
input      [7:0] data_i65;
input      [7:0] data_i66;
input      [7:0] data_i67;
input      [7:0] data_i68;
input      [7:0] data_i69;
input      [7:0] data_i7;
input      [7:0] data_i70;
input      [7:0] data_i71;
input      [7:0] data_i72;
input      [7:0] data_i73;
input      [7:0] data_i74;
input      [7:0] data_i75;
input      [7:0] data_i76;
input      [7:0] data_i77;
input      [7:0] data_i78;
input      [7:0] data_i79;
input      [7:0] data_i8;
input      [7:0] data_i80;
input      [7:0] data_i81;
input      [7:0] data_i82;
input      [7:0] data_i83;
input      [7:0] data_i84;
input      [7:0] data_i85;
input      [7:0] data_i86;
input      [7:0] data_i87;
input      [7:0] data_i88;
input      [7:0] data_i89;
input      [7:0] data_i9;
input      [7:0] data_i90;
input      [7:0] data_i91;
input      [7:0] data_i92;
input      [7:0] data_i93;
input      [7:0] data_i94;
input      [7:0] data_i95;
input      [7:0] data_i96;
input      [7:0] data_i97;
input      [7:0] data_i98;
input      [7:0] data_i99;
input    [127:0] data_mask_i;
input      [8:0] data_pd_i;
input            data_valid_i;
input    [175:0] nondet_muladd_0_n65;
input    [175:0] nondet_muladd_1_n67;
input    [175:0] nondet_muladd_2_n69;
input    [175:0] nondet_muladd_3_n71;
input    [175:0] nondet_muladd_4_n73;
input    [175:0] nondet_muladd_5_n75;
input    [175:0] nondet_muladd_6_n77;
input    [175:0] nondet_muladd_7_n79;
input            rst;
input      [7:0] weight_i0;
input      [7:0] weight_i1;
input      [7:0] weight_i10;
input      [7:0] weight_i100;
input      [7:0] weight_i101;
input      [7:0] weight_i102;
input      [7:0] weight_i103;
input      [7:0] weight_i104;
input      [7:0] weight_i105;
input      [7:0] weight_i106;
input      [7:0] weight_i107;
input      [7:0] weight_i108;
input      [7:0] weight_i109;
input      [7:0] weight_i11;
input      [7:0] weight_i110;
input      [7:0] weight_i111;
input      [7:0] weight_i112;
input      [7:0] weight_i113;
input      [7:0] weight_i114;
input      [7:0] weight_i115;
input      [7:0] weight_i116;
input      [7:0] weight_i117;
input      [7:0] weight_i118;
input      [7:0] weight_i119;
input      [7:0] weight_i12;
input      [7:0] weight_i120;
input      [7:0] weight_i121;
input      [7:0] weight_i122;
input      [7:0] weight_i123;
input      [7:0] weight_i124;
input      [7:0] weight_i125;
input      [7:0] weight_i126;
input      [7:0] weight_i127;
input      [7:0] weight_i13;
input      [7:0] weight_i14;
input      [7:0] weight_i15;
input      [7:0] weight_i16;
input      [7:0] weight_i17;
input      [7:0] weight_i18;
input      [7:0] weight_i19;
input      [7:0] weight_i2;
input      [7:0] weight_i20;
input      [7:0] weight_i21;
input      [7:0] weight_i22;
input      [7:0] weight_i23;
input      [7:0] weight_i24;
input      [7:0] weight_i25;
input      [7:0] weight_i26;
input      [7:0] weight_i27;
input      [7:0] weight_i28;
input      [7:0] weight_i29;
input      [7:0] weight_i3;
input      [7:0] weight_i30;
input      [7:0] weight_i31;
input      [7:0] weight_i32;
input      [7:0] weight_i33;
input      [7:0] weight_i34;
input      [7:0] weight_i35;
input      [7:0] weight_i36;
input      [7:0] weight_i37;
input      [7:0] weight_i38;
input      [7:0] weight_i39;
input      [7:0] weight_i4;
input      [7:0] weight_i40;
input      [7:0] weight_i41;
input      [7:0] weight_i42;
input      [7:0] weight_i43;
input      [7:0] weight_i44;
input      [7:0] weight_i45;
input      [7:0] weight_i46;
input      [7:0] weight_i47;
input      [7:0] weight_i48;
input      [7:0] weight_i49;
input      [7:0] weight_i5;
input      [7:0] weight_i50;
input      [7:0] weight_i51;
input      [7:0] weight_i52;
input      [7:0] weight_i53;
input      [7:0] weight_i54;
input      [7:0] weight_i55;
input      [7:0] weight_i56;
input      [7:0] weight_i57;
input      [7:0] weight_i58;
input      [7:0] weight_i59;
input      [7:0] weight_i6;
input      [7:0] weight_i60;
input      [7:0] weight_i61;
input      [7:0] weight_i62;
input      [7:0] weight_i63;
input      [7:0] weight_i64;
input      [7:0] weight_i65;
input      [7:0] weight_i66;
input      [7:0] weight_i67;
input      [7:0] weight_i68;
input      [7:0] weight_i69;
input      [7:0] weight_i7;
input      [7:0] weight_i70;
input      [7:0] weight_i71;
input      [7:0] weight_i72;
input      [7:0] weight_i73;
input      [7:0] weight_i74;
input      [7:0] weight_i75;
input      [7:0] weight_i76;
input      [7:0] weight_i77;
input      [7:0] weight_i78;
input      [7:0] weight_i79;
input      [7:0] weight_i8;
input      [7:0] weight_i80;
input      [7:0] weight_i81;
input      [7:0] weight_i82;
input      [7:0] weight_i83;
input      [7:0] weight_i84;
input      [7:0] weight_i85;
input      [7:0] weight_i86;
input      [7:0] weight_i87;
input      [7:0] weight_i88;
input      [7:0] weight_i89;
input      [7:0] weight_i9;
input      [7:0] weight_i90;
input      [7:0] weight_i91;
input      [7:0] weight_i92;
input      [7:0] weight_i93;
input      [7:0] weight_i94;
input      [7:0] weight_i95;
input      [7:0] weight_i96;
input      [7:0] weight_i97;
input      [7:0] weight_i98;
input      [7:0] weight_i99;
input    [127:0] weight_mask_i;
input      [7:0] weight_sel_i;
input            weight_valid_i;
output      [5:0] __ILA_NVDLA_CMAC_acc_decode__;
output            __ILA_NVDLA_CMAC_decode_of_compute__;
output            __ILA_NVDLA_CMAC_decode_of_set__SPACE__cfg_0__;
output            __ILA_NVDLA_CMAC_decode_of_set__SPACE__cfg_1__;
output            __ILA_NVDLA_CMAC_decode_of_set__SPACE__op_enable_0__;
output            __ILA_NVDLA_CMAC_decode_of_set__SPACE__op_enable_1__;
output            __ILA_NVDLA_CMAC_decode_of_set__SPACE__pointer__;
output            __ILA_NVDLA_CMAC_valid__;
output reg            producer;
output reg            consumer;
output reg            conv_mode0;
output reg            conv_mode1;
output reg      [1:0] proc_precision0;
output reg      [1:0] proc_precision1;
output reg            op_en0;
output reg            op_en1;
output reg            data_ready_o;
output reg            csb_req_ready_o;
output reg            csb_resp_valid_o;
output reg     [33:0] csb_resp_pd_o;
output reg    [127:0] data_mask_o;
output reg            data_valid_o;
output reg    [175:0] act_data_o0;
output reg    [175:0] act_data_o1;
output reg    [175:0] act_data_o2;
output reg    [175:0] act_data_o3;
output reg    [175:0] act_data_o4;
output reg    [175:0] act_data_o5;
output reg    [175:0] act_data_o6;
output reg    [175:0] act_data_o7;
output reg      [7:0] act_mask_o;
output reg      [8:0] act_pd_o;
wire      [5:0] __ILA_NVDLA_CMAC_acc_decode__;
wire            __ILA_NVDLA_CMAC_decode_of_compute__;
wire            __ILA_NVDLA_CMAC_decode_of_set__SPACE__cfg_0__;
wire            __ILA_NVDLA_CMAC_decode_of_set__SPACE__cfg_1__;
wire            __ILA_NVDLA_CMAC_decode_of_set__SPACE__op_enable_0__;
wire            __ILA_NVDLA_CMAC_decode_of_set__SPACE__op_enable_1__;
wire            __ILA_NVDLA_CMAC_decode_of_set__SPACE__pointer__;
wire      [5:0] __ILA_NVDLA_CMAC_grant__;
wire            __ILA_NVDLA_CMAC_valid__;
wire     [11:0] bv_12_12_n25;
wire     [11:0] bv_12_4_n5;
wire     [11:0] bv_12_8_n14;
wire            bv_1_1_n8;
wire      [1:0] bv_2_0_n2;
wire      [7:0] bv_8_255_n81;
wire            clk;
wire     [62:0] csb_req_pd;
wire            csb_req_valid_i;
wire      [7:0] data_i0;
wire      [7:0] data_i1;
wire      [7:0] data_i10;
wire      [7:0] data_i100;
wire      [7:0] data_i101;
wire      [7:0] data_i102;
wire      [7:0] data_i103;
wire      [7:0] data_i104;
wire      [7:0] data_i105;
wire      [7:0] data_i106;
wire      [7:0] data_i107;
wire      [7:0] data_i108;
wire      [7:0] data_i109;
wire      [7:0] data_i11;
wire      [7:0] data_i110;
wire      [7:0] data_i111;
wire      [7:0] data_i112;
wire      [7:0] data_i113;
wire      [7:0] data_i114;
wire      [7:0] data_i115;
wire      [7:0] data_i116;
wire      [7:0] data_i117;
wire      [7:0] data_i118;
wire      [7:0] data_i119;
wire      [7:0] data_i12;
wire      [7:0] data_i120;
wire      [7:0] data_i121;
wire      [7:0] data_i122;
wire      [7:0] data_i123;
wire      [7:0] data_i124;
wire      [7:0] data_i125;
wire      [7:0] data_i126;
wire      [7:0] data_i127;
wire      [7:0] data_i13;
wire      [7:0] data_i14;
wire      [7:0] data_i15;
wire      [7:0] data_i16;
wire      [7:0] data_i17;
wire      [7:0] data_i18;
wire      [7:0] data_i19;
wire      [7:0] data_i2;
wire      [7:0] data_i20;
wire      [7:0] data_i21;
wire      [7:0] data_i22;
wire      [7:0] data_i23;
wire      [7:0] data_i24;
wire      [7:0] data_i25;
wire      [7:0] data_i26;
wire      [7:0] data_i27;
wire      [7:0] data_i28;
wire      [7:0] data_i29;
wire      [7:0] data_i3;
wire      [7:0] data_i30;
wire      [7:0] data_i31;
wire      [7:0] data_i32;
wire      [7:0] data_i33;
wire      [7:0] data_i34;
wire      [7:0] data_i35;
wire      [7:0] data_i36;
wire      [7:0] data_i37;
wire      [7:0] data_i38;
wire      [7:0] data_i39;
wire      [7:0] data_i4;
wire      [7:0] data_i40;
wire      [7:0] data_i41;
wire      [7:0] data_i42;
wire      [7:0] data_i43;
wire      [7:0] data_i44;
wire      [7:0] data_i45;
wire      [7:0] data_i46;
wire      [7:0] data_i47;
wire      [7:0] data_i48;
wire      [7:0] data_i49;
wire      [7:0] data_i5;
wire      [7:0] data_i50;
wire      [7:0] data_i51;
wire      [7:0] data_i52;
wire      [7:0] data_i53;
wire      [7:0] data_i54;
wire      [7:0] data_i55;
wire      [7:0] data_i56;
wire      [7:0] data_i57;
wire      [7:0] data_i58;
wire      [7:0] data_i59;
wire      [7:0] data_i6;
wire      [7:0] data_i60;
wire      [7:0] data_i61;
wire      [7:0] data_i62;
wire      [7:0] data_i63;
wire      [7:0] data_i64;
wire      [7:0] data_i65;
wire      [7:0] data_i66;
wire      [7:0] data_i67;
wire      [7:0] data_i68;
wire      [7:0] data_i69;
wire      [7:0] data_i7;
wire      [7:0] data_i70;
wire      [7:0] data_i71;
wire      [7:0] data_i72;
wire      [7:0] data_i73;
wire      [7:0] data_i74;
wire      [7:0] data_i75;
wire      [7:0] data_i76;
wire      [7:0] data_i77;
wire      [7:0] data_i78;
wire      [7:0] data_i79;
wire      [7:0] data_i8;
wire      [7:0] data_i80;
wire      [7:0] data_i81;
wire      [7:0] data_i82;
wire      [7:0] data_i83;
wire      [7:0] data_i84;
wire      [7:0] data_i85;
wire      [7:0] data_i86;
wire      [7:0] data_i87;
wire      [7:0] data_i88;
wire      [7:0] data_i89;
wire      [7:0] data_i9;
wire      [7:0] data_i90;
wire      [7:0] data_i91;
wire      [7:0] data_i92;
wire      [7:0] data_i93;
wire      [7:0] data_i94;
wire      [7:0] data_i95;
wire      [7:0] data_i96;
wire      [7:0] data_i97;
wire      [7:0] data_i98;
wire      [7:0] data_i99;
wire    [127:0] data_mask_i;
wire      [8:0] data_pd_i;
wire            data_valid_i;
wire     [21:0] n0;
wire     [21:0] n1;
wire            n10;
wire            n11;
wire            n12;
wire     [11:0] n13;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire     [11:0] n24;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire     [23:0] n3;
wire            n30;
wire            n31;
wire            n32;
wire            n33;
wire            n34;
wire     [11:0] n35;
wire            n36;
wire            n37;
wire            n38;
wire            n39;
wire     [11:0] n4;
wire            n40;
wire            n41;
wire            n42;
wire            n43;
wire            n44;
wire     [11:0] n45;
wire            n46;
wire            n47;
wire            n48;
wire            n49;
wire            n50;
wire            n51;
wire            n52;
wire            n53;
wire            n54;
wire            n55;
wire            n56;
wire     [31:0] n57;
wire            n58;
wire            n59;
wire            n6;
wire            n60;
wire      [1:0] n61;
wire      [1:0] n62;
wire            n63;
wire            n64;
wire    [175:0] n66;
wire    [175:0] n68;
wire            n7;
wire    [175:0] n70;
wire    [175:0] n72;
wire    [175:0] n74;
wire    [175:0] n76;
wire    [175:0] n78;
wire    [175:0] n80;
wire            n9;
wire    [175:0] nondet_muladd_0_n65;
wire    [175:0] nondet_muladd_1_n67;
wire    [175:0] nondet_muladd_2_n69;
wire    [175:0] nondet_muladd_3_n71;
wire    [175:0] nondet_muladd_4_n73;
wire    [175:0] nondet_muladd_5_n75;
wire    [175:0] nondet_muladd_6_n77;
wire    [175:0] nondet_muladd_7_n79;
wire            rst;
wire      [7:0] weight_i0;
wire      [7:0] weight_i1;
wire      [7:0] weight_i10;
wire      [7:0] weight_i100;
wire      [7:0] weight_i101;
wire      [7:0] weight_i102;
wire      [7:0] weight_i103;
wire      [7:0] weight_i104;
wire      [7:0] weight_i105;
wire      [7:0] weight_i106;
wire      [7:0] weight_i107;
wire      [7:0] weight_i108;
wire      [7:0] weight_i109;
wire      [7:0] weight_i11;
wire      [7:0] weight_i110;
wire      [7:0] weight_i111;
wire      [7:0] weight_i112;
wire      [7:0] weight_i113;
wire      [7:0] weight_i114;
wire      [7:0] weight_i115;
wire      [7:0] weight_i116;
wire      [7:0] weight_i117;
wire      [7:0] weight_i118;
wire      [7:0] weight_i119;
wire      [7:0] weight_i12;
wire      [7:0] weight_i120;
wire      [7:0] weight_i121;
wire      [7:0] weight_i122;
wire      [7:0] weight_i123;
wire      [7:0] weight_i124;
wire      [7:0] weight_i125;
wire      [7:0] weight_i126;
wire      [7:0] weight_i127;
wire      [7:0] weight_i13;
wire      [7:0] weight_i14;
wire      [7:0] weight_i15;
wire      [7:0] weight_i16;
wire      [7:0] weight_i17;
wire      [7:0] weight_i18;
wire      [7:0] weight_i19;
wire      [7:0] weight_i2;
wire      [7:0] weight_i20;
wire      [7:0] weight_i21;
wire      [7:0] weight_i22;
wire      [7:0] weight_i23;
wire      [7:0] weight_i24;
wire      [7:0] weight_i25;
wire      [7:0] weight_i26;
wire      [7:0] weight_i27;
wire      [7:0] weight_i28;
wire      [7:0] weight_i29;
wire      [7:0] weight_i3;
wire      [7:0] weight_i30;
wire      [7:0] weight_i31;
wire      [7:0] weight_i32;
wire      [7:0] weight_i33;
wire      [7:0] weight_i34;
wire      [7:0] weight_i35;
wire      [7:0] weight_i36;
wire      [7:0] weight_i37;
wire      [7:0] weight_i38;
wire      [7:0] weight_i39;
wire      [7:0] weight_i4;
wire      [7:0] weight_i40;
wire      [7:0] weight_i41;
wire      [7:0] weight_i42;
wire      [7:0] weight_i43;
wire      [7:0] weight_i44;
wire      [7:0] weight_i45;
wire      [7:0] weight_i46;
wire      [7:0] weight_i47;
wire      [7:0] weight_i48;
wire      [7:0] weight_i49;
wire      [7:0] weight_i5;
wire      [7:0] weight_i50;
wire      [7:0] weight_i51;
wire      [7:0] weight_i52;
wire      [7:0] weight_i53;
wire      [7:0] weight_i54;
wire      [7:0] weight_i55;
wire      [7:0] weight_i56;
wire      [7:0] weight_i57;
wire      [7:0] weight_i58;
wire      [7:0] weight_i59;
wire      [7:0] weight_i6;
wire      [7:0] weight_i60;
wire      [7:0] weight_i61;
wire      [7:0] weight_i62;
wire      [7:0] weight_i63;
wire      [7:0] weight_i64;
wire      [7:0] weight_i65;
wire      [7:0] weight_i66;
wire      [7:0] weight_i67;
wire      [7:0] weight_i68;
wire      [7:0] weight_i69;
wire      [7:0] weight_i7;
wire      [7:0] weight_i70;
wire      [7:0] weight_i71;
wire      [7:0] weight_i72;
wire      [7:0] weight_i73;
wire      [7:0] weight_i74;
wire      [7:0] weight_i75;
wire      [7:0] weight_i76;
wire      [7:0] weight_i77;
wire      [7:0] weight_i78;
wire      [7:0] weight_i79;
wire      [7:0] weight_i8;
wire      [7:0] weight_i80;
wire      [7:0] weight_i81;
wire      [7:0] weight_i82;
wire      [7:0] weight_i83;
wire      [7:0] weight_i84;
wire      [7:0] weight_i85;
wire      [7:0] weight_i86;
wire      [7:0] weight_i87;
wire      [7:0] weight_i88;
wire      [7:0] weight_i89;
wire      [7:0] weight_i9;
wire      [7:0] weight_i90;
wire      [7:0] weight_i91;
wire      [7:0] weight_i92;
wire      [7:0] weight_i93;
wire      [7:0] weight_i94;
wire      [7:0] weight_i95;
wire      [7:0] weight_i96;
wire      [7:0] weight_i97;
wire      [7:0] weight_i98;
wire      [7:0] weight_i99;
wire    [127:0] weight_mask_i;
wire      [7:0] weight_sel_i;
wire            weight_valid_i;
assign __ILA_NVDLA_CMAC_valid__ = 1'b1 ;
assign n0 = csb_req_pd[21:0] ;
assign n1 = n0[21:0] ;
assign bv_2_0_n2 = 2'h0 ;
assign n3 =  { ( n1 ) , ( bv_2_0_n2 ) }  ;
assign n4 = n3[11:0] ;
assign bv_12_4_n5 = 12'h4 ;
assign n6 =  ( n4 ) == ( bv_12_4_n5 )  ;
assign n7 = csb_req_pd[54:54] ;
assign bv_1_1_n8 = 1'h1 ;
assign n9 =  ( n7 ) == ( bv_1_1_n8 )  ;
assign n10 =  ( n6 ) & (n9 )  ;
assign n11 =  ( n10 ) & (csb_req_valid_i )  ;
assign n12 =  ( n11 ) & (csb_req_ready_o )  ;
assign __ILA_NVDLA_CMAC_decode_of_set__SPACE__pointer__ = n12 ;
assign __ILA_NVDLA_CMAC_acc_decode__[0] = __ILA_NVDLA_CMAC_decode_of_set__SPACE__pointer__ ;
assign n13 = n3[11:0] ;
assign bv_12_8_n14 = 12'h8 ;
assign n15 =  ( n13 ) == ( bv_12_8_n14 )  ;
assign n16 =  ( producer ) == ( 1'b0 )  ;
assign n17 =  ( n15 ) & (n16 )  ;
assign n18 =  ( op_en0 ) == ( 1'b0 )  ;
assign n19 =  ( n17 ) & (n18 )  ;
assign n20 =  ( n7 ) == ( bv_1_1_n8 )  ;
assign n21 =  ( n19 ) & (n20 )  ;
assign n22 =  ( n21 ) & (csb_req_valid_i )  ;
assign n23 =  ( n22 ) & (csb_req_ready_o )  ;
assign __ILA_NVDLA_CMAC_decode_of_set__SPACE__op_enable_0__ = n23 ;
assign __ILA_NVDLA_CMAC_acc_decode__[1] = __ILA_NVDLA_CMAC_decode_of_set__SPACE__op_enable_0__ ;
assign n24 = n3[11:0] ;
assign bv_12_12_n25 = 12'hc ;
assign n26 =  ( n24 ) == ( bv_12_12_n25 )  ;
assign n27 =  ( producer ) == ( 1'b0 )  ;
assign n28 =  ( n26 ) & (n27 )  ;
assign n29 =  ( op_en0 ) == ( 1'b0 )  ;
assign n30 =  ( n28 ) & (n29 )  ;
assign n31 =  ( n7 ) == ( bv_1_1_n8 )  ;
assign n32 =  ( n30 ) & (n31 )  ;
assign n33 =  ( n32 ) & (csb_req_valid_i )  ;
assign n34 =  ( n33 ) & (csb_req_ready_o )  ;
assign __ILA_NVDLA_CMAC_decode_of_set__SPACE__cfg_0__ = n34 ;
assign __ILA_NVDLA_CMAC_acc_decode__[2] = __ILA_NVDLA_CMAC_decode_of_set__SPACE__cfg_0__ ;
assign n35 = n3[11:0] ;
assign n36 =  ( n35 ) == ( bv_12_8_n14 )  ;
assign n37 =  ( producer ) == ( 1'b1 )  ;
assign n38 =  ( n36 ) & (n37 )  ;
assign n39 =  ( op_en1 ) == ( 1'b0 )  ;
assign n40 =  ( n38 ) & (n39 )  ;
assign n41 =  ( n7 ) == ( bv_1_1_n8 )  ;
assign n42 =  ( n40 ) & (n41 )  ;
assign n43 =  ( n42 ) & (csb_req_valid_i )  ;
assign n44 =  ( n43 ) & (csb_req_ready_o )  ;
assign __ILA_NVDLA_CMAC_decode_of_set__SPACE__op_enable_1__ = n44 ;
assign __ILA_NVDLA_CMAC_acc_decode__[3] = __ILA_NVDLA_CMAC_decode_of_set__SPACE__op_enable_1__ ;
assign n45 = n3[11:0] ;
assign n46 =  ( n45 ) == ( bv_12_12_n25 )  ;
assign n47 =  ( producer ) == ( 1'b1 )  ;
assign n48 =  ( n46 ) & (n47 )  ;
assign n49 =  ( op_en1 ) == ( 1'b0 )  ;
assign n50 =  ( n48 ) & (n49 )  ;
assign n51 =  ( n7 ) == ( bv_1_1_n8 )  ;
assign n52 =  ( n50 ) & (n51 )  ;
assign n53 =  ( n52 ) & (csb_req_valid_i )  ;
assign n54 =  ( n53 ) & (csb_req_ready_o )  ;
assign __ILA_NVDLA_CMAC_decode_of_set__SPACE__cfg_1__ = n54 ;
assign __ILA_NVDLA_CMAC_acc_decode__[4] = __ILA_NVDLA_CMAC_decode_of_set__SPACE__cfg_1__ ;
assign n55 =  ( data_valid_i ) & (weight_valid_i )  ;
assign n56 =  ( n55 ) & (data_ready_o )  ;
assign __ILA_NVDLA_CMAC_decode_of_compute__ = n56 ;
assign __ILA_NVDLA_CMAC_acc_decode__[5] = __ILA_NVDLA_CMAC_decode_of_compute__ ;
assign n57 = csb_req_pd[53:22] ;
assign n58 = n57[0:0] ;
assign n59 = n57[0:0] ;
assign n60 = n57[0:0] ;
assign n61 = n57[13:12] ;
assign n62 = n57[13:12] ;
assign n63 = n57[0:0] ;
assign n64 = n57[0:0] ;
assign n66 = nondet_muladd_0_n65 ;
assign n68 = nondet_muladd_1_n67 ;
assign n70 = nondet_muladd_2_n69 ;
assign n72 = nondet_muladd_3_n71 ;
assign n74 = nondet_muladd_4_n73 ;
assign n76 = nondet_muladd_5_n75 ;
assign n78 = nondet_muladd_6_n77 ;
assign n80 = nondet_muladd_7_n79 ;
assign bv_8_255_n81 = 8'hff ;
always @(posedge clk) begin
   if(rst) begin
   end
   else if(__ILA_NVDLA_CMAC_valid__) begin
       if ( __ILA_NVDLA_CMAC_decode_of_set__SPACE__pointer__ && __ILA_NVDLA_CMAC_grant__[0] ) begin
           producer <= n58;
       end
       if ( __ILA_NVDLA_CMAC_decode_of_set__SPACE__cfg_0__ && __ILA_NVDLA_CMAC_grant__[2] ) begin
           conv_mode0 <= n59;
       end
       if ( __ILA_NVDLA_CMAC_decode_of_set__SPACE__cfg_1__ && __ILA_NVDLA_CMAC_grant__[4] ) begin
           conv_mode1 <= n60;
       end
       if ( __ILA_NVDLA_CMAC_decode_of_set__SPACE__cfg_0__ && __ILA_NVDLA_CMAC_grant__[2] ) begin
           proc_precision0 <= n61;
       end
       if ( __ILA_NVDLA_CMAC_decode_of_set__SPACE__cfg_1__ && __ILA_NVDLA_CMAC_grant__[4] ) begin
           proc_precision1 <= n62;
       end
       if ( __ILA_NVDLA_CMAC_decode_of_set__SPACE__op_enable_0__ && __ILA_NVDLA_CMAC_grant__[1] ) begin
           op_en0 <= n63;
       end
       if ( __ILA_NVDLA_CMAC_decode_of_set__SPACE__op_enable_1__ && __ILA_NVDLA_CMAC_grant__[3] ) begin
           op_en1 <= n64;
       end
       if ( __ILA_NVDLA_CMAC_decode_of_compute__ && __ILA_NVDLA_CMAC_grant__[5] ) begin
           data_valid_o <= data_valid_i;
       end
       if ( __ILA_NVDLA_CMAC_decode_of_compute__ && __ILA_NVDLA_CMAC_grant__[5] ) begin
           act_data_o0 <= n66;
       end
       if ( __ILA_NVDLA_CMAC_decode_of_compute__ && __ILA_NVDLA_CMAC_grant__[5] ) begin
           act_data_o1 <= n68;
       end
       if ( __ILA_NVDLA_CMAC_decode_of_compute__ && __ILA_NVDLA_CMAC_grant__[5] ) begin
           act_data_o2 <= n70;
       end
       if ( __ILA_NVDLA_CMAC_decode_of_compute__ && __ILA_NVDLA_CMAC_grant__[5] ) begin
           act_data_o3 <= n72;
       end
       if ( __ILA_NVDLA_CMAC_decode_of_compute__ && __ILA_NVDLA_CMAC_grant__[5] ) begin
           act_data_o4 <= n74;
       end
       if ( __ILA_NVDLA_CMAC_decode_of_compute__ && __ILA_NVDLA_CMAC_grant__[5] ) begin
           act_data_o5 <= n76;
       end
       if ( __ILA_NVDLA_CMAC_decode_of_compute__ && __ILA_NVDLA_CMAC_grant__[5] ) begin
           act_data_o6 <= n78;
       end
       if ( __ILA_NVDLA_CMAC_decode_of_compute__ && __ILA_NVDLA_CMAC_grant__[5] ) begin
           act_data_o7 <= n80;
       end
       if ( __ILA_NVDLA_CMAC_decode_of_compute__ && __ILA_NVDLA_CMAC_grant__[5] ) begin
           act_mask_o <= bv_8_255_n81;
       end
       if ( __ILA_NVDLA_CMAC_decode_of_compute__ && __ILA_NVDLA_CMAC_grant__[5] ) begin
           act_pd_o <= data_pd_i;
       end
   end
end
endmodule
